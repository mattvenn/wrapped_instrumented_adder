magic
tech sky130A
magscale 1 2
timestamp 1654174883
<< viali >>
rect 13369 47209 13403 47243
rect 19441 47141 19475 47175
rect 29929 47141 29963 47175
rect 48145 47141 48179 47175
rect 20085 47073 20119 47107
rect 30757 47073 30791 47107
rect 47041 47073 47075 47107
rect 2053 47005 2087 47039
rect 2973 47005 3007 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6837 47005 6871 47039
rect 7757 47005 7791 47039
rect 9137 47005 9171 47039
rect 11713 47005 11747 47039
rect 11989 47005 12023 47039
rect 13093 47005 13127 47039
rect 15301 47005 15335 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 19257 47005 19291 47039
rect 20361 47005 20395 47039
rect 24777 47005 24811 47039
rect 25421 47005 25455 47039
rect 28641 47005 28675 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38301 47005 38335 47039
rect 41889 47005 41923 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47961 47005 47995 47039
rect 2329 46937 2363 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 7941 46937 7975 46971
rect 14565 46937 14599 46971
rect 14749 46937 14783 46971
rect 15485 46937 15519 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 42809 46937 42843 46971
rect 44465 46937 44499 46971
rect 45385 46937 45419 46971
rect 3157 46869 3191 46903
rect 6929 46869 6963 46903
rect 9321 46869 9355 46903
rect 28457 46869 28491 46903
rect 28457 46597 28491 46631
rect 30113 46597 30147 46631
rect 1409 46529 1443 46563
rect 24593 46529 24627 46563
rect 28273 46529 28307 46563
rect 38117 46529 38151 46563
rect 41705 46529 41739 46563
rect 42441 46529 42475 46563
rect 47869 46529 47903 46563
rect 2973 46461 3007 46495
rect 3433 46461 3467 46495
rect 3617 46461 3651 46495
rect 4169 46461 4203 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 11989 46461 12023 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19441 46461 19475 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41797 46461 41831 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 1593 46325 1627 46359
rect 2329 46325 2363 46359
rect 22017 46325 22051 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 3893 46121 3927 46155
rect 11253 46121 11287 46155
rect 14289 46121 14323 46155
rect 20177 46121 20211 46155
rect 24685 46121 24719 46155
rect 38301 46121 38335 46155
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41337 45985 41371 46019
rect 41981 45985 42015 46019
rect 47041 45985 47075 46019
rect 2789 45917 2823 45951
rect 3801 45917 3835 45951
rect 11161 45917 11195 45951
rect 20085 45917 20119 45951
rect 24593 45917 24627 45951
rect 38209 45917 38243 45951
rect 44005 45917 44039 45951
rect 45569 45917 45603 45951
rect 46305 45917 46339 45951
rect 20913 45849 20947 45883
rect 25421 45849 25455 45883
rect 41521 45849 41555 45883
rect 46489 45849 46523 45883
rect 2881 45781 2915 45815
rect 44097 45781 44131 45815
rect 45753 45781 45787 45815
rect 13829 45577 13863 45611
rect 20913 45577 20947 45611
rect 25329 45577 25363 45611
rect 32229 45577 32263 45611
rect 41429 45577 41463 45611
rect 2145 45509 2179 45543
rect 42809 45509 42843 45543
rect 46949 45509 46983 45543
rect 47961 45509 47995 45543
rect 1961 45441 1995 45475
rect 13737 45441 13771 45475
rect 20269 45441 20303 45475
rect 20821 45441 20855 45475
rect 25237 45441 25271 45475
rect 32137 45441 32171 45475
rect 41337 45441 41371 45475
rect 42717 45441 42751 45475
rect 43821 45441 43855 45475
rect 46857 45441 46891 45475
rect 2789 45373 2823 45407
rect 44557 45373 44591 45407
rect 44741 45373 44775 45407
rect 45661 45373 45695 45407
rect 44005 45237 44039 45271
rect 48053 45237 48087 45271
rect 42901 45033 42935 45067
rect 44465 45033 44499 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 46949 44489 46983 44523
rect 45109 44353 45143 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 47685 44149 47719 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 47777 43265 47811 43299
rect 1593 43197 1627 43231
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 2237 41225 2271 41259
rect 46857 41225 46891 41259
rect 2145 41089 2179 41123
rect 46765 41089 46799 41123
rect 47961 41089 47995 41123
rect 48145 40953 48179 40987
rect 47685 40681 47719 40715
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 47777 39797 47811 39831
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 46489 39321 46523 39355
rect 46949 39049 46983 39083
rect 46857 38913 46891 38947
rect 47685 38913 47719 38947
rect 47869 38845 47903 38879
rect 26617 38505 26651 38539
rect 27537 38369 27571 38403
rect 22661 38301 22695 38335
rect 26341 38301 26375 38335
rect 27353 38301 27387 38335
rect 46305 38301 46339 38335
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 22477 38165 22511 38199
rect 26157 38165 26191 38199
rect 26985 38165 27019 38199
rect 27445 38165 27479 38199
rect 47685 37961 47719 37995
rect 22845 37893 22879 37927
rect 27261 37893 27295 37927
rect 47593 37825 47627 37859
rect 22569 37757 22603 37791
rect 26985 37757 27019 37791
rect 28733 37757 28767 37791
rect 24317 37621 24351 37655
rect 22293 37417 22327 37451
rect 24961 37417 24995 37451
rect 27353 37417 27387 37451
rect 47685 37417 47719 37451
rect 22937 37281 22971 37315
rect 24501 37281 24535 37315
rect 26985 37281 27019 37315
rect 23673 37213 23707 37247
rect 23765 37213 23799 37247
rect 24593 37213 24627 37247
rect 25421 37213 25455 37247
rect 27077 37213 27111 37247
rect 27905 37213 27939 37247
rect 27997 37213 28031 37247
rect 22661 37145 22695 37179
rect 22753 37145 22787 37179
rect 25513 37077 25547 37111
rect 28549 36737 28583 36771
rect 24501 36669 24535 36703
rect 24777 36669 24811 36703
rect 28825 36669 28859 36703
rect 26249 36533 26283 36567
rect 30297 36533 30331 36567
rect 24501 36329 24535 36363
rect 26157 36329 26191 36363
rect 28457 36329 28491 36363
rect 29745 36329 29779 36363
rect 2789 36193 2823 36227
rect 21741 36193 21775 36227
rect 22661 36193 22695 36227
rect 25789 36193 25823 36227
rect 27077 36193 27111 36227
rect 1409 36125 1443 36159
rect 21005 36125 21039 36159
rect 22385 36125 22419 36159
rect 24501 36125 24535 36159
rect 24685 36125 24719 36159
rect 25421 36125 25455 36159
rect 25605 36125 25639 36159
rect 25697 36125 25731 36159
rect 25973 36125 26007 36159
rect 26801 36125 26835 36159
rect 26985 36125 27019 36159
rect 28089 36125 28123 36159
rect 28457 36125 28491 36159
rect 29653 36125 29687 36159
rect 1593 36057 1627 36091
rect 20821 35989 20855 36023
rect 22017 35989 22051 36023
rect 22477 35989 22511 36023
rect 26617 35989 26651 36023
rect 28641 35989 28675 36023
rect 25237 35785 25271 35819
rect 26249 35785 26283 35819
rect 28825 35785 28859 35819
rect 29285 35785 29319 35819
rect 27169 35717 27203 35751
rect 31493 35717 31527 35751
rect 2053 35649 2087 35683
rect 22017 35649 22051 35683
rect 24869 35649 24903 35683
rect 25697 35649 25731 35683
rect 26065 35649 26099 35683
rect 27445 35649 27479 35683
rect 28089 35649 28123 35683
rect 28273 35649 28307 35683
rect 28365 35649 28399 35683
rect 28641 35649 28675 35683
rect 29469 35649 29503 35683
rect 31401 35649 31435 35683
rect 19533 35581 19567 35615
rect 19809 35581 19843 35615
rect 21281 35581 21315 35615
rect 21925 35581 21959 35615
rect 22385 35581 22419 35615
rect 24961 35581 24995 35615
rect 27353 35581 27387 35615
rect 28457 35581 28491 35615
rect 29745 35581 29779 35615
rect 32137 35581 32171 35615
rect 32413 35581 32447 35615
rect 25053 35445 25087 35479
rect 25789 35445 25823 35479
rect 27169 35445 27203 35479
rect 27629 35445 27663 35479
rect 29653 35445 29687 35479
rect 33885 35445 33919 35479
rect 2237 35241 2271 35275
rect 19993 35241 20027 35275
rect 28181 35241 28215 35275
rect 32873 35241 32907 35275
rect 23397 35105 23431 35139
rect 27445 35105 27479 35139
rect 27997 35105 28031 35139
rect 29653 35105 29687 35139
rect 31953 35105 31987 35139
rect 33333 35105 33367 35139
rect 35081 35105 35115 35139
rect 1593 35037 1627 35071
rect 2145 35037 2179 35071
rect 19901 35037 19935 35071
rect 23305 35037 23339 35071
rect 24409 35037 24443 35071
rect 26065 35037 26099 35071
rect 26249 35037 26283 35071
rect 27077 35037 27111 35071
rect 27261 35037 27295 35071
rect 27905 35037 27939 35071
rect 28181 35037 28215 35071
rect 32045 35037 32079 35071
rect 33057 35037 33091 35071
rect 33241 35037 33275 35071
rect 34897 35037 34931 35071
rect 35173 35037 35207 35071
rect 35633 35037 35667 35071
rect 47317 35037 47351 35071
rect 47593 35037 47627 35071
rect 29929 34969 29963 35003
rect 1409 34901 1443 34935
rect 23673 34901 23707 34935
rect 24593 34901 24627 34935
rect 26433 34901 26467 34935
rect 28365 34901 28399 34935
rect 31401 34901 31435 34935
rect 32413 34901 32447 34935
rect 34713 34901 34747 34935
rect 35725 34901 35759 34935
rect 25973 34697 26007 34731
rect 27721 34697 27755 34731
rect 29561 34697 29595 34731
rect 30941 34697 30975 34731
rect 32873 34697 32907 34731
rect 23305 34629 23339 34663
rect 23521 34629 23555 34663
rect 27261 34629 27295 34663
rect 34253 34629 34287 34663
rect 18797 34561 18831 34595
rect 27537 34561 27571 34595
rect 28273 34561 28307 34595
rect 29745 34561 29779 34595
rect 30849 34561 30883 34595
rect 33057 34561 33091 34595
rect 33149 34561 33183 34595
rect 33425 34561 33459 34595
rect 48145 34561 48179 34595
rect 24225 34493 24259 34527
rect 27353 34493 27387 34527
rect 28549 34493 28583 34527
rect 30021 34493 30055 34527
rect 33977 34493 34011 34527
rect 33333 34425 33367 34459
rect 18981 34357 19015 34391
rect 23489 34357 23523 34391
rect 23673 34357 23707 34391
rect 24482 34357 24516 34391
rect 27537 34357 27571 34391
rect 29929 34357 29963 34391
rect 35725 34357 35759 34391
rect 47961 34357 47995 34391
rect 22385 34153 22419 34187
rect 25789 34153 25823 34187
rect 35173 34153 35207 34187
rect 35725 34153 35759 34187
rect 27169 34085 27203 34119
rect 29009 34085 29043 34119
rect 28549 34017 28583 34051
rect 34805 34017 34839 34051
rect 36185 34017 36219 34051
rect 46305 34017 46339 34051
rect 19349 33949 19383 33983
rect 20637 33949 20671 33983
rect 20730 33949 20764 33983
rect 20913 33949 20947 33983
rect 21102 33949 21136 33983
rect 21741 33949 21775 33983
rect 21889 33949 21923 33983
rect 22206 33949 22240 33983
rect 23213 33949 23247 33983
rect 23361 33949 23395 33983
rect 23489 33949 23523 33983
rect 23581 33949 23615 33983
rect 23719 33949 23753 33983
rect 25697 33949 25731 33983
rect 26801 33949 26835 33983
rect 28641 33949 28675 33983
rect 34897 33949 34931 33983
rect 35909 33949 35943 33983
rect 36001 33949 36035 33983
rect 36277 33949 36311 33983
rect 21005 33881 21039 33915
rect 22017 33881 22051 33915
rect 22109 33881 22143 33915
rect 26985 33881 27019 33915
rect 46489 33881 46523 33915
rect 48145 33881 48179 33915
rect 19441 33813 19475 33847
rect 21281 33813 21315 33847
rect 23857 33813 23891 33847
rect 24593 33609 24627 33643
rect 28641 33609 28675 33643
rect 48053 33609 48087 33643
rect 20913 33541 20947 33575
rect 21129 33541 21163 33575
rect 22109 33541 22143 33575
rect 25881 33541 25915 33575
rect 18521 33473 18555 33507
rect 21833 33473 21867 33507
rect 24133 33473 24167 33507
rect 24409 33473 24443 33507
rect 26065 33473 26099 33507
rect 27537 33473 27571 33507
rect 27629 33473 27663 33507
rect 28273 33473 28307 33507
rect 34713 33473 34747 33507
rect 47869 33473 47903 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 18797 33405 18831 33439
rect 24317 33405 24351 33439
rect 27813 33405 27847 33439
rect 28365 33405 28399 33439
rect 34989 33405 35023 33439
rect 26249 33337 26283 33371
rect 34805 33337 34839 33371
rect 20269 33269 20303 33303
rect 21097 33269 21131 33303
rect 21281 33269 21315 33303
rect 23581 33269 23615 33303
rect 24409 33269 24443 33303
rect 27721 33269 27755 33303
rect 28365 33269 28399 33303
rect 34897 33269 34931 33303
rect 21005 33065 21039 33099
rect 22661 33065 22695 33099
rect 25145 33065 25179 33099
rect 26157 33065 26191 33099
rect 28457 33065 28491 33099
rect 23029 32997 23063 33031
rect 25421 32997 25455 33031
rect 27721 32997 27755 33031
rect 29837 32997 29871 33031
rect 1409 32929 1443 32963
rect 16957 32929 16991 32963
rect 22937 32929 22971 32963
rect 25145 32929 25179 32963
rect 28917 32929 28951 32963
rect 30757 32929 30791 32963
rect 31769 32929 31803 32963
rect 35265 32929 35299 32963
rect 19257 32861 19291 32895
rect 20361 32861 20395 32895
rect 20545 32861 20579 32895
rect 21281 32861 21315 32895
rect 21370 32858 21404 32892
rect 21465 32861 21499 32895
rect 21649 32861 21683 32895
rect 22845 32861 22879 32895
rect 23121 32861 23155 32895
rect 23305 32861 23339 32895
rect 25237 32861 25271 32895
rect 25973 32861 26007 32895
rect 27997 32861 28031 32895
rect 28641 32861 28675 32895
rect 28733 32861 28767 32895
rect 29009 32861 29043 32895
rect 30481 32861 30515 32895
rect 30573 32861 30607 32895
rect 30849 32861 30883 32895
rect 31493 32861 31527 32895
rect 31677 32861 31711 32895
rect 32229 32861 32263 32895
rect 32413 32861 32447 32895
rect 35081 32861 35115 32895
rect 35357 32861 35391 32895
rect 35817 32861 35851 32895
rect 46305 32861 46339 32895
rect 1593 32793 1627 32827
rect 3249 32793 3283 32827
rect 17233 32793 17267 32827
rect 19349 32793 19383 32827
rect 24961 32793 24995 32827
rect 27721 32793 27755 32827
rect 29653 32793 29687 32827
rect 30297 32793 30331 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 18705 32725 18739 32759
rect 20453 32725 20487 32759
rect 27905 32725 27939 32759
rect 31309 32725 31343 32759
rect 32321 32725 32355 32759
rect 34897 32725 34931 32759
rect 35909 32725 35943 32759
rect 18521 32521 18555 32555
rect 22293 32521 22327 32555
rect 23213 32521 23247 32555
rect 26249 32521 26283 32555
rect 28089 32521 28123 32555
rect 33793 32521 33827 32555
rect 47685 32521 47719 32555
rect 2145 32453 2179 32487
rect 22201 32453 22235 32487
rect 24593 32453 24627 32487
rect 27997 32453 28031 32487
rect 28917 32453 28951 32487
rect 30113 32453 30147 32487
rect 35081 32453 35115 32487
rect 17785 32385 17819 32419
rect 17969 32385 18003 32419
rect 18337 32385 18371 32419
rect 22845 32385 22879 32419
rect 23029 32385 23063 32419
rect 23857 32385 23891 32419
rect 24869 32385 24903 32419
rect 25973 32385 26007 32419
rect 27261 32385 27295 32419
rect 28733 32385 28767 32419
rect 32413 32385 32447 32419
rect 32781 32385 32815 32419
rect 33609 32385 33643 32419
rect 34805 32385 34839 32419
rect 47041 32385 47075 32419
rect 47593 32385 47627 32419
rect 1961 32317 1995 32351
rect 3801 32317 3835 32351
rect 18061 32317 18095 32351
rect 18153 32317 18187 32351
rect 24133 32317 24167 32351
rect 24777 32317 24811 32351
rect 29837 32317 29871 32351
rect 31585 32317 31619 32351
rect 33425 32317 33459 32351
rect 25053 32249 25087 32283
rect 32965 32249 32999 32283
rect 23673 32181 23707 32215
rect 24041 32181 24075 32215
rect 24777 32181 24811 32215
rect 27353 32181 27387 32215
rect 32505 32181 32539 32215
rect 36553 32181 36587 32215
rect 46857 32181 46891 32215
rect 1409 31977 1443 32011
rect 22201 31977 22235 32011
rect 23397 31977 23431 32011
rect 26525 31977 26559 32011
rect 31493 31977 31527 32011
rect 33793 31977 33827 32011
rect 34713 31977 34747 32011
rect 35173 31977 35207 32011
rect 35725 31977 35759 32011
rect 47685 31977 47719 32011
rect 23581 31909 23615 31943
rect 25605 31909 25639 31943
rect 25145 31841 25179 31875
rect 27261 31841 27295 31875
rect 29837 31841 29871 31875
rect 31217 31841 31251 31875
rect 32505 31841 32539 31875
rect 32597 31841 32631 31875
rect 34805 31841 34839 31875
rect 36185 31841 36219 31875
rect 1593 31773 1627 31807
rect 2329 31773 2363 31807
rect 2973 31773 3007 31807
rect 20545 31773 20579 31807
rect 22201 31773 22235 31807
rect 22385 31773 22419 31807
rect 23029 31773 23063 31807
rect 23305 31773 23339 31807
rect 25237 31773 25271 31807
rect 26341 31773 26375 31807
rect 31125 31773 31159 31807
rect 32229 31773 32263 31807
rect 32413 31773 32447 31807
rect 32781 31773 32815 31807
rect 33609 31773 33643 31807
rect 34989 31773 35023 31807
rect 35909 31773 35943 31807
rect 36001 31773 36035 31807
rect 36277 31773 36311 31807
rect 20913 31705 20947 31739
rect 27537 31705 27571 31739
rect 29653 31705 29687 31739
rect 33425 31705 33459 31739
rect 34713 31705 34747 31739
rect 3065 31637 3099 31671
rect 29009 31637 29043 31671
rect 32965 31637 32999 31671
rect 22661 31433 22695 31467
rect 27905 31433 27939 31467
rect 31217 31433 31251 31467
rect 34345 31433 34379 31467
rect 35173 31433 35207 31467
rect 35725 31433 35759 31467
rect 2237 31365 2271 31399
rect 21833 31365 21867 31399
rect 32873 31365 32907 31399
rect 2053 31297 2087 31331
rect 17325 31297 17359 31331
rect 19533 31297 19567 31331
rect 20269 31297 20303 31331
rect 20453 31297 20487 31331
rect 20913 31297 20947 31331
rect 21097 31297 21131 31331
rect 21281 31297 21315 31331
rect 22017 31297 22051 31331
rect 22109 31297 22143 31331
rect 22569 31297 22603 31331
rect 23949 31297 23983 31331
rect 25421 31297 25455 31331
rect 27268 31297 27302 31331
rect 27409 31297 27443 31331
rect 27537 31297 27571 31331
rect 27629 31297 27663 31331
rect 27767 31297 27801 31331
rect 28365 31297 28399 31331
rect 29193 31297 29227 31331
rect 31125 31297 31159 31331
rect 32597 31297 32631 31331
rect 34805 31297 34839 31331
rect 34897 31297 34931 31331
rect 35633 31297 35667 31331
rect 35817 31297 35851 31331
rect 2789 31229 2823 31263
rect 17601 31229 17635 31263
rect 25513 31229 25547 31263
rect 25697 31229 25731 31263
rect 29377 31161 29411 31195
rect 19073 31093 19107 31127
rect 19625 31093 19659 31127
rect 20361 31093 20395 31127
rect 21833 31093 21867 31127
rect 24041 31093 24075 31127
rect 25053 31093 25087 31127
rect 28549 31093 28583 31127
rect 34805 31093 34839 31127
rect 18521 30889 18555 30923
rect 19257 30889 19291 30923
rect 21281 30889 21315 30923
rect 28365 30889 28399 30923
rect 33517 30889 33551 30923
rect 19625 30821 19659 30855
rect 19717 30753 19751 30787
rect 22293 30753 22327 30787
rect 18429 30685 18463 30719
rect 19441 30685 19475 30719
rect 20453 30685 20487 30719
rect 20545 30685 20579 30719
rect 20729 30685 20763 30719
rect 20821 30685 20855 30719
rect 21281 30685 21315 30719
rect 21373 30685 21407 30719
rect 22569 30685 22603 30719
rect 24593 30685 24627 30719
rect 28181 30685 28215 30719
rect 30021 30685 30055 30719
rect 32321 30685 32355 30719
rect 32413 30685 32447 30719
rect 32597 30685 32631 30719
rect 32689 30685 32723 30719
rect 33425 30685 33459 30719
rect 20269 30617 20303 30651
rect 23673 30617 23707 30651
rect 25973 30617 26007 30651
rect 30757 30617 30791 30651
rect 30941 30617 30975 30651
rect 21649 30549 21683 30583
rect 23765 30549 23799 30583
rect 24409 30549 24443 30583
rect 27261 30549 27295 30583
rect 30113 30549 30147 30583
rect 32137 30549 32171 30583
rect 19625 30345 19659 30379
rect 25881 30277 25915 30311
rect 30389 30277 30423 30311
rect 20545 30209 20579 30243
rect 20729 30209 20763 30243
rect 20821 30209 20855 30243
rect 21097 30209 21131 30243
rect 21833 30209 21867 30243
rect 22569 30209 22603 30243
rect 25789 30209 25823 30243
rect 26985 30209 27019 30243
rect 27261 30209 27295 30243
rect 28641 30209 28675 30243
rect 29377 30209 29411 30243
rect 30205 30209 30239 30243
rect 33517 30209 33551 30243
rect 17877 30141 17911 30175
rect 18153 30141 18187 30175
rect 20913 30141 20947 30175
rect 23213 30141 23247 30175
rect 23489 30141 23523 30175
rect 24961 30141 24995 30175
rect 26065 30141 26099 30175
rect 21281 30073 21315 30107
rect 25421 30073 25455 30107
rect 21925 30005 21959 30039
rect 22661 30005 22695 30039
rect 28825 30005 28859 30039
rect 29561 30005 29595 30039
rect 33609 30005 33643 30039
rect 20729 29801 20763 29835
rect 26341 29801 26375 29835
rect 28365 29801 28399 29835
rect 34161 29801 34195 29835
rect 20821 29733 20855 29767
rect 28549 29733 28583 29767
rect 20913 29665 20947 29699
rect 24501 29665 24535 29699
rect 47593 29665 47627 29699
rect 20637 29597 20671 29631
rect 21005 29597 21039 29631
rect 24409 29597 24443 29631
rect 24593 29597 24627 29631
rect 25145 29597 25179 29631
rect 26249 29597 26283 29631
rect 26433 29597 26467 29631
rect 29561 29597 29595 29631
rect 29654 29597 29688 29631
rect 30067 29597 30101 29631
rect 30757 29597 30791 29631
rect 30941 29597 30975 29631
rect 32413 29597 32447 29631
rect 47317 29597 47351 29631
rect 28181 29529 28215 29563
rect 29837 29529 29871 29563
rect 29929 29529 29963 29563
rect 32689 29529 32723 29563
rect 25237 29461 25271 29495
rect 28381 29461 28415 29495
rect 30205 29461 30239 29495
rect 24409 29257 24443 29291
rect 26157 29257 26191 29291
rect 29193 29257 29227 29291
rect 20361 29189 20395 29223
rect 21833 29189 21867 29223
rect 22753 29189 22787 29223
rect 30113 29189 30147 29223
rect 33149 29189 33183 29223
rect 17049 29121 17083 29155
rect 20085 29121 20119 29155
rect 20269 29121 20303 29155
rect 20453 29121 20487 29155
rect 22017 29121 22051 29155
rect 23581 29121 23615 29155
rect 24317 29121 24351 29155
rect 25421 29121 25455 29155
rect 26065 29121 26099 29155
rect 27169 29121 27203 29155
rect 27261 29121 27295 29155
rect 27445 29121 27479 29155
rect 27537 29121 27571 29155
rect 28825 29121 28859 29155
rect 29837 29121 29871 29155
rect 32413 29121 32447 29155
rect 32597 29121 32631 29155
rect 32965 29121 32999 29155
rect 14289 29053 14323 29087
rect 14473 29053 14507 29087
rect 14749 29053 14783 29087
rect 17325 29053 17359 29087
rect 22201 29053 22235 29087
rect 28733 29053 28767 29087
rect 31585 29053 31619 29087
rect 32689 29053 32723 29087
rect 32781 29053 32815 29087
rect 22937 28985 22971 29019
rect 23765 28985 23799 29019
rect 25605 28985 25639 29019
rect 18797 28917 18831 28951
rect 20637 28917 20671 28951
rect 26985 28917 27019 28951
rect 14749 28713 14783 28747
rect 18429 28713 18463 28747
rect 21281 28713 21315 28747
rect 28549 28713 28583 28747
rect 31309 28713 31343 28747
rect 26801 28645 26835 28679
rect 15853 28577 15887 28611
rect 17969 28577 18003 28611
rect 20177 28577 20211 28611
rect 21373 28577 21407 28611
rect 24869 28577 24903 28611
rect 25053 28577 25087 28611
rect 27629 28577 27663 28611
rect 14657 28509 14691 28543
rect 15393 28509 15427 28543
rect 17693 28509 17727 28543
rect 17877 28509 17911 28543
rect 18061 28509 18095 28543
rect 18245 28509 18279 28543
rect 20085 28509 20119 28543
rect 21097 28509 21131 28543
rect 22017 28509 22051 28543
rect 22201 28509 22235 28543
rect 22293 28509 22327 28543
rect 23397 28509 23431 28543
rect 23673 28509 23707 28543
rect 24777 28509 24811 28543
rect 25697 28509 25731 28543
rect 25789 28509 25823 28543
rect 26617 28509 26651 28543
rect 26893 28509 26927 28543
rect 28365 28509 28399 28543
rect 31217 28509 31251 28543
rect 15577 28441 15611 28475
rect 25973 28441 26007 28475
rect 27445 28441 27479 28475
rect 28181 28441 28215 28475
rect 20453 28373 20487 28407
rect 20913 28373 20947 28407
rect 21833 28373 21867 28407
rect 23213 28373 23247 28407
rect 23581 28373 23615 28407
rect 24409 28373 24443 28407
rect 26433 28373 26467 28407
rect 15577 28169 15611 28203
rect 27169 28169 27203 28203
rect 28089 28169 28123 28203
rect 29009 28169 29043 28203
rect 31217 28169 31251 28203
rect 19257 28101 19291 28135
rect 22937 28101 22971 28135
rect 30297 28101 30331 28135
rect 30481 28101 30515 28135
rect 31033 28101 31067 28135
rect 32207 28101 32241 28135
rect 15485 28033 15519 28067
rect 18981 28033 19015 28067
rect 21833 28033 21867 28067
rect 22661 28033 22695 28067
rect 23949 28033 23983 28067
rect 24133 28033 24167 28067
rect 26249 28033 26283 28067
rect 26985 28033 27019 28067
rect 27261 28033 27295 28067
rect 27721 28033 27755 28067
rect 28549 28033 28583 28067
rect 28825 28033 28859 28067
rect 29653 28033 29687 28067
rect 30573 28033 30607 28067
rect 31309 28033 31343 28067
rect 32505 28033 32539 28067
rect 46765 28033 46799 28067
rect 12265 27965 12299 27999
rect 12541 27965 12575 27999
rect 14013 27965 14047 27999
rect 16681 27965 16715 27999
rect 16865 27965 16899 27999
rect 17141 27965 17175 27999
rect 20729 27965 20763 27999
rect 21925 27965 21959 27999
rect 27813 27965 27847 27999
rect 28641 27965 28675 27999
rect 29469 27965 29503 27999
rect 32137 27965 32171 27999
rect 32321 27965 32355 27999
rect 22201 27897 22235 27931
rect 22753 27897 22787 27931
rect 24317 27897 24351 27931
rect 26985 27897 27019 27931
rect 30297 27897 30331 27931
rect 21833 27829 21867 27863
rect 22845 27829 22879 27863
rect 26341 27829 26375 27863
rect 27905 27829 27939 27863
rect 28825 27829 28859 27863
rect 29837 27829 29871 27863
rect 31033 27829 31067 27863
rect 32413 27829 32447 27863
rect 46857 27829 46891 27863
rect 47777 27829 47811 27863
rect 11529 27625 11563 27659
rect 12541 27625 12575 27659
rect 17233 27625 17267 27659
rect 25776 27625 25810 27659
rect 27261 27625 27295 27659
rect 29929 27625 29963 27659
rect 31290 27625 31324 27659
rect 14197 27557 14231 27591
rect 18245 27557 18279 27591
rect 19349 27557 19383 27591
rect 21925 27557 21959 27591
rect 27905 27557 27939 27591
rect 12357 27489 12391 27523
rect 13185 27489 13219 27523
rect 16497 27489 16531 27523
rect 22017 27489 22051 27523
rect 27997 27489 28031 27523
rect 29837 27489 29871 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 11437 27421 11471 27455
rect 12265 27421 12299 27455
rect 13093 27421 13127 27455
rect 13277 27421 13311 27455
rect 14105 27421 14139 27455
rect 14841 27421 14875 27455
rect 17141 27421 17175 27455
rect 18153 27421 18187 27455
rect 19257 27421 19291 27455
rect 20453 27421 20487 27455
rect 20821 27421 20855 27455
rect 21796 27421 21830 27455
rect 25513 27421 25547 27455
rect 27721 27421 27755 27455
rect 27813 27421 27847 27455
rect 28641 27421 28675 27455
rect 29009 27421 29043 27455
rect 29561 27421 29595 27455
rect 31033 27421 31067 27455
rect 15025 27353 15059 27387
rect 20637 27353 20671 27387
rect 21649 27353 21683 27387
rect 28825 27353 28859 27387
rect 22293 27285 22327 27319
rect 30113 27285 30147 27319
rect 32781 27285 32815 27319
rect 15025 27081 15059 27115
rect 26249 27081 26283 27115
rect 22017 27013 22051 27047
rect 23489 27013 23523 27047
rect 24961 27013 24995 27047
rect 29377 27013 29411 27047
rect 30113 27013 30147 27047
rect 32229 27013 32263 27047
rect 10333 26945 10367 26979
rect 12541 26945 12575 26979
rect 12725 26945 12759 26979
rect 14933 26945 14967 26979
rect 20821 26945 20855 26979
rect 21005 26945 21039 26979
rect 21281 26945 21315 26979
rect 21925 26945 21959 26979
rect 22201 26945 22235 26979
rect 22477 26945 22511 26979
rect 23305 26945 23339 26979
rect 24777 26945 24811 26979
rect 26065 26945 26099 26979
rect 28641 26945 28675 26979
rect 28829 26943 28863 26977
rect 28917 26945 28951 26979
rect 29055 26945 29089 26979
rect 29193 26945 29227 26979
rect 32137 26945 32171 26979
rect 7849 26877 7883 26911
rect 8033 26877 8067 26911
rect 8309 26877 8343 26911
rect 10425 26877 10459 26911
rect 20913 26877 20947 26911
rect 22109 26877 22143 26911
rect 29837 26877 29871 26911
rect 10701 26741 10735 26775
rect 12541 26741 12575 26775
rect 20545 26741 20579 26775
rect 21097 26741 21131 26775
rect 22311 26741 22345 26775
rect 31585 26741 31619 26775
rect 8125 26537 8159 26571
rect 12541 26537 12575 26571
rect 19441 26537 19475 26571
rect 22017 26537 22051 26571
rect 31125 26537 31159 26571
rect 14289 26469 14323 26503
rect 26525 26469 26559 26503
rect 9689 26401 9723 26435
rect 11161 26401 11195 26435
rect 12357 26401 12391 26435
rect 13001 26401 13035 26435
rect 23489 26401 23523 26435
rect 7389 26333 7423 26367
rect 8033 26333 8067 26367
rect 9413 26333 9447 26367
rect 12173 26333 12207 26367
rect 12265 26333 12299 26367
rect 12541 26333 12575 26367
rect 13369 26333 13403 26367
rect 13553 26333 13587 26367
rect 14657 26333 14691 26367
rect 19257 26333 19291 26367
rect 21649 26333 21683 26367
rect 22661 26333 22695 26367
rect 22937 26333 22971 26367
rect 23397 26333 23431 26367
rect 23581 26333 23615 26367
rect 26525 26333 26559 26367
rect 26709 26333 26743 26367
rect 26801 26333 26835 26367
rect 27261 26333 27295 26367
rect 27445 26333 27479 26367
rect 31033 26333 31067 26367
rect 13185 26265 13219 26299
rect 14841 26265 14875 26299
rect 21833 26265 21867 26299
rect 22477 26265 22511 26299
rect 27353 26265 27387 26299
rect 7481 26197 7515 26231
rect 13277 26197 13311 26231
rect 14473 26197 14507 26231
rect 14565 26197 14599 26231
rect 22845 26197 22879 26231
rect 10517 25993 10551 26027
rect 15669 25993 15703 26027
rect 24225 25993 24259 26027
rect 27537 25993 27571 26027
rect 8217 25925 8251 25959
rect 22753 25925 22787 25959
rect 26065 25925 26099 25959
rect 26249 25925 26283 25959
rect 27169 25925 27203 25959
rect 10425 25857 10459 25891
rect 17141 25857 17175 25891
rect 17325 25857 17359 25891
rect 23029 25857 23063 25891
rect 23118 25857 23152 25891
rect 23218 25857 23252 25891
rect 23397 25857 23431 25891
rect 24041 25857 24075 25891
rect 24317 25857 24351 25891
rect 26985 25857 27019 25891
rect 27261 25857 27295 25891
rect 27353 25857 27387 25891
rect 28917 25857 28951 25891
rect 8033 25789 8067 25823
rect 8493 25789 8527 25823
rect 11713 25789 11747 25823
rect 11989 25789 12023 25823
rect 13921 25789 13955 25823
rect 14197 25789 14231 25823
rect 19533 25789 19567 25823
rect 19809 25789 19843 25823
rect 13461 25653 13495 25687
rect 17141 25653 17175 25687
rect 21281 25653 21315 25687
rect 23857 25653 23891 25687
rect 26433 25653 26467 25687
rect 29009 25653 29043 25687
rect 47777 25653 47811 25687
rect 9505 25449 9539 25483
rect 11621 25449 11655 25483
rect 13185 25449 13219 25483
rect 14105 25449 14139 25483
rect 14473 25449 14507 25483
rect 15117 25449 15151 25483
rect 16129 25449 16163 25483
rect 20177 25449 20211 25483
rect 22661 25449 22695 25483
rect 27629 25449 27663 25483
rect 27905 25449 27939 25483
rect 28733 25381 28767 25415
rect 14565 25313 14599 25347
rect 17141 25313 17175 25347
rect 22017 25313 22051 25347
rect 22502 25313 22536 25347
rect 30021 25313 30055 25347
rect 46305 25313 46339 25347
rect 1409 25245 1443 25279
rect 9505 25245 9539 25279
rect 10057 25245 10091 25279
rect 10241 25245 10275 25279
rect 11621 25245 11655 25279
rect 13093 25245 13127 25279
rect 14289 25245 14323 25279
rect 15025 25245 15059 25279
rect 16129 25245 16163 25279
rect 16405 25245 16439 25279
rect 16865 25245 16899 25279
rect 19257 25245 19291 25279
rect 20085 25245 20119 25279
rect 20729 25245 20763 25279
rect 21557 25245 21591 25279
rect 22293 25245 22327 25279
rect 25789 25245 25823 25279
rect 26617 25245 26651 25279
rect 27629 25245 27663 25279
rect 27721 25245 27755 25279
rect 28641 25245 28675 25279
rect 28825 25245 28859 25279
rect 28917 25245 28951 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 29837 25245 29871 25279
rect 30113 25245 30147 25279
rect 30573 25245 30607 25279
rect 48145 25245 48179 25279
rect 1685 25177 1719 25211
rect 22385 25177 22419 25211
rect 26801 25177 26835 25211
rect 27445 25177 27479 25211
rect 46489 25177 46523 25211
rect 10149 25109 10183 25143
rect 16313 25109 16347 25143
rect 18613 25109 18647 25143
rect 19349 25109 19383 25143
rect 20821 25109 20855 25143
rect 21373 25109 21407 25143
rect 25605 25109 25639 25143
rect 26985 25109 27019 25143
rect 28457 25109 28491 25143
rect 30665 25109 30699 25143
rect 14565 24905 14599 24939
rect 15853 24905 15887 24939
rect 15945 24905 15979 24939
rect 16865 24905 16899 24939
rect 22109 24905 22143 24939
rect 30941 24905 30975 24939
rect 15761 24837 15795 24871
rect 8309 24769 8343 24803
rect 13185 24769 13219 24803
rect 13829 24769 13863 24803
rect 14013 24769 14047 24803
rect 14473 24769 14507 24803
rect 15577 24769 15611 24803
rect 16681 24769 16715 24803
rect 18245 24769 18279 24803
rect 18337 24769 18371 24803
rect 22477 24769 22511 24803
rect 22569 24769 22603 24803
rect 27629 24769 27663 24803
rect 46857 24769 46891 24803
rect 47593 24769 47627 24803
rect 47685 24769 47719 24803
rect 8401 24701 8435 24735
rect 8861 24701 8895 24735
rect 9137 24701 9171 24735
rect 18981 24701 19015 24735
rect 19165 24701 19199 24735
rect 20821 24701 20855 24735
rect 22753 24701 22787 24735
rect 23305 24701 23339 24735
rect 23581 24701 23615 24735
rect 25053 24701 25087 24735
rect 27721 24701 27755 24735
rect 29193 24701 29227 24735
rect 29469 24701 29503 24735
rect 13369 24633 13403 24667
rect 16129 24633 16163 24667
rect 10609 24565 10643 24599
rect 13921 24565 13955 24599
rect 23121 24565 23155 24599
rect 27905 24565 27939 24599
rect 46949 24565 46983 24599
rect 9965 24361 9999 24395
rect 18521 24361 18555 24395
rect 19809 24361 19843 24395
rect 22109 24361 22143 24395
rect 26433 24361 26467 24395
rect 27537 24361 27571 24395
rect 28549 24361 28583 24395
rect 28917 24361 28951 24395
rect 29929 24361 29963 24395
rect 16037 24225 16071 24259
rect 17049 24225 17083 24259
rect 20361 24225 20395 24259
rect 24685 24225 24719 24259
rect 24961 24225 24995 24259
rect 27997 24225 28031 24259
rect 29009 24225 29043 24259
rect 30021 24225 30055 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 9873 24157 9907 24191
rect 12449 24157 12483 24191
rect 13185 24157 13219 24191
rect 15853 24157 15887 24191
rect 16313 24157 16347 24191
rect 16773 24157 16807 24191
rect 19625 24157 19659 24191
rect 27721 24157 27755 24191
rect 27813 24157 27847 24191
rect 28089 24157 28123 24191
rect 28733 24157 28767 24191
rect 29745 24157 29779 24191
rect 46305 24157 46339 24191
rect 13369 24089 13403 24123
rect 20637 24089 20671 24123
rect 12541 24021 12575 24055
rect 16221 24021 16255 24055
rect 29561 24021 29595 24055
rect 1593 23817 1627 23851
rect 12817 23817 12851 23851
rect 14565 23817 14599 23851
rect 15669 23817 15703 23851
rect 15853 23817 15887 23851
rect 16865 23817 16899 23851
rect 18337 23817 18371 23851
rect 24409 23817 24443 23851
rect 25697 23817 25731 23851
rect 28733 23817 28767 23851
rect 9413 23749 9447 23783
rect 11529 23749 11563 23783
rect 11745 23749 11779 23783
rect 13645 23749 13679 23783
rect 14657 23749 14691 23783
rect 15301 23749 15335 23783
rect 26341 23749 26375 23783
rect 45385 23749 45419 23783
rect 1409 23681 1443 23715
rect 8493 23681 8527 23715
rect 9597 23681 9631 23715
rect 9689 23681 9723 23715
rect 10149 23681 10183 23715
rect 12633 23681 12667 23715
rect 13277 23681 13311 23715
rect 13461 23681 13495 23715
rect 14473 23681 14507 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 16681 23681 16715 23715
rect 18245 23681 18279 23715
rect 18889 23681 18923 23715
rect 24317 23681 24351 23715
rect 25605 23681 25639 23715
rect 26249 23681 26283 23715
rect 26985 23681 27019 23715
rect 47777 23681 47811 23715
rect 12449 23613 12483 23647
rect 14289 23613 14323 23647
rect 27261 23613 27295 23647
rect 45201 23613 45235 23647
rect 46765 23613 46799 23647
rect 9413 23545 9447 23579
rect 11897 23545 11931 23579
rect 8309 23477 8343 23511
rect 10241 23477 10275 23511
rect 11713 23477 11747 23511
rect 14841 23477 14875 23511
rect 18981 23477 19015 23511
rect 9505 23273 9539 23307
rect 10241 23273 10275 23307
rect 10425 23273 10459 23307
rect 11897 23273 11931 23307
rect 15485 23273 15519 23307
rect 19441 23273 19475 23307
rect 22017 23205 22051 23239
rect 13277 23137 13311 23171
rect 27353 23137 27387 23171
rect 46305 23137 46339 23171
rect 46857 23137 46891 23171
rect 9134 23069 9168 23103
rect 9597 23069 9631 23103
rect 13185 23069 13219 23103
rect 14289 23069 14323 23103
rect 14841 23069 14875 23103
rect 15669 23069 15703 23103
rect 15945 23069 15979 23103
rect 19257 23069 19291 23103
rect 22293 23069 22327 23103
rect 22753 23069 22787 23103
rect 27169 23069 27203 23103
rect 44465 23069 44499 23103
rect 45385 23069 45419 23103
rect 45569 23069 45603 23103
rect 10057 23001 10091 23035
rect 10977 23001 11011 23035
rect 11161 23001 11195 23035
rect 11805 23001 11839 23035
rect 15853 23001 15887 23035
rect 22017 23001 22051 23035
rect 29009 23001 29043 23035
rect 46489 23001 46523 23035
rect 8953 22933 8987 22967
rect 9137 22933 9171 22967
rect 10257 22933 10291 22967
rect 13553 22933 13587 22967
rect 14289 22933 14323 22967
rect 14933 22933 14967 22967
rect 22201 22933 22235 22967
rect 22845 22933 22879 22967
rect 44281 22933 44315 22967
rect 45477 22933 45511 22967
rect 9781 22729 9815 22763
rect 10451 22729 10485 22763
rect 11989 22729 12023 22763
rect 15117 22729 15151 22763
rect 23949 22729 23983 22763
rect 47685 22729 47719 22763
rect 8309 22661 8343 22695
rect 10241 22661 10275 22695
rect 11621 22661 11655 22695
rect 11837 22661 11871 22695
rect 13645 22661 13679 22695
rect 21189 22661 21223 22695
rect 22477 22661 22511 22695
rect 26433 22661 26467 22695
rect 12633 22593 12667 22627
rect 15853 22593 15887 22627
rect 18521 22593 18555 22627
rect 19349 22593 19383 22627
rect 21097 22593 21131 22627
rect 21281 22593 21315 22627
rect 24593 22593 24627 22627
rect 29469 22593 29503 22627
rect 44649 22593 44683 22627
rect 44925 22593 44959 22627
rect 46489 22593 46523 22627
rect 47593 22593 47627 22627
rect 8033 22525 8067 22559
rect 13369 22525 13403 22559
rect 22201 22525 22235 22559
rect 24777 22525 24811 22559
rect 27629 22525 27663 22559
rect 27813 22525 27847 22559
rect 46213 22525 46247 22559
rect 10609 22457 10643 22491
rect 45109 22457 45143 22491
rect 10425 22389 10459 22423
rect 11805 22389 11839 22423
rect 12817 22389 12851 22423
rect 15669 22389 15703 22423
rect 18705 22389 18739 22423
rect 19441 22389 19475 22423
rect 14289 22185 14323 22219
rect 22201 22185 22235 22219
rect 22845 22185 22879 22219
rect 15209 22049 15243 22083
rect 16957 22049 16991 22083
rect 17969 22049 18003 22083
rect 18429 22049 18463 22083
rect 19533 22049 19567 22083
rect 21005 22049 21039 22083
rect 24961 22049 24995 22083
rect 29745 22049 29779 22083
rect 44373 22049 44407 22083
rect 46305 22049 46339 22083
rect 46949 22049 46983 22083
rect 9873 21981 9907 22015
rect 10149 21981 10183 22015
rect 10609 21981 10643 22015
rect 14105 21981 14139 22015
rect 18061 21981 18095 22015
rect 19257 21981 19291 22015
rect 22845 21981 22879 22015
rect 24869 21981 24903 22015
rect 25513 21981 25547 22015
rect 27353 21981 27387 22015
rect 28733 21981 28767 22015
rect 29561 21981 29595 22015
rect 43453 21981 43487 22015
rect 43637 21981 43671 22015
rect 45293 21981 45327 22015
rect 45569 21981 45603 22015
rect 10885 21913 10919 21947
rect 15485 21913 15519 21947
rect 22017 21913 22051 21947
rect 25697 21913 25731 21947
rect 27905 21913 27939 21947
rect 31401 21913 31435 21947
rect 45661 21913 45695 21947
rect 46489 21913 46523 21947
rect 9689 21845 9723 21879
rect 10057 21845 10091 21879
rect 12357 21845 12391 21879
rect 22217 21845 22251 21879
rect 22385 21845 22419 21879
rect 27997 21845 28031 21879
rect 28825 21845 28859 21879
rect 10885 21641 10919 21675
rect 16773 21641 16807 21675
rect 22477 21641 22511 21675
rect 22569 21641 22603 21675
rect 26249 21641 26283 21675
rect 29929 21641 29963 21675
rect 44005 21641 44039 21675
rect 44649 21641 44683 21675
rect 9781 21573 9815 21607
rect 22385 21573 22419 21607
rect 47961 21573 47995 21607
rect 10793 21505 10827 21539
rect 11897 21505 11931 21539
rect 14381 21505 14415 21539
rect 15301 21505 15335 21539
rect 16681 21505 16715 21539
rect 17325 21505 17359 21539
rect 18337 21505 18371 21539
rect 19533 21505 19567 21539
rect 20269 21505 20303 21539
rect 21097 21505 21131 21539
rect 23397 21505 23431 21539
rect 25513 21505 25547 21539
rect 26157 21505 26191 21539
rect 27537 21505 27571 21539
rect 29009 21505 29043 21539
rect 29377 21505 29411 21539
rect 29837 21505 29871 21539
rect 39129 21505 39163 21539
rect 44465 21505 44499 21539
rect 45201 21505 45235 21539
rect 45661 21505 45695 21539
rect 15393 21437 15427 21471
rect 15669 21437 15703 21471
rect 20361 21437 20395 21471
rect 22753 21437 22787 21471
rect 23213 21437 23247 21471
rect 28273 21437 28307 21471
rect 39313 21437 39347 21471
rect 39589 21437 39623 21471
rect 44373 21437 44407 21471
rect 10057 21369 10091 21403
rect 12081 21369 12115 21403
rect 18521 21369 18555 21403
rect 22201 21369 22235 21403
rect 48145 21369 48179 21403
rect 10241 21301 10275 21335
rect 14473 21301 14507 21335
rect 17417 21301 17451 21335
rect 19533 21301 19567 21335
rect 20637 21301 20671 21335
rect 21189 21301 21223 21335
rect 23581 21301 23615 21335
rect 25605 21301 25639 21335
rect 46673 21301 46707 21335
rect 45753 21097 45787 21131
rect 11253 21029 11287 21063
rect 22385 21029 22419 21063
rect 8125 20961 8159 20995
rect 8401 20961 8435 20995
rect 9229 20961 9263 20995
rect 14105 20961 14139 20995
rect 14289 20961 14323 20995
rect 15485 20961 15519 20995
rect 16865 20961 16899 20995
rect 17049 20961 17083 20995
rect 20177 20961 20211 20995
rect 20453 20961 20487 20995
rect 25789 20961 25823 20995
rect 27445 20961 27479 20995
rect 29561 20961 29595 20995
rect 30481 20961 30515 20995
rect 48145 20961 48179 20995
rect 8033 20893 8067 20927
rect 8953 20893 8987 20927
rect 11437 20893 11471 20927
rect 19257 20893 19291 20927
rect 22661 20893 22695 20927
rect 23121 20893 23155 20927
rect 24409 20893 24443 20927
rect 25605 20893 25639 20927
rect 27905 20893 27939 20927
rect 45385 20893 45419 20927
rect 46305 20893 46339 20927
rect 18705 20825 18739 20859
rect 22385 20825 22419 20859
rect 28733 20825 28767 20859
rect 29745 20825 29779 20859
rect 45569 20825 45603 20859
rect 46489 20825 46523 20859
rect 10701 20757 10735 20791
rect 19349 20757 19383 20791
rect 21925 20757 21959 20791
rect 22569 20757 22603 20791
rect 23305 20757 23339 20791
rect 24501 20757 24535 20791
rect 43729 20553 43763 20587
rect 47685 20553 47719 20587
rect 9965 20485 9999 20519
rect 15669 20485 15703 20519
rect 18429 20485 18463 20519
rect 27905 20485 27939 20519
rect 45385 20485 45419 20519
rect 7573 20417 7607 20451
rect 9873 20417 9907 20451
rect 10701 20417 10735 20451
rect 11805 20417 11839 20451
rect 12633 20417 12667 20451
rect 15301 20417 15335 20451
rect 16865 20417 16899 20451
rect 18245 20417 18279 20451
rect 20545 20417 20579 20451
rect 22569 20417 22603 20451
rect 22753 20417 22787 20451
rect 23213 20417 23247 20451
rect 26065 20417 26099 20451
rect 27077 20417 27111 20451
rect 43821 20417 43855 20451
rect 44189 20417 44223 20451
rect 47593 20417 47627 20451
rect 45201 20383 45235 20417
rect 7757 20349 7791 20383
rect 8033 20349 8067 20383
rect 12817 20349 12851 20383
rect 14381 20349 14415 20383
rect 17049 20349 17083 20383
rect 18705 20349 18739 20383
rect 22661 20349 22695 20383
rect 23489 20349 23523 20383
rect 24961 20349 24995 20383
rect 27721 20349 27755 20383
rect 28181 20349 28215 20383
rect 44649 20349 44683 20383
rect 46673 20349 46707 20383
rect 10517 20281 10551 20315
rect 11989 20213 12023 20247
rect 20637 20213 20671 20247
rect 26157 20213 26191 20247
rect 27169 20213 27203 20247
rect 7941 20009 7975 20043
rect 8953 20009 8987 20043
rect 12817 20009 12851 20043
rect 25145 19941 25179 19975
rect 45385 19941 45419 19975
rect 16405 19873 16439 19907
rect 19533 19873 19567 19907
rect 19717 19873 19751 19907
rect 22937 19873 22971 19907
rect 23213 19873 23247 19907
rect 40785 19873 40819 19907
rect 43637 19873 43671 19907
rect 45477 19873 45511 19907
rect 46489 19873 46523 19907
rect 2053 19805 2087 19839
rect 7849 19805 7883 19839
rect 9137 19805 9171 19839
rect 12725 19805 12759 19839
rect 15209 19805 15243 19839
rect 16129 19805 16163 19839
rect 17417 19805 17451 19839
rect 22017 19805 22051 19839
rect 22845 19805 22879 19839
rect 23673 19805 23707 19839
rect 24961 19805 24995 19839
rect 25881 19805 25915 19839
rect 27169 19805 27203 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 43821 19805 43855 19839
rect 46305 19805 46339 19839
rect 18245 19737 18279 19771
rect 21373 19737 21407 19771
rect 26525 19737 26559 19771
rect 27997 19737 28031 19771
rect 29009 19737 29043 19771
rect 30021 19737 30055 19771
rect 40969 19737 41003 19771
rect 42625 19737 42659 19771
rect 45017 19737 45051 19771
rect 48145 19737 48179 19771
rect 15393 19669 15427 19703
rect 22109 19669 22143 19703
rect 23765 19669 23799 19703
rect 30113 19669 30147 19703
rect 44465 19669 44499 19703
rect 40877 19465 40911 19499
rect 44005 19465 44039 19499
rect 46213 19465 46247 19499
rect 47685 19465 47719 19499
rect 8217 19397 8251 19431
rect 14381 19397 14415 19431
rect 16773 19397 16807 19431
rect 19257 19397 19291 19431
rect 23397 19397 23431 19431
rect 27169 19397 27203 19431
rect 27353 19397 27387 19431
rect 1777 19329 1811 19363
rect 8033 19329 8067 19363
rect 11897 19329 11931 19363
rect 12449 19329 12483 19363
rect 13185 19329 13219 19363
rect 14197 19329 14231 19363
rect 16681 19329 16715 19363
rect 17417 19329 17451 19363
rect 19717 19329 19751 19363
rect 21925 19329 21959 19363
rect 23121 19329 23155 19363
rect 25789 19329 25823 19363
rect 26157 19329 26191 19363
rect 28365 19329 28399 19363
rect 28549 19329 28583 19363
rect 29653 19329 29687 19363
rect 30757 19329 30791 19363
rect 30941 19329 30975 19363
rect 31309 19329 31343 19363
rect 32137 19329 32171 19363
rect 40785 19329 40819 19363
rect 43913 19329 43947 19363
rect 44097 19329 44131 19363
rect 44833 19329 44867 19363
rect 46121 19329 46155 19363
rect 46305 19329 46339 19363
rect 47593 19329 47627 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 8585 19261 8619 19295
rect 14657 19261 14691 19295
rect 17601 19261 17635 19295
rect 27537 19261 27571 19295
rect 29745 19261 29779 19295
rect 30205 19261 30239 19295
rect 45109 19261 45143 19295
rect 45661 19261 45695 19295
rect 24869 19193 24903 19227
rect 28457 19193 28491 19227
rect 47041 19193 47075 19227
rect 11713 19125 11747 19159
rect 12633 19125 12667 19159
rect 13277 19125 13311 19159
rect 19901 19125 19935 19159
rect 22017 19125 22051 19159
rect 31217 19125 31251 19159
rect 32229 19125 32263 19159
rect 2237 18921 2271 18955
rect 8309 18921 8343 18955
rect 33333 18921 33367 18955
rect 44281 18921 44315 18955
rect 18337 18853 18371 18887
rect 31125 18853 31159 18887
rect 43269 18853 43303 18887
rect 11805 18785 11839 18819
rect 19257 18785 19291 18819
rect 19441 18785 19475 18819
rect 21925 18785 21959 18819
rect 22293 18785 22327 18819
rect 28089 18785 28123 18819
rect 29837 18785 29871 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 8217 18717 8251 18751
rect 9137 18717 9171 18751
rect 14473 18717 14507 18751
rect 15301 18717 15335 18751
rect 16589 18717 16623 18751
rect 21741 18717 21775 18751
rect 25053 18717 25087 18751
rect 25237 18717 25271 18751
rect 25697 18717 25731 18751
rect 26709 18717 26743 18751
rect 27169 18717 27203 18751
rect 27445 18717 27479 18751
rect 27813 18717 27847 18751
rect 28641 18717 28675 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 30205 18717 30239 18751
rect 30389 18717 30423 18751
rect 30849 18717 30883 18751
rect 31677 18717 31711 18751
rect 32597 18717 32631 18751
rect 43269 18717 43303 18751
rect 43453 18717 43487 18751
rect 44189 18717 44223 18751
rect 44373 18717 44407 18751
rect 45017 18717 45051 18751
rect 45201 18717 45235 18751
rect 46305 18717 46339 18751
rect 9413 18649 9447 18683
rect 12081 18649 12115 18683
rect 15669 18649 15703 18683
rect 16865 18649 16899 18683
rect 21097 18649 21131 18683
rect 25973 18649 26007 18683
rect 45385 18649 45419 18683
rect 46489 18649 46523 18683
rect 10885 18581 10919 18615
rect 13553 18581 13587 18615
rect 14657 18581 14691 18615
rect 9045 18377 9079 18411
rect 9597 18377 9631 18411
rect 10885 18377 10919 18411
rect 11897 18377 11931 18411
rect 12081 18377 12115 18411
rect 17509 18377 17543 18411
rect 18153 18377 18187 18411
rect 46029 18377 46063 18411
rect 47685 18377 47719 18411
rect 16129 18309 16163 18343
rect 29837 18309 29871 18343
rect 32321 18309 32355 18343
rect 1409 18241 1443 18275
rect 2145 18241 2179 18275
rect 9045 18241 9079 18275
rect 9781 18241 9815 18275
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 10793 18241 10827 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 11805 18241 11839 18275
rect 12725 18241 12759 18275
rect 13553 18241 13587 18275
rect 14289 18241 14323 18275
rect 16681 18241 16715 18275
rect 17417 18241 17451 18275
rect 18061 18241 18095 18275
rect 20453 18241 20487 18275
rect 21833 18241 21867 18275
rect 26065 18241 26099 18275
rect 32137 18241 32171 18275
rect 44189 18241 44223 18275
rect 44649 18241 44683 18275
rect 45017 18241 45051 18275
rect 45937 18241 45971 18275
rect 46121 18241 46155 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 12633 18173 12667 18207
rect 13093 18173 13127 18207
rect 14473 18173 14507 18207
rect 20545 18173 20579 18207
rect 26157 18173 26191 18207
rect 27169 18173 27203 18207
rect 27353 18173 27387 18207
rect 27905 18173 27939 18207
rect 29653 18173 29687 18207
rect 31493 18173 31527 18207
rect 33977 18173 34011 18207
rect 45293 18173 45327 18207
rect 1593 18105 1627 18139
rect 26433 18105 26467 18139
rect 45385 18105 45419 18139
rect 2237 18037 2271 18071
rect 13645 18037 13679 18071
rect 16865 18037 16899 18071
rect 20821 18037 20855 18071
rect 21925 18037 21959 18071
rect 14657 17833 14691 17867
rect 23581 17833 23615 17867
rect 27261 17833 27295 17867
rect 27813 17833 27847 17867
rect 28917 17833 28951 17867
rect 30021 17833 30055 17867
rect 44465 17833 44499 17867
rect 45293 17833 45327 17867
rect 10793 17765 10827 17799
rect 29929 17765 29963 17799
rect 21189 17697 21223 17731
rect 25605 17697 25639 17731
rect 26341 17697 26375 17731
rect 2053 17629 2087 17663
rect 10977 17629 11011 17663
rect 11345 17629 11379 17663
rect 11805 17629 11839 17663
rect 14565 17629 14599 17663
rect 17601 17629 17635 17663
rect 20729 17629 20763 17663
rect 23397 17629 23431 17663
rect 26893 17629 26927 17663
rect 27077 17629 27111 17663
rect 27721 17629 27755 17663
rect 28825 17629 28859 17663
rect 29561 17629 29595 17663
rect 44097 17629 44131 17663
rect 44281 17629 44315 17663
rect 46305 17629 46339 17663
rect 11069 17561 11103 17595
rect 12081 17561 12115 17595
rect 15209 17561 15243 17595
rect 20913 17561 20947 17595
rect 23029 17561 23063 17595
rect 23213 17561 23247 17595
rect 45017 17561 45051 17595
rect 45201 17561 45235 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 11161 17493 11195 17527
rect 13553 17493 13587 17527
rect 16497 17493 16531 17527
rect 17601 17493 17635 17527
rect 23305 17493 23339 17527
rect 11897 17289 11931 17323
rect 13185 17289 13219 17323
rect 21189 17289 21223 17323
rect 23137 17289 23171 17323
rect 25513 17289 25547 17323
rect 27169 17289 27203 17323
rect 46213 17289 46247 17323
rect 47685 17289 47719 17323
rect 1961 17221 1995 17255
rect 11529 17221 11563 17255
rect 11745 17221 11779 17255
rect 22937 17221 22971 17255
rect 23949 17221 23983 17255
rect 44373 17221 44407 17255
rect 1777 17153 1811 17187
rect 12357 17153 12391 17187
rect 12541 17153 12575 17187
rect 12633 17153 12667 17187
rect 13093 17153 13127 17187
rect 14381 17153 14415 17187
rect 15209 17153 15243 17187
rect 16865 17153 16899 17187
rect 23765 17153 23799 17187
rect 24041 17153 24075 17187
rect 25421 17153 25455 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 44281 17153 44315 17187
rect 44465 17153 44499 17187
rect 46397 17153 46431 17187
rect 47041 17153 47075 17187
rect 47593 17153 47627 17187
rect 2789 17085 2823 17119
rect 15945 17085 15979 17119
rect 17141 17085 17175 17119
rect 18613 17085 18647 17119
rect 19441 17085 19475 17119
rect 19717 17085 19751 17119
rect 11713 16949 11747 16983
rect 12357 16949 12391 16983
rect 14473 16949 14507 16983
rect 23121 16949 23155 16983
rect 23305 16949 23339 16983
rect 23765 16949 23799 16983
rect 11897 16745 11931 16779
rect 16957 16745 16991 16779
rect 19533 16745 19567 16779
rect 14381 16609 14415 16643
rect 14565 16609 14599 16643
rect 22109 16609 22143 16643
rect 22385 16609 22419 16643
rect 25881 16609 25915 16643
rect 27537 16609 27571 16643
rect 46305 16609 46339 16643
rect 11897 16541 11931 16575
rect 12081 16541 12115 16575
rect 16773 16541 16807 16575
rect 17509 16541 17543 16575
rect 18521 16541 18555 16575
rect 18613 16541 18647 16575
rect 19349 16541 19383 16575
rect 20361 16541 20395 16575
rect 20453 16541 20487 16575
rect 21189 16541 21223 16575
rect 22017 16541 22051 16575
rect 22837 16541 22871 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 24409 16541 24443 16575
rect 28825 16541 28859 16575
rect 29561 16541 29595 16575
rect 31401 16541 31435 16575
rect 16221 16473 16255 16507
rect 26065 16473 26099 16507
rect 28917 16473 28951 16507
rect 29745 16473 29779 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 17601 16405 17635 16439
rect 21281 16405 21315 16439
rect 22937 16405 22971 16439
rect 23581 16405 23615 16439
rect 24501 16405 24535 16439
rect 18337 16201 18371 16235
rect 46857 16201 46891 16235
rect 16865 16133 16899 16167
rect 11713 16065 11747 16099
rect 12265 16065 12299 16099
rect 14657 16065 14691 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 16681 16065 16715 16099
rect 17049 16065 17083 16099
rect 17693 16065 17727 16099
rect 17877 16065 17911 16099
rect 18521 16065 18555 16099
rect 19073 16065 19107 16099
rect 20913 16065 20947 16099
rect 22845 16065 22879 16099
rect 25237 16065 25271 16099
rect 25973 16065 26007 16099
rect 26065 16065 26099 16099
rect 28181 16065 28215 16099
rect 30021 16065 30055 16099
rect 46765 16065 46799 16099
rect 47777 16065 47811 16099
rect 16037 15997 16071 16031
rect 17509 15997 17543 16031
rect 23121 15997 23155 16031
rect 24593 15997 24627 16031
rect 28365 15997 28399 16031
rect 11529 15861 11563 15895
rect 12357 15861 12391 15895
rect 14749 15861 14783 15895
rect 19165 15861 19199 15895
rect 21097 15861 21131 15895
rect 25329 15861 25363 15895
rect 22845 15657 22879 15691
rect 10609 15589 10643 15623
rect 10333 15521 10367 15555
rect 11069 15521 11103 15555
rect 11345 15521 11379 15555
rect 13093 15521 13127 15555
rect 15669 15521 15703 15555
rect 17141 15521 17175 15555
rect 21097 15521 21131 15555
rect 21373 15521 21407 15555
rect 25329 15521 25363 15555
rect 26709 15521 26743 15555
rect 2053 15453 2087 15487
rect 10241 15453 10275 15487
rect 15393 15453 15427 15487
rect 17233 15453 17267 15487
rect 18061 15453 18095 15487
rect 25145 15453 25179 15487
rect 14565 15385 14599 15419
rect 14841 15317 14875 15351
rect 17601 15317 17635 15351
rect 18245 15317 18279 15351
rect 15025 15113 15059 15147
rect 19809 15113 19843 15147
rect 15117 15045 15151 15079
rect 18337 15045 18371 15079
rect 1777 14977 1811 15011
rect 11713 14977 11747 15011
rect 12541 14977 12575 15011
rect 13185 14977 13219 15011
rect 15209 14977 15243 15011
rect 16129 14977 16163 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 18061 14977 18095 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 12357 14909 12391 14943
rect 15393 14909 15427 14943
rect 16957 14909 16991 14943
rect 17141 14909 17175 14943
rect 14841 14841 14875 14875
rect 11529 14773 11563 14807
rect 12725 14773 12759 14807
rect 13277 14773 13311 14807
rect 15945 14773 15979 14807
rect 16681 14773 16715 14807
rect 2237 14569 2271 14603
rect 15945 14501 15979 14535
rect 17233 14501 17267 14535
rect 11437 14433 11471 14467
rect 2145 14365 2179 14399
rect 15117 14365 15151 14399
rect 16221 14365 16255 14399
rect 16313 14365 16347 14399
rect 18061 14365 18095 14399
rect 19349 14365 19383 14399
rect 11713 14297 11747 14331
rect 14933 14297 14967 14331
rect 15301 14297 15335 14331
rect 16129 14297 16163 14331
rect 16957 14297 16991 14331
rect 13185 14229 13219 14263
rect 15209 14229 15243 14263
rect 15485 14229 15519 14263
rect 16497 14229 16531 14263
rect 17417 14229 17451 14263
rect 17877 14229 17911 14263
rect 19533 14229 19567 14263
rect 11897 14025 11931 14059
rect 14105 14025 14139 14059
rect 19073 14025 19107 14059
rect 13737 13957 13771 13991
rect 13953 13957 13987 13991
rect 17601 13957 17635 13991
rect 12081 13889 12115 13923
rect 12357 13889 12391 13923
rect 12541 13889 12575 13923
rect 17325 13821 17359 13855
rect 13921 13685 13955 13719
rect 12633 13481 12667 13515
rect 15669 13481 15703 13515
rect 15853 13481 15887 13515
rect 17417 13481 17451 13515
rect 18521 13481 18555 13515
rect 12817 13413 12851 13447
rect 16589 13277 16623 13311
rect 17233 13277 17267 13311
rect 18429 13277 18463 13311
rect 12449 13209 12483 13243
rect 15485 13209 15519 13243
rect 15701 13209 15735 13243
rect 12659 13141 12693 13175
rect 16681 13141 16715 13175
rect 1593 12937 1627 12971
rect 1409 12801 1443 12835
rect 11989 12801 12023 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 12081 12733 12115 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 12357 12665 12391 12699
rect 14565 12597 14599 12631
rect 15209 12597 15243 12631
rect 47777 12597 47811 12631
rect 12725 12393 12759 12427
rect 14197 12393 14231 12427
rect 16313 12325 16347 12359
rect 16037 12257 16071 12291
rect 16773 12257 16807 12291
rect 17049 12257 17083 12291
rect 46305 12257 46339 12291
rect 48145 12257 48179 12291
rect 12725 12189 12759 12223
rect 14105 12189 14139 12223
rect 14841 12189 14875 12223
rect 15945 12189 15979 12223
rect 46489 12121 46523 12155
rect 14933 12053 14967 12087
rect 18521 12053 18555 12087
rect 17969 11849 18003 11883
rect 47685 11849 47719 11883
rect 15577 11781 15611 11815
rect 12265 11713 12299 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13737 11713 13771 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 16681 11713 16715 11747
rect 17877 11713 17911 11747
rect 46765 11713 46799 11747
rect 47593 11713 47627 11747
rect 15577 11577 15611 11611
rect 12265 11509 12299 11543
rect 12909 11509 12943 11543
rect 13829 11509 13863 11543
rect 16773 11509 16807 11543
rect 46857 11509 46891 11543
rect 12173 11169 12207 11203
rect 14933 11169 14967 11203
rect 15209 11169 15243 11203
rect 16681 11169 16715 11203
rect 46489 11169 46523 11203
rect 12081 11101 12115 11135
rect 46305 11101 46339 11135
rect 48145 11033 48179 11067
rect 12449 10965 12483 10999
rect 12541 10693 12575 10727
rect 14933 10693 14967 10727
rect 12265 10625 12299 10659
rect 47777 10625 47811 10659
rect 45201 10557 45235 10591
rect 45385 10557 45419 10591
rect 46765 10557 46799 10591
rect 15117 10489 15151 10523
rect 14013 10421 14047 10455
rect 15025 10081 15059 10115
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 14381 10013 14415 10047
rect 15209 9945 15243 9979
rect 16865 9945 16899 9979
rect 46489 9945 46523 9979
rect 14473 9877 14507 9911
rect 14473 9605 14507 9639
rect 16773 9605 16807 9639
rect 47685 9605 47719 9639
rect 13001 9537 13035 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 16681 9537 16715 9571
rect 47041 9537 47075 9571
rect 47593 9537 47627 9571
rect 14749 9469 14783 9503
rect 13093 9333 13127 9367
rect 13737 9333 13771 9367
rect 11713 8993 11747 9027
rect 11897 8993 11931 9027
rect 14289 8993 14323 9027
rect 14749 8993 14783 9027
rect 16589 8993 16623 9027
rect 17969 8993 18003 9027
rect 47317 8993 47351 9027
rect 47593 8925 47627 8959
rect 13553 8857 13587 8891
rect 14473 8857 14507 8891
rect 16773 8857 16807 8891
rect 14289 8517 14323 8551
rect 47777 8517 47811 8551
rect 11713 8449 11747 8483
rect 14105 8449 14139 8483
rect 11897 8381 11931 8415
rect 12449 8381 12483 8415
rect 14841 8381 14875 8415
rect 47961 8313 47995 8347
rect 11805 8041 11839 8075
rect 14565 8041 14599 8075
rect 15209 8041 15243 8075
rect 46305 7905 46339 7939
rect 46765 7905 46799 7939
rect 11713 7837 11747 7871
rect 14473 7837 14507 7871
rect 15117 7837 15151 7871
rect 46489 7769 46523 7803
rect 45017 7429 45051 7463
rect 48145 7361 48179 7395
rect 44925 7293 44959 7327
rect 45201 7293 45235 7327
rect 47961 7225 47995 7259
rect 47317 6817 47351 6851
rect 47593 6817 47627 6851
rect 48145 6273 48179 6307
rect 47961 6069 47995 6103
rect 47317 5729 47351 5763
rect 47593 5661 47627 5695
rect 45661 5253 45695 5287
rect 16681 5185 16715 5219
rect 20085 5185 20119 5219
rect 20729 5185 20763 5219
rect 47869 5185 47903 5219
rect 45569 5117 45603 5151
rect 45845 5117 45879 5151
rect 16773 4981 16807 5015
rect 20177 4981 20211 5015
rect 20821 4981 20855 5015
rect 48053 4981 48087 5015
rect 20729 4777 20763 4811
rect 21373 4777 21407 4811
rect 15301 4641 15335 4675
rect 45845 4641 45879 4675
rect 46305 4641 46339 4675
rect 9597 4573 9631 4607
rect 17601 4573 17635 4607
rect 19349 4573 19383 4607
rect 19993 4573 20027 4607
rect 20085 4573 20119 4607
rect 20637 4573 20671 4607
rect 21281 4573 21315 4607
rect 21925 4573 21959 4607
rect 42901 4573 42935 4607
rect 45385 4573 45419 4607
rect 15485 4505 15519 4539
rect 17141 4505 17175 4539
rect 46029 4505 46063 4539
rect 17693 4437 17727 4471
rect 19441 4437 19475 4471
rect 22017 4437 22051 4471
rect 9413 4097 9447 4131
rect 10425 4097 10459 4131
rect 11529 4097 11563 4131
rect 13737 4097 13771 4131
rect 15945 4097 15979 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 18337 4097 18371 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 20821 4097 20855 4131
rect 22201 4097 22235 4131
rect 22845 4097 22879 4131
rect 25697 4097 25731 4131
rect 33149 4097 33183 4131
rect 39773 4097 39807 4131
rect 42625 4097 42659 4131
rect 43269 4097 43303 4131
rect 46121 4097 46155 4131
rect 46765 4097 46799 4131
rect 47869 4097 47903 4131
rect 2145 4029 2179 4063
rect 2329 4029 2363 4063
rect 3249 4029 3283 4063
rect 7113 4029 7147 4063
rect 7297 4029 7331 4063
rect 8309 4029 8343 4063
rect 29561 4029 29595 4063
rect 29745 4029 29779 4063
rect 31401 4029 31435 4063
rect 43453 4029 43487 4063
rect 44189 4029 44223 4063
rect 46949 3961 46983 3995
rect 9505 3893 9539 3927
rect 10517 3893 10551 3927
rect 11621 3893 11655 3927
rect 13829 3893 13863 3927
rect 16037 3893 16071 3927
rect 17141 3893 17175 3927
rect 17785 3893 17819 3927
rect 18429 3893 18463 3927
rect 19073 3893 19107 3927
rect 19717 3893 19751 3927
rect 20913 3893 20947 3927
rect 22293 3893 22327 3927
rect 22937 3893 22971 3927
rect 25789 3893 25823 3927
rect 33241 3893 33275 3927
rect 39865 3893 39899 3927
rect 42717 3893 42751 3927
rect 46213 3893 46247 3927
rect 48053 3893 48087 3927
rect 3157 3689 3191 3723
rect 3985 3689 4019 3723
rect 8217 3689 8251 3723
rect 17785 3689 17819 3723
rect 18429 3689 18463 3723
rect 19349 3689 19383 3723
rect 6469 3553 6503 3587
rect 9413 3553 9447 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 15393 3553 15427 3587
rect 15853 3553 15887 3587
rect 20269 3553 20303 3587
rect 20545 3553 20579 3587
rect 25329 3553 25363 3587
rect 25605 3553 25639 3587
rect 42625 3553 42659 3587
rect 42809 3553 42843 3587
rect 43177 3553 43211 3587
rect 45201 3553 45235 3587
rect 46489 3553 46523 3587
rect 1685 3485 1719 3519
rect 2145 3485 2179 3519
rect 3065 3485 3099 3519
rect 5181 3485 5215 3519
rect 5825 3485 5859 3519
rect 8125 3485 8159 3519
rect 11897 3485 11931 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 16313 3485 16347 3519
rect 16957 3485 16991 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 19257 3485 19291 3519
rect 20085 3485 20119 3519
rect 22569 3485 22603 3519
rect 23029 3485 23063 3519
rect 23121 3485 23155 3519
rect 23673 3485 23707 3519
rect 24685 3485 24719 3519
rect 25145 3485 25179 3519
rect 33333 3485 33367 3519
rect 36001 3485 36035 3519
rect 37841 3485 37875 3519
rect 39129 3485 39163 3519
rect 40049 3485 40083 3519
rect 40325 3485 40359 3519
rect 41337 3485 41371 3519
rect 41521 3485 41555 3519
rect 45661 3485 45695 3519
rect 46305 3485 46339 3519
rect 5273 3417 5307 3451
rect 6009 3417 6043 3451
rect 36185 3417 36219 3451
rect 48145 3417 48179 3451
rect 2237 3349 2271 3383
rect 16405 3349 16439 3383
rect 17049 3349 17083 3383
rect 23765 3349 23799 3383
rect 39221 3349 39255 3383
rect 41981 3349 42015 3383
rect 45753 3349 45787 3383
rect 16773 3145 16807 3179
rect 17417 3145 17451 3179
rect 19165 3145 19199 3179
rect 20821 3145 20855 3179
rect 1961 3077 1995 3111
rect 8217 3077 8251 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 22293 3077 22327 3111
rect 33241 3077 33275 3111
rect 39037 3077 39071 3111
rect 42625 3077 42659 3111
rect 45385 3077 45419 3111
rect 47777 3077 47811 3111
rect 1777 3009 1811 3043
rect 6561 3009 6595 3043
rect 7389 3009 7423 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 16681 3009 16715 3043
rect 17325 3009 17359 3043
rect 17969 3009 18003 3043
rect 19073 3009 19107 3043
rect 20269 3009 20303 3043
rect 20729 3009 20763 3043
rect 22109 3009 22143 3043
rect 28549 3009 28583 3043
rect 33057 3009 33091 3043
rect 37749 3009 37783 3043
rect 37841 3009 37875 3043
rect 39497 3009 39531 3043
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 2237 2941 2271 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 22569 2941 22603 2975
rect 24409 2941 24443 2975
rect 24593 2941 24627 2975
rect 26157 2941 26191 2975
rect 28733 2941 28767 2975
rect 30389 2941 30423 2975
rect 33517 2941 33551 2975
rect 38393 2941 38427 2975
rect 38577 2941 38611 2975
rect 39681 2941 39715 2975
rect 41337 2941 41371 2975
rect 44281 2941 44315 2975
rect 47041 2941 47075 2975
rect 47961 2873 47995 2907
rect 18061 2805 18095 2839
rect 17509 2601 17543 2635
rect 18153 2601 18187 2635
rect 19717 2601 19751 2635
rect 20453 2601 20487 2635
rect 21925 2601 21959 2635
rect 23673 2601 23707 2635
rect 24961 2601 24995 2635
rect 35725 2601 35759 2635
rect 36277 2601 36311 2635
rect 39221 2601 39255 2635
rect 40417 2601 40451 2635
rect 42993 2601 43027 2635
rect 2145 2533 2179 2567
rect 8217 2533 8251 2567
rect 16865 2533 16899 2567
rect 26433 2533 26467 2567
rect 47961 2533 47995 2567
rect 15577 2465 15611 2499
rect 27629 2465 27663 2499
rect 30021 2465 30055 2499
rect 38393 2465 38427 2499
rect 41337 2465 41371 2499
rect 43913 2465 43947 2499
rect 46213 2465 46247 2499
rect 5457 2397 5491 2431
rect 15301 2397 15335 2431
rect 16681 2397 16715 2431
rect 17417 2397 17451 2431
rect 18061 2397 18095 2431
rect 19625 2397 19659 2431
rect 21281 2397 21315 2431
rect 21925 2397 21959 2431
rect 23029 2397 23063 2431
rect 23857 2397 23891 2431
rect 29745 2397 29779 2431
rect 36461 2397 36495 2431
rect 39129 2397 39163 2431
rect 41061 2397 41095 2431
rect 42901 2397 42935 2431
rect 43637 2397 43671 2431
rect 46489 2397 46523 2431
rect 1869 2329 1903 2363
rect 2789 2329 2823 2363
rect 9413 2329 9447 2363
rect 9781 2329 9815 2363
rect 20361 2329 20395 2363
rect 21097 2329 21131 2363
rect 24869 2329 24903 2363
rect 26249 2329 26283 2363
rect 27445 2329 27479 2363
rect 28549 2329 28583 2363
rect 35633 2329 35667 2363
rect 38209 2329 38243 2363
rect 40325 2329 40359 2363
rect 45385 2329 45419 2363
rect 47777 2329 47811 2363
rect 3065 2261 3099 2295
rect 5273 2261 5307 2295
rect 28641 2261 28675 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 13357 47243 13415 47249
rect 13357 47209 13369 47243
rect 13403 47240 13415 47243
rect 19978 47240 19984 47252
rect 13403 47212 19984 47240
rect 13403 47209 13415 47212
rect 13357 47203 13415 47209
rect 19978 47200 19984 47212
rect 20036 47200 20042 47252
rect 19429 47175 19487 47181
rect 19429 47141 19441 47175
rect 19475 47172 19487 47175
rect 20254 47172 20260 47184
rect 19475 47144 20260 47172
rect 19475 47141 19487 47144
rect 19429 47135 19487 47141
rect 20254 47132 20260 47144
rect 20312 47132 20318 47184
rect 29362 47132 29368 47184
rect 29420 47172 29426 47184
rect 29917 47175 29975 47181
rect 29917 47172 29929 47175
rect 29420 47144 29929 47172
rect 29420 47132 29426 47144
rect 29917 47141 29929 47144
rect 29963 47141 29975 47175
rect 48133 47175 48191 47181
rect 48133 47172 48145 47175
rect 29917 47135 29975 47141
rect 30024 47144 48145 47172
rect 3050 47064 3056 47116
rect 3108 47104 3114 47116
rect 20070 47104 20076 47116
rect 3108 47076 19380 47104
rect 20031 47076 20076 47104
rect 3108 47064 3114 47076
rect 1946 46996 1952 47048
rect 2004 47036 2010 47048
rect 2041 47039 2099 47045
rect 2041 47036 2053 47039
rect 2004 47008 2053 47036
rect 2004 46996 2010 47008
rect 2041 47005 2053 47008
rect 2087 47005 2099 47039
rect 2041 46999 2099 47005
rect 2774 46996 2780 47048
rect 2832 47036 2838 47048
rect 2961 47039 3019 47045
rect 2961 47036 2973 47039
rect 2832 47008 2973 47036
rect 2832 46996 2838 47008
rect 2961 47005 2973 47008
rect 3007 47005 3019 47039
rect 2961 46999 3019 47005
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6825 47039 6883 47045
rect 6825 47036 6837 47039
rect 5868 47008 6837 47036
rect 5868 46996 5874 47008
rect 6825 47005 6837 47008
rect 6871 47005 6883 47039
rect 6825 46999 6883 47005
rect 7098 46996 7104 47048
rect 7156 47036 7162 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7156 47008 7757 47036
rect 7156 46996 7162 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 7745 46999 7803 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9125 47039 9183 47045
rect 9125 47036 9137 47039
rect 9088 47008 9137 47036
rect 9088 46996 9094 47008
rect 9125 47005 9137 47008
rect 9171 47005 9183 47039
rect 9125 46999 9183 47005
rect 11606 46996 11612 47048
rect 11664 47036 11670 47048
rect 11701 47039 11759 47045
rect 11701 47036 11713 47039
rect 11664 47008 11713 47036
rect 11664 46996 11670 47008
rect 11701 47005 11713 47008
rect 11747 47005 11759 47039
rect 11974 47036 11980 47048
rect 11935 47008 11980 47036
rect 11701 46999 11759 47005
rect 11974 46996 11980 47008
rect 12032 46996 12038 47048
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 15289 47039 15347 47045
rect 15289 47036 15301 47039
rect 13872 47008 15301 47036
rect 13872 46996 13878 47008
rect 15289 47005 15301 47008
rect 15335 47005 15347 47039
rect 15289 46999 15347 47005
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16942 47036 16948 47048
rect 16903 47008 16948 47036
rect 16669 46999 16727 47005
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 19245 46999 19303 47005
rect 2314 46968 2320 46980
rect 2275 46940 2320 46968
rect 2314 46928 2320 46940
rect 2372 46928 2378 46980
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 7834 46928 7840 46980
rect 7892 46968 7898 46980
rect 7929 46971 7987 46977
rect 7929 46968 7941 46971
rect 7892 46940 7941 46968
rect 7892 46928 7898 46940
rect 7929 46937 7941 46940
rect 7975 46937 7987 46971
rect 14553 46971 14611 46977
rect 14553 46968 14565 46971
rect 7929 46931 7987 46937
rect 13464 46940 14565 46968
rect 3142 46900 3148 46912
rect 3103 46872 3148 46900
rect 3142 46860 3148 46872
rect 3200 46860 3206 46912
rect 6914 46860 6920 46912
rect 6972 46900 6978 46912
rect 9306 46900 9312 46912
rect 6972 46872 7017 46900
rect 9267 46872 9312 46900
rect 6972 46860 6978 46872
rect 9306 46860 9312 46872
rect 9364 46860 9370 46912
rect 12250 46860 12256 46912
rect 12308 46900 12314 46912
rect 13464 46900 13492 46940
rect 14553 46937 14565 46940
rect 14599 46937 14611 46971
rect 14553 46931 14611 46937
rect 14642 46928 14648 46980
rect 14700 46968 14706 46980
rect 14737 46971 14795 46977
rect 14737 46968 14749 46971
rect 14700 46940 14749 46968
rect 14700 46928 14706 46940
rect 14737 46937 14749 46940
rect 14783 46937 14795 46971
rect 14737 46931 14795 46937
rect 15378 46928 15384 46980
rect 15436 46968 15442 46980
rect 15473 46971 15531 46977
rect 15473 46968 15485 46971
rect 15436 46940 15485 46968
rect 15436 46928 15442 46940
rect 15473 46937 15485 46940
rect 15519 46937 15531 46971
rect 19352 46968 19380 47076
rect 20070 47064 20076 47076
rect 20128 47064 20134 47116
rect 26602 47064 26608 47116
rect 26660 47104 26666 47116
rect 30024 47104 30052 47144
rect 48133 47141 48145 47144
rect 48179 47141 48191 47175
rect 48133 47135 48191 47141
rect 30742 47104 30748 47116
rect 26660 47076 30052 47104
rect 30703 47076 30748 47104
rect 26660 47064 26666 47076
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 46750 47104 46756 47116
rect 35866 47076 46756 47104
rect 20346 47036 20352 47048
rect 20307 47008 20352 47036
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 24578 46996 24584 47048
rect 24636 47036 24642 47048
rect 24765 47039 24823 47045
rect 24765 47036 24777 47039
rect 24636 47008 24777 47036
rect 24636 46996 24642 47008
rect 24765 47005 24777 47008
rect 24811 47005 24823 47039
rect 25406 47036 25412 47048
rect 25367 47008 25412 47036
rect 24765 46999 24823 47005
rect 25406 46996 25412 47008
rect 25464 46996 25470 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28629 47039 28687 47045
rect 28629 47036 28641 47039
rect 28408 47008 28641 47036
rect 28408 46996 28414 47008
rect 28629 47005 28641 47008
rect 28675 47005 28687 47039
rect 28629 46999 28687 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 31018 47036 31024 47048
rect 30979 47008 31024 47036
rect 29733 46999 29791 47005
rect 31018 46996 31024 47008
rect 31076 46996 31082 47048
rect 22186 46968 22192 46980
rect 19352 46940 22192 46968
rect 15473 46931 15531 46937
rect 22186 46928 22192 46940
rect 22244 46928 22250 46980
rect 26694 46928 26700 46980
rect 26752 46968 26758 46980
rect 35866 46968 35894 47076
rect 46750 47064 46756 47076
rect 46808 47064 46814 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38289 47039 38347 47045
rect 38289 47036 38301 47039
rect 38160 47008 38301 47036
rect 38160 46996 38166 47008
rect 38289 47005 38301 47008
rect 38335 47005 38347 47039
rect 41874 47036 41880 47048
rect 41835 47008 41880 47036
rect 38289 46999 38347 47005
rect 41874 46996 41880 47008
rect 41932 46996 41938 47048
rect 42610 47036 42616 47048
rect 42571 47008 42616 47036
rect 42610 46996 42616 47008
rect 42668 46996 42674 47048
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47949 47039 48007 47045
rect 47949 47036 47961 47039
rect 47728 47008 47961 47036
rect 47728 46996 47734 47008
rect 47949 47005 47961 47008
rect 47995 47005 48007 47039
rect 47949 46999 48007 47005
rect 26752 46940 35894 46968
rect 40313 46971 40371 46977
rect 26752 46928 26758 46940
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 12308 46872 13492 46900
rect 12308 46860 12314 46872
rect 28258 46860 28264 46912
rect 28316 46900 28322 46912
rect 28445 46903 28503 46909
rect 28445 46900 28457 46903
rect 28316 46872 28457 46900
rect 28316 46860 28322 46872
rect 28445 46869 28457 46872
rect 28491 46869 28503 46903
rect 28445 46863 28503 46869
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 42794 46968 42800 46980
rect 42755 46940 42800 46968
rect 40497 46931 40555 46937
rect 42794 46928 42800 46940
rect 42852 46928 42858 46980
rect 44453 46971 44511 46977
rect 44453 46937 44465 46971
rect 44499 46937 44511 46971
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 44453 46931 44511 46937
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 43162 46860 43168 46912
rect 43220 46900 43226 46912
rect 44468 46900 44496 46931
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 43220 46872 44496 46900
rect 43220 46860 43226 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 3142 46588 3148 46640
rect 3200 46628 3206 46640
rect 28445 46631 28503 46637
rect 28445 46628 28457 46631
rect 3200 46600 28457 46628
rect 3200 46588 3206 46600
rect 28445 46597 28457 46600
rect 28491 46597 28503 46631
rect 28445 46591 28503 46597
rect 30101 46631 30159 46637
rect 30101 46597 30113 46631
rect 30147 46628 30159 46631
rect 30147 46600 35894 46628
rect 30147 46597 30159 46600
rect 30101 46591 30159 46597
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 24578 46560 24584 46572
rect 24539 46532 24584 46560
rect 24578 46520 24584 46532
rect 24636 46520 24642 46572
rect 28258 46560 28264 46572
rect 28219 46532 28264 46560
rect 28258 46520 28264 46532
rect 28316 46520 28322 46572
rect 2961 46495 3019 46501
rect 2961 46461 2973 46495
rect 3007 46492 3019 46495
rect 3421 46495 3479 46501
rect 3421 46492 3433 46495
rect 3007 46464 3433 46492
rect 3007 46461 3019 46464
rect 2961 46455 3019 46461
rect 3421 46461 3433 46464
rect 3467 46461 3479 46495
rect 3421 46455 3479 46461
rect 3605 46495 3663 46501
rect 3605 46461 3617 46495
rect 3651 46492 3663 46495
rect 3878 46492 3884 46504
rect 3651 46464 3884 46492
rect 3651 46461 3663 46464
rect 3605 46455 3663 46461
rect 3878 46452 3884 46464
rect 3936 46452 3942 46504
rect 3970 46452 3976 46504
rect 4028 46492 4034 46504
rect 4157 46495 4215 46501
rect 4157 46492 4169 46495
rect 4028 46464 4169 46492
rect 4028 46452 4034 46464
rect 4157 46461 4169 46464
rect 4203 46461 4215 46495
rect 4157 46455 4215 46461
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11698 46492 11704 46504
rect 11659 46464 11704 46492
rect 11517 46455 11575 46461
rect 11698 46452 11704 46464
rect 11756 46452 11762 46504
rect 11977 46495 12035 46501
rect 11977 46461 11989 46495
rect 12023 46461 12035 46495
rect 13814 46492 13820 46504
rect 13775 46464 13820 46492
rect 11977 46455 12035 46461
rect 11992 46424 12020 46455
rect 13814 46452 13820 46464
rect 13872 46452 13878 46504
rect 13998 46492 14004 46504
rect 13959 46464 14004 46492
rect 13998 46452 14004 46464
rect 14056 46452 14062 46504
rect 14182 46452 14188 46504
rect 14240 46492 14246 46504
rect 14277 46495 14335 46501
rect 14277 46492 14289 46495
rect 14240 46464 14289 46492
rect 14240 46452 14246 46464
rect 14277 46461 14289 46464
rect 14323 46461 14335 46495
rect 19426 46492 19432 46504
rect 19387 46464 19432 46492
rect 14277 46455 14335 46461
rect 19426 46452 19432 46464
rect 19484 46452 19490 46504
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20162 46492 20168 46504
rect 19659 46464 20168 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 20162 46452 20168 46464
rect 20220 46452 20226 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 32585 46455 32643 46461
rect 10980 46396 12020 46424
rect 10980 46368 11008 46396
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 32272 46396 32628 46424
rect 35866 46424 35894 46600
rect 38378 46588 38384 46640
rect 38436 46628 38442 46640
rect 46750 46628 46756 46640
rect 38436 46600 46756 46628
rect 38436 46588 38442 46600
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 41708 46569 41736 46600
rect 46750 46588 46756 46600
rect 46808 46588 46814 46640
rect 41693 46563 41751 46569
rect 41693 46529 41705 46563
rect 41739 46529 41751 46563
rect 41693 46523 41751 46529
rect 41874 46520 41880 46572
rect 41932 46560 41938 46572
rect 42429 46563 42487 46569
rect 42429 46560 42441 46563
rect 41932 46532 42441 46560
rect 41932 46520 41938 46532
rect 42429 46529 42441 46532
rect 42475 46529 42487 46563
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 42429 46523 42487 46529
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41785 46495 41843 46501
rect 41785 46461 41797 46495
rect 41831 46492 41843 46495
rect 42613 46495 42671 46501
rect 42613 46492 42625 46495
rect 41831 46464 42625 46492
rect 41831 46461 41843 46464
rect 41785 46455 41843 46461
rect 42613 46461 42625 46464
rect 42659 46461 42671 46495
rect 42613 46455 42671 46461
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46290 46492 46296 46504
rect 45419 46464 46296 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 35866 46396 41460 46424
rect 32272 46384 32278 46396
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 1670 46356 1676 46368
rect 1627 46328 1676 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 1946 46316 1952 46368
rect 2004 46356 2010 46368
rect 2317 46359 2375 46365
rect 2317 46356 2329 46359
rect 2004 46328 2329 46356
rect 2004 46316 2010 46328
rect 2317 46325 2329 46328
rect 2363 46325 2375 46359
rect 2317 46319 2375 46325
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 20714 46316 20720 46368
rect 20772 46356 20778 46368
rect 22005 46359 22063 46365
rect 22005 46356 22017 46359
rect 20772 46328 22017 46356
rect 20772 46316 20778 46328
rect 22005 46325 22017 46328
rect 22051 46325 22063 46359
rect 22005 46319 22063 46325
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 41432 46356 41460 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 42576 46396 42932 46424
rect 45204 46424 45232 46455
rect 46290 46452 46296 46464
rect 46348 46452 46354 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 47762 46424 47768 46436
rect 45204 46396 47768 46424
rect 42576 46384 42582 46396
rect 47762 46384 47768 46396
rect 47820 46384 47826 46436
rect 43530 46356 43536 46368
rect 41432 46328 43536 46356
rect 43530 46316 43536 46328
rect 43588 46316 43594 46368
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3878 46152 3884 46164
rect 3839 46124 3884 46152
rect 3878 46112 3884 46124
rect 3936 46112 3942 46164
rect 11241 46155 11299 46161
rect 11241 46121 11253 46155
rect 11287 46152 11299 46155
rect 11698 46152 11704 46164
rect 11287 46124 11704 46152
rect 11287 46121 11299 46124
rect 11241 46115 11299 46121
rect 11698 46112 11704 46124
rect 11756 46112 11762 46164
rect 13814 46112 13820 46164
rect 13872 46152 13878 46164
rect 14277 46155 14335 46161
rect 14277 46152 14289 46155
rect 13872 46124 14289 46152
rect 13872 46112 13878 46124
rect 14277 46121 14289 46124
rect 14323 46121 14335 46155
rect 20162 46152 20168 46164
rect 20123 46124 20168 46152
rect 14277 46115 14335 46121
rect 20162 46112 20168 46124
rect 20220 46112 20226 46164
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 20714 46016 20720 46028
rect 20675 45988 20720 46016
rect 20714 45976 20720 45988
rect 20772 45976 20778 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25406 46016 25412 46028
rect 25271 45988 25412 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25406 45976 25412 45988
rect 25464 45976 25470 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 41322 46016 41328 46028
rect 41283 45988 41328 46016
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41966 46016 41972 46028
rect 41927 45988 41972 46016
rect 41966 45976 41972 45988
rect 42024 45976 42030 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 2777 45951 2835 45957
rect 2777 45917 2789 45951
rect 2823 45948 2835 45951
rect 3789 45951 3847 45957
rect 3789 45948 3801 45951
rect 2823 45920 3801 45948
rect 2823 45917 2835 45920
rect 2777 45911 2835 45917
rect 3789 45917 3801 45920
rect 3835 45948 3847 45951
rect 11149 45951 11207 45957
rect 3835 45920 6914 45948
rect 3835 45917 3847 45920
rect 3789 45911 3847 45917
rect 2866 45812 2872 45824
rect 2827 45784 2872 45812
rect 2866 45772 2872 45784
rect 2924 45772 2930 45824
rect 6886 45812 6914 45920
rect 11149 45917 11161 45951
rect 11195 45948 11207 45951
rect 14090 45948 14096 45960
rect 11195 45920 14096 45948
rect 11195 45917 11207 45920
rect 11149 45911 11207 45917
rect 14090 45908 14096 45920
rect 14148 45908 14154 45960
rect 20070 45948 20076 45960
rect 20031 45920 20076 45948
rect 20070 45908 20076 45920
rect 20128 45908 20134 45960
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45948 24639 45951
rect 24670 45948 24676 45960
rect 24627 45920 24676 45948
rect 24627 45917 24639 45920
rect 24581 45911 24639 45917
rect 24670 45908 24676 45920
rect 24728 45908 24734 45960
rect 38194 45948 38200 45960
rect 38107 45920 38200 45948
rect 38194 45908 38200 45920
rect 38252 45948 38258 45960
rect 38378 45948 38384 45960
rect 38252 45920 38384 45948
rect 38252 45908 38258 45920
rect 38378 45908 38384 45920
rect 38436 45908 38442 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43993 45951 44051 45957
rect 43993 45948 44005 45951
rect 43864 45920 44005 45948
rect 43864 45908 43870 45920
rect 43993 45917 44005 45920
rect 44039 45917 44051 45951
rect 43993 45911 44051 45917
rect 45557 45951 45615 45957
rect 45557 45917 45569 45951
rect 45603 45948 45615 45951
rect 45738 45948 45744 45960
rect 45603 45920 45744 45948
rect 45603 45917 45615 45920
rect 45557 45911 45615 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 45830 45908 45836 45960
rect 45888 45948 45894 45960
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45888 45920 46305 45948
rect 45888 45908 45894 45920
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 41506 45880 41512 45892
rect 41467 45852 41512 45880
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 25314 45812 25320 45824
rect 6886 45784 25320 45812
rect 25314 45772 25320 45784
rect 25372 45772 25378 45824
rect 33318 45772 33324 45824
rect 33376 45812 33382 45824
rect 44085 45815 44143 45821
rect 44085 45812 44097 45815
rect 33376 45784 44097 45812
rect 33376 45772 33382 45784
rect 44085 45781 44097 45784
rect 44131 45781 44143 45815
rect 44085 45775 44143 45781
rect 45554 45772 45560 45824
rect 45612 45812 45618 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 45612 45784 45753 45812
rect 45612 45772 45618 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 13817 45611 13875 45617
rect 13817 45577 13829 45611
rect 13863 45608 13875 45611
rect 13998 45608 14004 45620
rect 13863 45580 14004 45608
rect 13863 45577 13875 45580
rect 13817 45571 13875 45577
rect 13998 45568 14004 45580
rect 14056 45568 14062 45620
rect 14090 45568 14096 45620
rect 14148 45608 14154 45620
rect 20898 45608 20904 45620
rect 14148 45580 20760 45608
rect 20859 45580 20904 45608
rect 14148 45568 14154 45580
rect 2133 45543 2191 45549
rect 2133 45509 2145 45543
rect 2179 45540 2191 45543
rect 2866 45540 2872 45552
rect 2179 45512 2872 45540
rect 2179 45509 2191 45512
rect 2133 45503 2191 45509
rect 2866 45500 2872 45512
rect 2924 45500 2930 45552
rect 20732 45540 20760 45580
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 25317 45611 25375 45617
rect 25317 45577 25329 45611
rect 25363 45608 25375 45611
rect 25406 45608 25412 45620
rect 25363 45580 25412 45608
rect 25363 45577 25375 45580
rect 25317 45571 25375 45577
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 32217 45611 32275 45617
rect 32217 45577 32229 45611
rect 32263 45608 32275 45611
rect 32306 45608 32312 45620
rect 32263 45580 32312 45608
rect 32263 45577 32275 45580
rect 32217 45571 32275 45577
rect 32306 45568 32312 45580
rect 32364 45568 32370 45620
rect 41417 45611 41475 45617
rect 41417 45577 41429 45611
rect 41463 45608 41475 45611
rect 41506 45608 41512 45620
rect 41463 45580 41512 45608
rect 41463 45577 41475 45580
rect 41417 45571 41475 45577
rect 41506 45568 41512 45580
rect 41564 45568 41570 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45646 45608 45652 45620
rect 45152 45580 45652 45608
rect 45152 45568 45158 45580
rect 45646 45568 45652 45580
rect 45704 45568 45710 45620
rect 46382 45568 46388 45620
rect 46440 45608 46446 45620
rect 46440 45580 47992 45608
rect 46440 45568 46446 45580
rect 24670 45540 24676 45552
rect 20732 45512 24676 45540
rect 1946 45472 1952 45484
rect 1907 45444 1952 45472
rect 1946 45432 1952 45444
rect 2004 45432 2010 45484
rect 13722 45472 13728 45484
rect 13683 45444 13728 45472
rect 13722 45432 13728 45444
rect 13780 45432 13786 45484
rect 19426 45432 19432 45484
rect 19484 45472 19490 45484
rect 20824 45481 20852 45512
rect 24670 45500 24676 45512
rect 24728 45500 24734 45552
rect 40678 45540 40684 45552
rect 26206 45512 40684 45540
rect 20257 45475 20315 45481
rect 20257 45472 20269 45475
rect 19484 45444 20269 45472
rect 19484 45432 19490 45444
rect 20257 45441 20269 45444
rect 20303 45441 20315 45475
rect 20257 45435 20315 45441
rect 20809 45475 20867 45481
rect 20809 45441 20821 45475
rect 20855 45472 20867 45475
rect 25225 45475 25283 45481
rect 20855 45444 20889 45472
rect 20855 45441 20867 45444
rect 20809 45435 20867 45441
rect 25225 45441 25237 45475
rect 25271 45472 25283 45475
rect 25314 45472 25320 45484
rect 25271 45444 25320 45472
rect 25271 45441 25283 45444
rect 25225 45435 25283 45441
rect 25314 45432 25320 45444
rect 25372 45432 25378 45484
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 20070 45364 20076 45416
rect 20128 45404 20134 45416
rect 26206 45404 26234 45512
rect 40678 45500 40684 45512
rect 40736 45500 40742 45552
rect 42794 45540 42800 45552
rect 42755 45512 42800 45540
rect 42794 45500 42800 45512
rect 42852 45500 42858 45552
rect 45370 45500 45376 45552
rect 45428 45540 45434 45552
rect 47964 45549 47992 45580
rect 46937 45543 46995 45549
rect 46937 45540 46949 45543
rect 45428 45512 46949 45540
rect 45428 45500 45434 45512
rect 46937 45509 46949 45512
rect 46983 45509 46995 45543
rect 46937 45503 46995 45509
rect 47949 45543 48007 45549
rect 47949 45509 47961 45543
rect 47995 45509 48007 45543
rect 47949 45503 48007 45509
rect 32125 45475 32183 45481
rect 32125 45441 32137 45475
rect 32171 45472 32183 45475
rect 32214 45472 32220 45484
rect 32171 45444 32220 45472
rect 32171 45441 32183 45444
rect 32125 45435 32183 45441
rect 32214 45432 32220 45444
rect 32272 45432 32278 45484
rect 41325 45475 41383 45481
rect 41325 45441 41337 45475
rect 41371 45472 41383 45475
rect 42705 45475 42763 45481
rect 42705 45472 42717 45475
rect 41371 45444 42717 45472
rect 41371 45441 41383 45444
rect 41325 45435 41383 45441
rect 42705 45441 42717 45444
rect 42751 45441 42763 45475
rect 42705 45435 42763 45441
rect 43809 45475 43867 45481
rect 43809 45441 43821 45475
rect 43855 45472 43867 45475
rect 44174 45472 44180 45484
rect 43855 45444 44180 45472
rect 43855 45441 43867 45444
rect 43809 45435 43867 45441
rect 20128 45376 26234 45404
rect 20128 45364 20134 45376
rect 42720 45336 42748 45435
rect 44174 45432 44180 45444
rect 44232 45432 44238 45484
rect 46845 45475 46903 45481
rect 46845 45441 46857 45475
rect 46891 45472 46903 45475
rect 47578 45472 47584 45484
rect 46891 45444 47584 45472
rect 46891 45441 46903 45444
rect 46845 45435 46903 45441
rect 47578 45432 47584 45444
rect 47636 45432 47642 45484
rect 44450 45364 44456 45416
rect 44508 45404 44514 45416
rect 44545 45407 44603 45413
rect 44545 45404 44557 45407
rect 44508 45376 44557 45404
rect 44508 45364 44514 45376
rect 44545 45373 44557 45376
rect 44591 45373 44603 45407
rect 44545 45367 44603 45373
rect 44729 45407 44787 45413
rect 44729 45373 44741 45407
rect 44775 45404 44787 45407
rect 45094 45404 45100 45416
rect 44775 45376 45100 45404
rect 44775 45373 44787 45376
rect 44729 45367 44787 45373
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45646 45404 45652 45416
rect 45607 45376 45652 45404
rect 45646 45364 45652 45376
rect 45704 45364 45710 45416
rect 47394 45404 47400 45416
rect 45756 45376 47400 45404
rect 45756 45336 45784 45376
rect 47394 45364 47400 45376
rect 47452 45364 47458 45416
rect 42720 45308 45784 45336
rect 43990 45268 43996 45280
rect 43951 45240 43996 45268
rect 43990 45228 43996 45240
rect 44048 45228 44054 45280
rect 45462 45228 45468 45280
rect 45520 45268 45526 45280
rect 48041 45271 48099 45277
rect 48041 45268 48053 45271
rect 45520 45240 48053 45268
rect 45520 45228 45526 45240
rect 48041 45237 48053 45240
rect 48087 45237 48099 45271
rect 48041 45231 48099 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 42610 45024 42616 45076
rect 42668 45064 42674 45076
rect 42889 45067 42947 45073
rect 42889 45064 42901 45067
rect 42668 45036 42901 45064
rect 42668 45024 42674 45036
rect 42889 45033 42901 45036
rect 42935 45033 42947 45067
rect 44450 45064 44456 45076
rect 44411 45036 44456 45064
rect 42889 45027 42947 45033
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 40678 44956 40684 45008
rect 40736 44996 40742 45008
rect 47578 44996 47584 45008
rect 40736 44968 47584 44996
rect 40736 44956 40742 44968
rect 47578 44956 47584 44968
rect 47636 44956 47642 45008
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 44910 44820 44916 44872
rect 44968 44860 44974 44872
rect 45005 44863 45063 44869
rect 45005 44860 45017 44863
rect 44968 44832 45017 44860
rect 44968 44820 44974 44832
rect 45005 44829 45017 44832
rect 45051 44829 45063 44863
rect 45646 44860 45652 44872
rect 45607 44832 45652 44860
rect 45005 44823 45063 44829
rect 45646 44820 45652 44832
rect 45704 44820 45710 44872
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 46934 44792 46940 44804
rect 46523 44764 46940 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 46934 44752 46940 44764
rect 46992 44752 46998 44804
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 46290 44520 46296 44532
rect 46251 44492 46296 44520
rect 46290 44480 46296 44492
rect 46348 44480 46354 44532
rect 46934 44520 46940 44532
rect 46895 44492 46940 44520
rect 46934 44480 46940 44492
rect 46992 44480 46998 44532
rect 46014 44412 46020 44464
rect 46072 44452 46078 44464
rect 46072 44424 46888 44452
rect 46072 44412 46078 44424
rect 45097 44387 45155 44393
rect 45097 44353 45109 44387
rect 45143 44384 45155 44387
rect 45186 44384 45192 44396
rect 45143 44356 45192 44384
rect 45143 44353 45155 44356
rect 45097 44347 45155 44353
rect 45186 44344 45192 44356
rect 45244 44344 45250 44396
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46860 44393 46888 44424
rect 46201 44387 46259 44393
rect 46201 44353 46213 44387
rect 46247 44353 46259 44387
rect 46201 44347 46259 44353
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 45646 44276 45652 44328
rect 45704 44316 45710 44328
rect 46216 44316 46244 44347
rect 45704 44288 46244 44316
rect 45704 44276 45710 44288
rect 47670 44180 47676 44192
rect 47631 44152 47676 44180
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47670 43840 47676 43852
rect 46523 43812 47676 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47670 43800 47676 43812
rect 47728 43800 47734 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47762 43296 47768 43308
rect 47723 43268 47768 43296
rect 47762 43256 47768 43268
rect 47820 43256 47826 43308
rect 1486 43188 1492 43240
rect 1544 43228 1550 43240
rect 1581 43231 1639 43237
rect 1581 43228 1593 43231
rect 1544 43200 1593 43228
rect 1544 43188 1550 43200
rect 1581 43197 1593 43200
rect 1627 43197 1639 43231
rect 1581 43191 1639 43197
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47029 42171 47087 42177
rect 47394 42168 47400 42220
rect 47452 42208 47458 42220
rect 47581 42211 47639 42217
rect 47581 42208 47593 42211
rect 47452 42180 47593 42208
rect 47452 42168 47458 42180
rect 47581 42177 47593 42180
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 1636 41228 2237 41256
rect 1636 41216 1642 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 2225 41219 2283 41225
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46845 41259 46903 41265
rect 46845 41256 46857 41259
rect 46532 41228 46857 41256
rect 46532 41216 46538 41228
rect 46845 41225 46857 41228
rect 46891 41225 46903 41259
rect 46845 41219 46903 41225
rect 2133 41123 2191 41129
rect 2133 41089 2145 41123
rect 2179 41120 2191 41123
rect 2406 41120 2412 41132
rect 2179 41092 2412 41120
rect 2179 41089 2191 41092
rect 2133 41083 2191 41089
rect 2406 41080 2412 41092
rect 2464 41080 2470 41132
rect 46750 41120 46756 41132
rect 46711 41092 46756 41120
rect 46750 41080 46756 41092
rect 46808 41080 46814 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 45526 40956 48145 40984
rect 43438 40876 43444 40928
rect 43496 40916 43502 40928
rect 45526 40916 45554 40956
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 43496 40888 45554 40916
rect 43496 40876 43502 40888
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2038 40440 2044 40452
rect 1999 40412 2044 40440
rect 2038 40400 2044 40412
rect 2096 40400 2102 40452
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46934 39352 46940 39364
rect 46523 39324 46940 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46934 39312 46940 39324
rect 46992 39312 46998 39364
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 46934 39080 46940 39092
rect 46895 39052 46940 39080
rect 46934 39040 46940 39052
rect 46992 39040 46998 39092
rect 3510 38972 3516 39024
rect 3568 39012 3574 39024
rect 7558 39012 7564 39024
rect 3568 38984 7564 39012
rect 3568 38972 3574 38984
rect 7558 38972 7564 38984
rect 7616 38972 7622 39024
rect 46750 38904 46756 38956
rect 46808 38944 46814 38956
rect 46845 38947 46903 38953
rect 46845 38944 46857 38947
rect 46808 38916 46857 38944
rect 46808 38904 46814 38916
rect 46845 38913 46857 38916
rect 46891 38913 46903 38947
rect 47670 38944 47676 38956
rect 47631 38916 47676 38944
rect 46845 38907 46903 38913
rect 47670 38904 47676 38916
rect 47728 38904 47734 38956
rect 47854 38876 47860 38888
rect 47815 38848 47860 38876
rect 47854 38836 47860 38848
rect 47912 38836 47918 38888
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 26602 38536 26608 38548
rect 26563 38508 26608 38536
rect 26602 38496 26608 38508
rect 26660 38536 26666 38548
rect 26660 38508 27384 38536
rect 26660 38496 26666 38508
rect 22646 38332 22652 38344
rect 22607 38304 22652 38332
rect 22646 38292 22652 38304
rect 22704 38292 22710 38344
rect 27356 38341 27384 38508
rect 27522 38400 27528 38412
rect 27483 38372 27528 38400
rect 27522 38360 27528 38372
rect 27580 38360 27586 38412
rect 26329 38335 26387 38341
rect 26329 38301 26341 38335
rect 26375 38332 26387 38335
rect 27341 38335 27399 38341
rect 26375 38304 27016 38332
rect 26375 38301 26387 38304
rect 26329 38295 26387 38301
rect 22465 38199 22523 38205
rect 22465 38165 22477 38199
rect 22511 38196 22523 38199
rect 22830 38196 22836 38208
rect 22511 38168 22836 38196
rect 22511 38165 22523 38168
rect 22465 38159 22523 38165
rect 22830 38156 22836 38168
rect 22888 38156 22894 38208
rect 26142 38196 26148 38208
rect 26103 38168 26148 38196
rect 26142 38156 26148 38168
rect 26200 38156 26206 38208
rect 26988 38205 27016 38304
rect 27341 38301 27353 38335
rect 27387 38301 27399 38335
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 27341 38295 27399 38301
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 47670 38264 47676 38276
rect 46523 38236 47676 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 47670 38224 47676 38236
rect 47728 38224 47734 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 26973 38199 27031 38205
rect 26973 38165 26985 38199
rect 27019 38165 27031 38199
rect 26973 38159 27031 38165
rect 27430 38156 27436 38208
rect 27488 38196 27494 38208
rect 27488 38168 27533 38196
rect 27488 38156 27494 38168
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 47670 37992 47676 38004
rect 47631 37964 47676 37992
rect 47670 37952 47676 37964
rect 47728 37952 47734 38004
rect 22830 37924 22836 37936
rect 22791 37896 22836 37924
rect 22830 37884 22836 37896
rect 22888 37884 22894 37936
rect 23842 37884 23848 37936
rect 23900 37884 23906 37936
rect 26142 37884 26148 37936
rect 26200 37924 26206 37936
rect 27249 37927 27307 37933
rect 27249 37924 27261 37927
rect 26200 37896 27261 37924
rect 26200 37884 26206 37896
rect 27249 37893 27261 37896
rect 27295 37893 27307 37927
rect 27249 37887 27307 37893
rect 27982 37884 27988 37936
rect 28040 37884 28046 37936
rect 32214 37816 32220 37868
rect 32272 37856 32278 37868
rect 47581 37859 47639 37865
rect 47581 37856 47593 37859
rect 32272 37828 47593 37856
rect 32272 37816 32278 37828
rect 47581 37825 47593 37828
rect 47627 37825 47639 37859
rect 47581 37819 47639 37825
rect 22557 37791 22615 37797
rect 22557 37757 22569 37791
rect 22603 37788 22615 37791
rect 26973 37791 27031 37797
rect 22603 37760 22692 37788
rect 22603 37757 22615 37760
rect 22557 37751 22615 37757
rect 22664 37652 22692 37760
rect 26973 37757 26985 37791
rect 27019 37757 27031 37791
rect 26973 37751 27031 37757
rect 24210 37652 24216 37664
rect 22664 37624 24216 37652
rect 24210 37612 24216 37624
rect 24268 37612 24274 37664
rect 24302 37612 24308 37664
rect 24360 37652 24366 37664
rect 26988 37652 27016 37751
rect 27246 37748 27252 37800
rect 27304 37788 27310 37800
rect 28721 37791 28779 37797
rect 28721 37788 28733 37791
rect 27304 37760 28733 37788
rect 27304 37748 27310 37760
rect 28721 37757 28733 37760
rect 28767 37757 28779 37791
rect 28721 37751 28779 37757
rect 28534 37652 28540 37664
rect 24360 37624 24405 37652
rect 26988 37624 28540 37652
rect 24360 37612 24366 37624
rect 28534 37612 28540 37624
rect 28592 37612 28598 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 22281 37451 22339 37457
rect 22281 37417 22293 37451
rect 22327 37448 22339 37451
rect 22646 37448 22652 37460
rect 22327 37420 22652 37448
rect 22327 37417 22339 37420
rect 22281 37411 22339 37417
rect 22646 37408 22652 37420
rect 22704 37408 22710 37460
rect 23474 37408 23480 37460
rect 23532 37448 23538 37460
rect 24949 37451 25007 37457
rect 24949 37448 24961 37451
rect 23532 37420 24961 37448
rect 23532 37408 23538 37420
rect 24949 37417 24961 37420
rect 24995 37417 25007 37451
rect 24949 37411 25007 37417
rect 27341 37451 27399 37457
rect 27341 37417 27353 37451
rect 27387 37448 27399 37451
rect 27430 37448 27436 37460
rect 27387 37420 27436 37448
rect 27387 37417 27399 37420
rect 27341 37411 27399 37417
rect 27430 37408 27436 37420
rect 27488 37408 27494 37460
rect 46290 37408 46296 37460
rect 46348 37448 46354 37460
rect 47673 37451 47731 37457
rect 47673 37448 47685 37451
rect 46348 37420 47685 37448
rect 46348 37408 46354 37420
rect 47673 37417 47685 37420
rect 47719 37417 47731 37451
rect 47673 37411 47731 37417
rect 23382 37380 23388 37392
rect 22940 37352 23388 37380
rect 22940 37321 22968 37352
rect 23382 37340 23388 37352
rect 23440 37380 23446 37392
rect 27522 37380 27528 37392
rect 23440 37352 27528 37380
rect 23440 37340 23446 37352
rect 27522 37340 27528 37352
rect 27580 37340 27586 37392
rect 22925 37315 22983 37321
rect 22925 37281 22937 37315
rect 22971 37281 22983 37315
rect 24486 37312 24492 37324
rect 24447 37284 24492 37312
rect 22925 37275 22983 37281
rect 24486 37272 24492 37284
rect 24544 37272 24550 37324
rect 25222 37272 25228 37324
rect 25280 37312 25286 37324
rect 26973 37315 27031 37321
rect 26973 37312 26985 37315
rect 25280 37284 26985 37312
rect 25280 37272 25286 37284
rect 26973 37281 26985 37284
rect 27019 37281 27031 37315
rect 26973 37275 27031 37281
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37213 23719 37247
rect 23661 37207 23719 37213
rect 23753 37247 23811 37253
rect 23753 37213 23765 37247
rect 23799 37244 23811 37247
rect 23842 37244 23848 37256
rect 23799 37216 23848 37244
rect 23799 37213 23811 37216
rect 23753 37207 23811 37213
rect 11974 37136 11980 37188
rect 12032 37176 12038 37188
rect 22649 37179 22707 37185
rect 22649 37176 22661 37179
rect 12032 37148 22661 37176
rect 12032 37136 12038 37148
rect 22649 37145 22661 37148
rect 22695 37145 22707 37179
rect 22649 37139 22707 37145
rect 22741 37179 22799 37185
rect 22741 37145 22753 37179
rect 22787 37176 22799 37179
rect 23474 37176 23480 37188
rect 22787 37148 23480 37176
rect 22787 37145 22799 37148
rect 22741 37139 22799 37145
rect 23474 37136 23480 37148
rect 23532 37136 23538 37188
rect 23676 37108 23704 37207
rect 23842 37204 23848 37216
rect 23900 37204 23906 37256
rect 24302 37204 24308 37256
rect 24360 37244 24366 37256
rect 24578 37244 24584 37256
rect 24360 37216 24584 37244
rect 24360 37204 24366 37216
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25332 37216 25421 37244
rect 25332 37108 25360 37216
rect 25409 37213 25421 37216
rect 25455 37244 25467 37247
rect 25866 37244 25872 37256
rect 25455 37216 25872 37244
rect 25455 37213 25467 37216
rect 25409 37207 25467 37213
rect 25866 37204 25872 37216
rect 25924 37204 25930 37256
rect 27065 37247 27123 37253
rect 27065 37213 27077 37247
rect 27111 37244 27123 37247
rect 27246 37244 27252 37256
rect 27111 37216 27252 37244
rect 27111 37213 27123 37216
rect 27065 37207 27123 37213
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 27798 37204 27804 37256
rect 27856 37244 27862 37256
rect 27893 37247 27951 37253
rect 27893 37244 27905 37247
rect 27856 37216 27905 37244
rect 27856 37204 27862 37216
rect 27893 37213 27905 37216
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 27982 37204 27988 37256
rect 28040 37244 28046 37256
rect 28040 37216 28085 37244
rect 28040 37204 28046 37216
rect 25498 37108 25504 37120
rect 23676 37080 25360 37108
rect 25459 37080 25504 37108
rect 25498 37068 25504 37080
rect 25556 37068 25562 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 22554 36864 22560 36916
rect 22612 36904 22618 36916
rect 45554 36904 45560 36916
rect 22612 36876 45560 36904
rect 22612 36864 22618 36876
rect 45554 36864 45560 36876
rect 45612 36864 45618 36916
rect 25498 36796 25504 36848
rect 25556 36796 25562 36848
rect 29822 36796 29828 36848
rect 29880 36796 29886 36848
rect 28534 36768 28540 36780
rect 28495 36740 28540 36768
rect 28534 36728 28540 36740
rect 28592 36728 28598 36780
rect 24210 36660 24216 36712
rect 24268 36700 24274 36712
rect 24489 36703 24547 36709
rect 24489 36700 24501 36703
rect 24268 36672 24501 36700
rect 24268 36660 24274 36672
rect 24489 36669 24501 36672
rect 24535 36669 24547 36703
rect 24489 36663 24547 36669
rect 24765 36703 24823 36709
rect 24765 36669 24777 36703
rect 24811 36700 24823 36703
rect 26142 36700 26148 36712
rect 24811 36672 26148 36700
rect 24811 36669 24823 36672
rect 24765 36663 24823 36669
rect 26142 36660 26148 36672
rect 26200 36660 26206 36712
rect 28810 36700 28816 36712
rect 28771 36672 28816 36700
rect 28810 36660 28816 36672
rect 28868 36660 28874 36712
rect 28258 36632 28264 36644
rect 26160 36604 28264 36632
rect 25498 36524 25504 36576
rect 25556 36564 25562 36576
rect 26160 36564 26188 36604
rect 28258 36592 28264 36604
rect 28316 36592 28322 36644
rect 25556 36536 26188 36564
rect 26237 36567 26295 36573
rect 25556 36524 25562 36536
rect 26237 36533 26249 36567
rect 26283 36564 26295 36567
rect 26326 36564 26332 36576
rect 26283 36536 26332 36564
rect 26283 36533 26295 36536
rect 26237 36527 26295 36533
rect 26326 36524 26332 36536
rect 26384 36524 26390 36576
rect 30282 36564 30288 36576
rect 30243 36536 30288 36564
rect 30282 36524 30288 36536
rect 30340 36524 30346 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2038 36320 2044 36372
rect 2096 36360 2102 36372
rect 24486 36360 24492 36372
rect 2096 36332 6914 36360
rect 24447 36332 24492 36360
rect 2096 36320 2102 36332
rect 6886 36292 6914 36332
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 24578 36320 24584 36372
rect 24636 36360 24642 36372
rect 26142 36360 26148 36372
rect 24636 36332 26004 36360
rect 26103 36332 26148 36360
rect 24636 36320 24642 36332
rect 25976 36292 26004 36332
rect 26142 36320 26148 36332
rect 26200 36320 26206 36372
rect 28445 36363 28503 36369
rect 28445 36329 28457 36363
rect 28491 36360 28503 36363
rect 28718 36360 28724 36372
rect 28491 36332 28724 36360
rect 28491 36329 28503 36332
rect 28445 36323 28503 36329
rect 28718 36320 28724 36332
rect 28776 36320 28782 36372
rect 29733 36363 29791 36369
rect 29733 36329 29745 36363
rect 29779 36360 29791 36363
rect 29822 36360 29828 36372
rect 29779 36332 29828 36360
rect 29779 36329 29791 36332
rect 29733 36323 29791 36329
rect 29822 36320 29828 36332
rect 29880 36320 29886 36372
rect 26050 36292 26056 36304
rect 6886 36264 25820 36292
rect 25963 36264 26056 36292
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 21729 36227 21787 36233
rect 21729 36193 21741 36227
rect 21775 36224 21787 36227
rect 22554 36224 22560 36236
rect 21775 36196 22560 36224
rect 21775 36193 21787 36196
rect 21729 36187 21787 36193
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 22388 36165 22416 36196
rect 22554 36184 22560 36196
rect 22612 36184 22618 36236
rect 22649 36227 22707 36233
rect 22649 36193 22661 36227
rect 22695 36224 22707 36227
rect 23198 36224 23204 36236
rect 22695 36196 23204 36224
rect 22695 36193 22707 36196
rect 22649 36187 22707 36193
rect 23198 36184 23204 36196
rect 23256 36184 23262 36236
rect 25792 36233 25820 36264
rect 26050 36252 26056 36264
rect 26108 36292 26114 36304
rect 26108 36264 27108 36292
rect 26108 36252 26114 36264
rect 25777 36227 25835 36233
rect 25777 36193 25789 36227
rect 25823 36193 25835 36227
rect 26142 36224 26148 36236
rect 25777 36187 25835 36193
rect 25884 36196 26148 36224
rect 20993 36159 21051 36165
rect 20993 36125 21005 36159
rect 21039 36156 21051 36159
rect 22373 36159 22431 36165
rect 21039 36128 22048 36156
rect 21039 36125 21051 36128
rect 20993 36119 21051 36125
rect 1581 36091 1639 36097
rect 1581 36057 1593 36091
rect 1627 36088 1639 36091
rect 2222 36088 2228 36100
rect 1627 36060 2228 36088
rect 1627 36057 1639 36060
rect 1581 36051 1639 36057
rect 2222 36048 2228 36060
rect 2280 36048 2286 36100
rect 20806 36020 20812 36032
rect 20767 35992 20812 36020
rect 20806 35980 20812 35992
rect 20864 35980 20870 36032
rect 22020 36029 22048 36128
rect 22373 36125 22385 36159
rect 22419 36156 22431 36159
rect 24489 36159 24547 36165
rect 22419 36128 22453 36156
rect 22419 36125 22431 36128
rect 22373 36119 22431 36125
rect 24489 36125 24501 36159
rect 24535 36125 24547 36159
rect 24489 36119 24547 36125
rect 24673 36159 24731 36165
rect 24673 36125 24685 36159
rect 24719 36156 24731 36159
rect 25409 36159 25467 36165
rect 24719 36128 25360 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 24504 36088 24532 36119
rect 25038 36088 25044 36100
rect 24504 36060 25044 36088
rect 25038 36048 25044 36060
rect 25096 36048 25102 36100
rect 22005 36023 22063 36029
rect 22005 35989 22017 36023
rect 22051 35989 22063 36023
rect 22005 35983 22063 35989
rect 22462 35980 22468 36032
rect 22520 36020 22526 36032
rect 25332 36020 25360 36128
rect 25409 36125 25421 36159
rect 25455 36125 25467 36159
rect 25409 36119 25467 36125
rect 25424 36088 25452 36119
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 25593 36159 25651 36165
rect 25593 36156 25605 36159
rect 25556 36128 25605 36156
rect 25556 36116 25562 36128
rect 25593 36125 25605 36128
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 25685 36159 25743 36165
rect 25685 36125 25697 36159
rect 25731 36156 25743 36159
rect 25884 36156 25912 36196
rect 26142 36184 26148 36196
rect 26200 36184 26206 36236
rect 27080 36233 27108 36264
rect 27065 36227 27123 36233
rect 27065 36193 27077 36227
rect 27111 36193 27123 36227
rect 27065 36187 27123 36193
rect 25731 36128 25912 36156
rect 25731 36125 25743 36128
rect 25685 36119 25743 36125
rect 25958 36116 25964 36168
rect 26016 36156 26022 36168
rect 26016 36128 26061 36156
rect 26016 36116 26022 36128
rect 26326 36116 26332 36168
rect 26384 36156 26390 36168
rect 26789 36159 26847 36165
rect 26789 36156 26801 36159
rect 26384 36128 26801 36156
rect 26384 36116 26390 36128
rect 26789 36125 26801 36128
rect 26835 36125 26847 36159
rect 26789 36119 26847 36125
rect 26973 36159 27031 36165
rect 26973 36125 26985 36159
rect 27019 36125 27031 36159
rect 26973 36119 27031 36125
rect 28077 36159 28135 36165
rect 28077 36125 28089 36159
rect 28123 36156 28135 36159
rect 28166 36156 28172 36168
rect 28123 36128 28172 36156
rect 28123 36125 28135 36128
rect 28077 36119 28135 36125
rect 26234 36088 26240 36100
rect 25424 36060 26240 36088
rect 26234 36048 26240 36060
rect 26292 36048 26298 36100
rect 26988 36088 27016 36119
rect 28166 36116 28172 36128
rect 28224 36116 28230 36168
rect 28445 36159 28503 36165
rect 28445 36125 28457 36159
rect 28491 36156 28503 36159
rect 29270 36156 29276 36168
rect 28491 36128 29276 36156
rect 28491 36125 28503 36128
rect 28445 36119 28503 36125
rect 29270 36116 29276 36128
rect 29328 36116 29334 36168
rect 29641 36159 29699 36165
rect 29641 36125 29653 36159
rect 29687 36125 29699 36159
rect 29641 36119 29699 36125
rect 26344 36060 27016 36088
rect 26142 36020 26148 36032
rect 22520 35992 22565 36020
rect 25332 35992 26148 36020
rect 22520 35980 22526 35992
rect 26142 35980 26148 35992
rect 26200 36020 26206 36032
rect 26344 36020 26372 36060
rect 27798 36048 27804 36100
rect 27856 36088 27862 36100
rect 29656 36088 29684 36119
rect 27856 36060 29684 36088
rect 27856 36048 27862 36060
rect 26602 36020 26608 36032
rect 26200 35992 26372 36020
rect 26563 35992 26608 36020
rect 26200 35980 26206 35992
rect 26602 35980 26608 35992
rect 26660 35980 26666 36032
rect 28074 35980 28080 36032
rect 28132 36020 28138 36032
rect 28629 36023 28687 36029
rect 28629 36020 28641 36023
rect 28132 35992 28641 36020
rect 28132 35980 28138 35992
rect 28629 35989 28641 35992
rect 28675 35989 28687 36023
rect 29656 36020 29684 36060
rect 34514 36020 34520 36032
rect 29656 35992 34520 36020
rect 28629 35983 28687 35989
rect 34514 35980 34520 35992
rect 34572 35980 34578 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 25222 35816 25228 35828
rect 25183 35788 25228 35816
rect 25222 35776 25228 35788
rect 25280 35776 25286 35828
rect 26234 35816 26240 35828
rect 26195 35788 26240 35816
rect 26234 35776 26240 35788
rect 26292 35776 26298 35828
rect 27706 35816 27712 35828
rect 27172 35788 27712 35816
rect 27172 35760 27200 35788
rect 27706 35776 27712 35788
rect 27764 35776 27770 35828
rect 28810 35816 28816 35828
rect 28771 35788 28816 35816
rect 28810 35776 28816 35788
rect 28868 35776 28874 35828
rect 29270 35816 29276 35828
rect 29231 35788 29276 35816
rect 29270 35776 29276 35788
rect 29328 35776 29334 35828
rect 20254 35708 20260 35760
rect 20312 35708 20318 35760
rect 27154 35748 27160 35760
rect 27067 35720 27160 35748
rect 27154 35708 27160 35720
rect 27212 35708 27218 35760
rect 27246 35708 27252 35760
rect 27304 35708 27310 35760
rect 31481 35751 31539 35757
rect 28368 35720 29500 35748
rect 1394 35640 1400 35692
rect 1452 35680 1458 35692
rect 2041 35683 2099 35689
rect 2041 35680 2053 35683
rect 1452 35652 2053 35680
rect 1452 35640 1458 35652
rect 2041 35649 2053 35652
rect 2087 35649 2099 35683
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 2041 35643 2099 35649
rect 21284 35652 22017 35680
rect 19150 35572 19156 35624
rect 19208 35612 19214 35624
rect 19521 35615 19579 35621
rect 19521 35612 19533 35615
rect 19208 35584 19533 35612
rect 19208 35572 19214 35584
rect 19521 35581 19533 35584
rect 19567 35581 19579 35615
rect 19521 35575 19579 35581
rect 19797 35615 19855 35621
rect 19797 35581 19809 35615
rect 19843 35612 19855 35615
rect 20806 35612 20812 35624
rect 19843 35584 20812 35612
rect 19843 35581 19855 35584
rect 19797 35575 19855 35581
rect 20806 35572 20812 35584
rect 20864 35572 20870 35624
rect 21284 35621 21312 35652
rect 22005 35649 22017 35652
rect 22051 35680 22063 35683
rect 23106 35680 23112 35692
rect 22051 35652 23112 35680
rect 22051 35649 22063 35652
rect 22005 35643 22063 35649
rect 23106 35640 23112 35652
rect 23164 35640 23170 35692
rect 24854 35680 24860 35692
rect 24815 35652 24860 35680
rect 24854 35640 24860 35652
rect 24912 35640 24918 35692
rect 25682 35680 25688 35692
rect 25643 35652 25688 35680
rect 25682 35640 25688 35652
rect 25740 35640 25746 35692
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 26602 35680 26608 35692
rect 26099 35652 26608 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 26602 35640 26608 35652
rect 26660 35640 26666 35692
rect 27264 35680 27292 35708
rect 27433 35683 27491 35689
rect 27433 35680 27445 35683
rect 27264 35652 27445 35680
rect 27433 35649 27445 35652
rect 27479 35649 27491 35683
rect 28074 35680 28080 35692
rect 28035 35652 28080 35680
rect 27433 35643 27491 35649
rect 28074 35640 28080 35652
rect 28132 35640 28138 35692
rect 28258 35680 28264 35692
rect 28219 35652 28264 35680
rect 28258 35640 28264 35652
rect 28316 35640 28322 35692
rect 28368 35689 28396 35720
rect 28353 35683 28411 35689
rect 28353 35649 28365 35683
rect 28399 35649 28411 35683
rect 28626 35680 28632 35692
rect 28587 35652 28632 35680
rect 28353 35643 28411 35649
rect 21269 35615 21327 35621
rect 21269 35581 21281 35615
rect 21315 35581 21327 35615
rect 21269 35575 21327 35581
rect 21358 35572 21364 35624
rect 21416 35612 21422 35624
rect 21913 35615 21971 35621
rect 21913 35612 21925 35615
rect 21416 35584 21925 35612
rect 21416 35572 21422 35584
rect 21913 35581 21925 35584
rect 21959 35581 21971 35615
rect 21913 35575 21971 35581
rect 22373 35615 22431 35621
rect 22373 35581 22385 35615
rect 22419 35612 22431 35615
rect 22462 35612 22468 35624
rect 22419 35584 22468 35612
rect 22419 35581 22431 35584
rect 22373 35575 22431 35581
rect 22462 35572 22468 35584
rect 22520 35572 22526 35624
rect 23290 35572 23296 35624
rect 23348 35612 23354 35624
rect 24949 35615 25007 35621
rect 24949 35612 24961 35615
rect 23348 35584 24961 35612
rect 23348 35572 23354 35584
rect 24949 35581 24961 35584
rect 24995 35612 25007 35615
rect 25958 35612 25964 35624
rect 24995 35584 25964 35612
rect 24995 35581 25007 35584
rect 24949 35575 25007 35581
rect 25958 35572 25964 35584
rect 26016 35572 26022 35624
rect 27338 35612 27344 35624
rect 27251 35584 27344 35612
rect 27338 35572 27344 35584
rect 27396 35612 27402 35624
rect 28368 35612 28396 35643
rect 28626 35640 28632 35652
rect 28684 35640 28690 35692
rect 29472 35689 29500 35720
rect 31481 35717 31493 35751
rect 31527 35748 31539 35751
rect 31527 35720 32890 35748
rect 31527 35717 31539 35720
rect 31481 35711 31539 35717
rect 29457 35683 29515 35689
rect 29457 35649 29469 35683
rect 29503 35680 29515 35683
rect 30282 35680 30288 35692
rect 29503 35652 30288 35680
rect 29503 35649 29515 35652
rect 29457 35643 29515 35649
rect 30282 35640 30288 35652
rect 30340 35640 30346 35692
rect 31386 35680 31392 35692
rect 31347 35652 31392 35680
rect 31386 35640 31392 35652
rect 31444 35640 31450 35692
rect 27396 35584 28396 35612
rect 28445 35615 28503 35621
rect 27396 35572 27402 35584
rect 28445 35581 28457 35615
rect 28491 35581 28503 35615
rect 29733 35615 29791 35621
rect 29733 35612 29745 35615
rect 28445 35575 28503 35581
rect 28966 35584 29745 35612
rect 28460 35544 28488 35575
rect 28966 35544 28994 35584
rect 29733 35581 29745 35584
rect 29779 35612 29791 35615
rect 31202 35612 31208 35624
rect 29779 35584 31208 35612
rect 29779 35581 29791 35584
rect 29733 35575 29791 35581
rect 31202 35572 31208 35584
rect 31260 35572 31266 35624
rect 32122 35612 32128 35624
rect 32083 35584 32128 35612
rect 32122 35572 32128 35584
rect 32180 35572 32186 35624
rect 32401 35615 32459 35621
rect 32401 35581 32413 35615
rect 32447 35612 32459 35615
rect 32858 35612 32864 35624
rect 32447 35584 32864 35612
rect 32447 35581 32459 35584
rect 32401 35575 32459 35581
rect 32858 35572 32864 35584
rect 32916 35572 32922 35624
rect 20824 35516 28488 35544
rect 28552 35516 28994 35544
rect 19886 35436 19892 35488
rect 19944 35476 19950 35488
rect 20824 35476 20852 35516
rect 25038 35476 25044 35488
rect 19944 35448 20852 35476
rect 24951 35448 25044 35476
rect 19944 35436 19950 35448
rect 25038 35436 25044 35448
rect 25096 35476 25102 35488
rect 25406 35476 25412 35488
rect 25096 35448 25412 35476
rect 25096 35436 25102 35448
rect 25406 35436 25412 35448
rect 25464 35436 25470 35488
rect 25774 35476 25780 35488
rect 25735 35448 25780 35476
rect 25774 35436 25780 35448
rect 25832 35436 25838 35488
rect 25958 35436 25964 35488
rect 26016 35476 26022 35488
rect 27157 35479 27215 35485
rect 27157 35476 27169 35479
rect 26016 35448 27169 35476
rect 26016 35436 26022 35448
rect 27157 35445 27169 35448
rect 27203 35445 27215 35479
rect 27157 35439 27215 35445
rect 27246 35436 27252 35488
rect 27304 35476 27310 35488
rect 27617 35479 27675 35485
rect 27617 35476 27629 35479
rect 27304 35448 27629 35476
rect 27304 35436 27310 35448
rect 27617 35445 27629 35448
rect 27663 35445 27675 35479
rect 27617 35439 27675 35445
rect 27706 35436 27712 35488
rect 27764 35476 27770 35488
rect 28552 35476 28580 35516
rect 27764 35448 28580 35476
rect 27764 35436 27770 35448
rect 28626 35436 28632 35488
rect 28684 35476 28690 35488
rect 29641 35479 29699 35485
rect 29641 35476 29653 35479
rect 28684 35448 29653 35476
rect 28684 35436 28690 35448
rect 29641 35445 29653 35448
rect 29687 35476 29699 35479
rect 31938 35476 31944 35488
rect 29687 35448 31944 35476
rect 29687 35445 29699 35448
rect 29641 35439 29699 35445
rect 31938 35436 31944 35448
rect 31996 35436 32002 35488
rect 33134 35436 33140 35488
rect 33192 35476 33198 35488
rect 33873 35479 33931 35485
rect 33873 35476 33885 35479
rect 33192 35448 33885 35476
rect 33192 35436 33198 35448
rect 33873 35445 33885 35448
rect 33919 35445 33931 35479
rect 33873 35439 33931 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 19886 35272 19892 35284
rect 6886 35244 19892 35272
rect 2038 35164 2044 35216
rect 2096 35204 2102 35216
rect 6886 35204 6914 35244
rect 19886 35232 19892 35244
rect 19944 35232 19950 35284
rect 19981 35275 20039 35281
rect 19981 35241 19993 35275
rect 20027 35272 20039 35275
rect 20254 35272 20260 35284
rect 20027 35244 20260 35272
rect 20027 35241 20039 35244
rect 19981 35235 20039 35241
rect 20254 35232 20260 35244
rect 20312 35232 20318 35284
rect 28169 35275 28227 35281
rect 28169 35241 28181 35275
rect 28215 35272 28227 35275
rect 28350 35272 28356 35284
rect 28215 35244 28356 35272
rect 28215 35241 28227 35244
rect 28169 35235 28227 35241
rect 28350 35232 28356 35244
rect 28408 35232 28414 35284
rect 32858 35272 32864 35284
rect 32819 35244 32864 35272
rect 32858 35232 32864 35244
rect 32916 35232 32922 35284
rect 2096 35176 6914 35204
rect 2096 35164 2102 35176
rect 25682 35164 25688 35216
rect 25740 35204 25746 35216
rect 27614 35204 27620 35216
rect 25740 35176 27620 35204
rect 25740 35164 25746 35176
rect 27614 35164 27620 35176
rect 27672 35204 27678 35216
rect 32122 35204 32128 35216
rect 27672 35176 28120 35204
rect 27672 35164 27678 35176
rect 23385 35139 23443 35145
rect 23385 35105 23397 35139
rect 23431 35136 23443 35139
rect 24854 35136 24860 35148
rect 23431 35108 24860 35136
rect 23431 35105 23443 35108
rect 23385 35099 23443 35105
rect 24854 35096 24860 35108
rect 24912 35136 24918 35148
rect 27433 35139 27491 35145
rect 24912 35108 26188 35136
rect 24912 35096 24918 35108
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 2130 35068 2136 35080
rect 2091 35040 2136 35068
rect 2130 35028 2136 35040
rect 2188 35028 2194 35080
rect 19242 35028 19248 35080
rect 19300 35068 19306 35080
rect 19889 35071 19947 35077
rect 19889 35068 19901 35071
rect 19300 35040 19901 35068
rect 19300 35028 19306 35040
rect 19889 35037 19901 35040
rect 19935 35037 19947 35071
rect 23290 35068 23296 35080
rect 23251 35040 23296 35068
rect 19889 35031 19947 35037
rect 23290 35028 23296 35040
rect 23348 35028 23354 35080
rect 23934 35028 23940 35080
rect 23992 35068 23998 35080
rect 24397 35071 24455 35077
rect 24397 35068 24409 35071
rect 23992 35040 24409 35068
rect 23992 35028 23998 35040
rect 24397 35037 24409 35040
rect 24443 35068 24455 35071
rect 25774 35068 25780 35080
rect 24443 35040 25780 35068
rect 24443 35037 24455 35040
rect 24397 35031 24455 35037
rect 25774 35028 25780 35040
rect 25832 35028 25838 35080
rect 26050 35068 26056 35080
rect 26011 35040 26056 35068
rect 26050 35028 26056 35040
rect 26108 35028 26114 35080
rect 26160 35000 26188 35108
rect 27433 35105 27445 35139
rect 27479 35136 27491 35139
rect 27985 35139 28043 35145
rect 27985 35136 27997 35139
rect 27479 35108 27997 35136
rect 27479 35105 27491 35108
rect 27433 35099 27491 35105
rect 27985 35105 27997 35108
rect 28031 35105 28043 35139
rect 27985 35099 28043 35105
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35068 26295 35071
rect 26326 35068 26332 35080
rect 26283 35040 26332 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 27065 35071 27123 35077
rect 27065 35037 27077 35071
rect 27111 35068 27123 35071
rect 27154 35068 27160 35080
rect 27111 35040 27160 35068
rect 27111 35037 27123 35040
rect 27065 35031 27123 35037
rect 27154 35028 27160 35040
rect 27212 35028 27218 35080
rect 27249 35071 27307 35077
rect 27249 35037 27261 35071
rect 27295 35068 27307 35071
rect 27338 35068 27344 35080
rect 27295 35040 27344 35068
rect 27295 35037 27307 35040
rect 27249 35031 27307 35037
rect 27338 35028 27344 35040
rect 27396 35028 27402 35080
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35068 27951 35071
rect 28092 35068 28120 35176
rect 31726 35176 32128 35204
rect 28534 35096 28540 35148
rect 28592 35136 28598 35148
rect 29641 35139 29699 35145
rect 29641 35136 29653 35139
rect 28592 35108 29653 35136
rect 28592 35096 28598 35108
rect 29641 35105 29653 35108
rect 29687 35136 29699 35139
rect 31726 35136 31754 35176
rect 32122 35164 32128 35176
rect 32180 35204 32186 35216
rect 32950 35204 32956 35216
rect 32180 35176 32956 35204
rect 32180 35164 32186 35176
rect 32950 35164 32956 35176
rect 33008 35164 33014 35216
rect 34514 35164 34520 35216
rect 34572 35204 34578 35216
rect 34572 35176 35664 35204
rect 34572 35164 34578 35176
rect 31938 35136 31944 35148
rect 29687 35108 31754 35136
rect 31899 35108 31944 35136
rect 29687 35105 29699 35108
rect 29641 35099 29699 35105
rect 31938 35096 31944 35108
rect 31996 35096 32002 35148
rect 32766 35096 32772 35148
rect 32824 35136 32830 35148
rect 33321 35139 33379 35145
rect 33321 35136 33333 35139
rect 32824 35108 33333 35136
rect 32824 35096 32830 35108
rect 33321 35105 33333 35108
rect 33367 35136 33379 35139
rect 35069 35139 35127 35145
rect 33367 35108 35020 35136
rect 33367 35105 33379 35108
rect 33321 35099 33379 35105
rect 27939 35040 28120 35068
rect 28169 35071 28227 35077
rect 27939 35037 27951 35040
rect 27893 35031 27951 35037
rect 28169 35037 28181 35071
rect 28215 35037 28227 35071
rect 28169 35031 28227 35037
rect 26160 34972 27384 35000
rect 1397 34935 1455 34941
rect 1397 34901 1409 34935
rect 1443 34932 1455 34935
rect 1486 34932 1492 34944
rect 1443 34904 1492 34932
rect 1443 34901 1455 34904
rect 1397 34895 1455 34901
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 23474 34892 23480 34944
rect 23532 34932 23538 34944
rect 23661 34935 23719 34941
rect 23661 34932 23673 34935
rect 23532 34904 23673 34932
rect 23532 34892 23538 34904
rect 23661 34901 23673 34904
rect 23707 34901 23719 34935
rect 23661 34895 23719 34901
rect 24581 34935 24639 34941
rect 24581 34901 24593 34935
rect 24627 34932 24639 34935
rect 24762 34932 24768 34944
rect 24627 34904 24768 34932
rect 24627 34901 24639 34904
rect 24581 34895 24639 34901
rect 24762 34892 24768 34904
rect 24820 34892 24826 34944
rect 26421 34935 26479 34941
rect 26421 34901 26433 34935
rect 26467 34932 26479 34935
rect 26786 34932 26792 34944
rect 26467 34904 26792 34932
rect 26467 34901 26479 34904
rect 26421 34895 26479 34901
rect 26786 34892 26792 34904
rect 26844 34892 26850 34944
rect 27356 34932 27384 34972
rect 27706 34960 27712 35012
rect 27764 35000 27770 35012
rect 28184 35000 28212 35031
rect 31202 35028 31208 35080
rect 31260 35068 31266 35080
rect 32033 35071 32091 35077
rect 32033 35068 32045 35071
rect 31260 35040 32045 35068
rect 31260 35028 31266 35040
rect 32033 35037 32045 35040
rect 32079 35037 32091 35071
rect 32033 35031 32091 35037
rect 29914 35000 29920 35012
rect 27764 34972 28212 35000
rect 29875 34972 29920 35000
rect 27764 34960 27770 34972
rect 29914 34960 29920 34972
rect 29972 34960 29978 35012
rect 30926 34960 30932 35012
rect 30984 34960 30990 35012
rect 32048 35000 32076 35031
rect 32858 35028 32864 35080
rect 32916 35068 32922 35080
rect 33045 35071 33103 35077
rect 33045 35068 33057 35071
rect 32916 35040 33057 35068
rect 32916 35028 32922 35040
rect 33045 35037 33057 35040
rect 33091 35037 33103 35071
rect 33045 35031 33103 35037
rect 33229 35071 33287 35077
rect 33229 35037 33241 35071
rect 33275 35037 33287 35071
rect 33229 35031 33287 35037
rect 34885 35071 34943 35077
rect 34885 35037 34897 35071
rect 34931 35037 34943 35071
rect 34992 35068 35020 35108
rect 35069 35105 35081 35139
rect 35115 35136 35127 35139
rect 35342 35136 35348 35148
rect 35115 35108 35348 35136
rect 35115 35105 35127 35108
rect 35069 35099 35127 35105
rect 35342 35096 35348 35108
rect 35400 35096 35406 35148
rect 35161 35071 35219 35077
rect 35161 35068 35173 35071
rect 34992 35040 35173 35068
rect 34885 35031 34943 35037
rect 35161 35037 35173 35040
rect 35207 35068 35219 35071
rect 35434 35068 35440 35080
rect 35207 35040 35440 35068
rect 35207 35037 35219 35040
rect 35161 35031 35219 35037
rect 33134 35000 33140 35012
rect 32048 34972 33140 35000
rect 33134 34960 33140 34972
rect 33192 34960 33198 35012
rect 28166 34932 28172 34944
rect 27356 34904 28172 34932
rect 28166 34892 28172 34904
rect 28224 34932 28230 34944
rect 28353 34935 28411 34941
rect 28353 34932 28365 34935
rect 28224 34904 28365 34932
rect 28224 34892 28230 34904
rect 28353 34901 28365 34904
rect 28399 34901 28411 34935
rect 28353 34895 28411 34901
rect 28534 34892 28540 34944
rect 28592 34932 28598 34944
rect 31389 34935 31447 34941
rect 31389 34932 31401 34935
rect 28592 34904 31401 34932
rect 28592 34892 28598 34904
rect 31389 34901 31401 34904
rect 31435 34901 31447 34935
rect 31389 34895 31447 34901
rect 32401 34935 32459 34941
rect 32401 34901 32413 34935
rect 32447 34932 32459 34935
rect 33244 34932 33272 35031
rect 34900 35000 34928 35031
rect 35434 35028 35440 35040
rect 35492 35028 35498 35080
rect 35636 35077 35664 35176
rect 35621 35071 35679 35077
rect 35621 35037 35633 35071
rect 35667 35068 35679 35071
rect 35802 35068 35808 35080
rect 35667 35040 35808 35068
rect 35667 35037 35679 35040
rect 35621 35031 35679 35037
rect 35802 35028 35808 35040
rect 35860 35028 35866 35080
rect 47302 35068 47308 35080
rect 47263 35040 47308 35068
rect 47302 35028 47308 35040
rect 47360 35028 47366 35080
rect 47486 35028 47492 35080
rect 47544 35068 47550 35080
rect 47581 35071 47639 35077
rect 47581 35068 47593 35071
rect 47544 35040 47593 35068
rect 47544 35028 47550 35040
rect 47581 35037 47593 35040
rect 47627 35037 47639 35071
rect 47581 35031 47639 35037
rect 35526 35000 35532 35012
rect 34900 34972 35532 35000
rect 35526 34960 35532 34972
rect 35584 34960 35590 35012
rect 32447 34904 33272 34932
rect 32447 34901 32459 34904
rect 32401 34895 32459 34901
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 34701 34935 34759 34941
rect 34701 34932 34713 34935
rect 34572 34904 34713 34932
rect 34572 34892 34578 34904
rect 34701 34901 34713 34904
rect 34747 34901 34759 34935
rect 35710 34932 35716 34944
rect 35671 34904 35716 34932
rect 34701 34895 34759 34901
rect 35710 34892 35716 34904
rect 35768 34892 35774 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 25958 34728 25964 34740
rect 25919 34700 25964 34728
rect 25958 34688 25964 34700
rect 26016 34688 26022 34740
rect 26142 34688 26148 34740
rect 26200 34728 26206 34740
rect 27709 34731 27767 34737
rect 27709 34728 27721 34731
rect 26200 34700 27721 34728
rect 26200 34688 26206 34700
rect 27709 34697 27721 34700
rect 27755 34697 27767 34731
rect 29549 34731 29607 34737
rect 27709 34691 27767 34697
rect 28184 34700 29500 34728
rect 23290 34660 23296 34672
rect 23251 34632 23296 34660
rect 23290 34620 23296 34632
rect 23348 34620 23354 34672
rect 23509 34663 23567 34669
rect 23509 34629 23521 34663
rect 23555 34660 23567 34663
rect 23658 34660 23664 34672
rect 23555 34632 23664 34660
rect 23555 34629 23567 34632
rect 23509 34623 23567 34629
rect 23658 34620 23664 34632
rect 23716 34620 23722 34672
rect 25774 34660 25780 34672
rect 25714 34632 25780 34660
rect 25774 34620 25780 34632
rect 25832 34620 25838 34672
rect 27246 34660 27252 34672
rect 27207 34632 27252 34660
rect 27246 34620 27252 34632
rect 27304 34620 27310 34672
rect 28184 34660 28212 34700
rect 28534 34660 28540 34672
rect 27448 34632 28212 34660
rect 28276 34632 28540 34660
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34592 18843 34595
rect 19978 34592 19984 34604
rect 18831 34564 19984 34592
rect 18831 34561 18843 34564
rect 18785 34555 18843 34561
rect 19978 34552 19984 34564
rect 20036 34552 20042 34604
rect 25866 34552 25872 34604
rect 25924 34592 25930 34604
rect 27448 34592 27476 34632
rect 25924 34564 27476 34592
rect 27525 34595 27583 34601
rect 25924 34552 25930 34564
rect 27525 34561 27537 34595
rect 27571 34592 27583 34595
rect 27706 34592 27712 34604
rect 27571 34564 27712 34592
rect 27571 34561 27583 34564
rect 27525 34555 27583 34561
rect 27706 34552 27712 34564
rect 27764 34552 27770 34604
rect 28276 34601 28304 34632
rect 28534 34620 28540 34632
rect 28592 34620 28598 34672
rect 29472 34660 29500 34700
rect 29549 34697 29561 34731
rect 29595 34728 29607 34731
rect 29914 34728 29920 34740
rect 29595 34700 29920 34728
rect 29595 34697 29607 34700
rect 29549 34691 29607 34697
rect 29914 34688 29920 34700
rect 29972 34688 29978 34740
rect 30926 34728 30932 34740
rect 30887 34700 30932 34728
rect 30926 34688 30932 34700
rect 30984 34688 30990 34740
rect 32858 34728 32864 34740
rect 32819 34700 32864 34728
rect 32858 34688 32864 34700
rect 32916 34688 32922 34740
rect 36262 34728 36268 34740
rect 33520 34700 36268 34728
rect 31386 34660 31392 34672
rect 29472 34632 31392 34660
rect 28261 34595 28319 34601
rect 28261 34561 28273 34595
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 24210 34524 24216 34536
rect 24171 34496 24216 34524
rect 24210 34484 24216 34496
rect 24268 34484 24274 34536
rect 26786 34484 26792 34536
rect 26844 34524 26850 34536
rect 27341 34527 27399 34533
rect 27341 34524 27353 34527
rect 26844 34496 27353 34524
rect 26844 34484 26850 34496
rect 27341 34493 27353 34496
rect 27387 34493 27399 34527
rect 27341 34487 27399 34493
rect 28276 34456 28304 34555
rect 28442 34552 28448 34604
rect 28500 34592 28506 34604
rect 30852 34601 30880 34632
rect 31386 34620 31392 34632
rect 31444 34620 31450 34672
rect 29733 34595 29791 34601
rect 29733 34592 29745 34595
rect 28500 34564 29745 34592
rect 28500 34552 28506 34564
rect 29733 34561 29745 34564
rect 29779 34561 29791 34595
rect 29733 34555 29791 34561
rect 30837 34595 30895 34601
rect 30837 34561 30849 34595
rect 30883 34561 30895 34595
rect 33042 34592 33048 34604
rect 30837 34555 30895 34561
rect 31726 34564 33048 34592
rect 28350 34484 28356 34536
rect 28408 34524 28414 34536
rect 28537 34527 28595 34533
rect 28537 34524 28549 34527
rect 28408 34496 28549 34524
rect 28408 34484 28414 34496
rect 28537 34493 28549 34496
rect 28583 34493 28595 34527
rect 28537 34487 28595 34493
rect 29822 34484 29828 34536
rect 29880 34524 29886 34536
rect 30009 34527 30067 34533
rect 30009 34524 30021 34527
rect 29880 34496 30021 34524
rect 29880 34484 29886 34496
rect 30009 34493 30021 34496
rect 30055 34493 30067 34527
rect 30009 34487 30067 34493
rect 30466 34484 30472 34536
rect 30524 34524 30530 34536
rect 31726 34524 31754 34564
rect 33042 34552 33048 34564
rect 33100 34552 33106 34604
rect 33134 34552 33140 34604
rect 33192 34592 33198 34604
rect 33192 34564 33237 34592
rect 33192 34552 33198 34564
rect 33410 34552 33416 34604
rect 33468 34592 33474 34604
rect 33520 34592 33548 34700
rect 36262 34688 36268 34700
rect 36320 34688 36326 34740
rect 34241 34663 34299 34669
rect 34241 34629 34253 34663
rect 34287 34660 34299 34663
rect 34514 34660 34520 34672
rect 34287 34632 34520 34660
rect 34287 34629 34299 34632
rect 34241 34623 34299 34629
rect 34514 34620 34520 34632
rect 34572 34620 34578 34672
rect 35710 34660 35716 34672
rect 35466 34632 35716 34660
rect 35710 34620 35716 34632
rect 35768 34620 35774 34672
rect 48130 34592 48136 34604
rect 33468 34564 33561 34592
rect 48091 34564 48136 34592
rect 33468 34552 33474 34564
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 30524 34496 31754 34524
rect 30524 34484 30530 34496
rect 32950 34484 32956 34536
rect 33008 34524 33014 34536
rect 33965 34527 34023 34533
rect 33965 34524 33977 34527
rect 33008 34496 33977 34524
rect 33008 34484 33014 34496
rect 33965 34493 33977 34496
rect 34011 34493 34023 34527
rect 33965 34487 34023 34493
rect 33318 34456 33324 34468
rect 27540 34428 28304 34456
rect 33279 34428 33324 34456
rect 18969 34391 19027 34397
rect 18969 34357 18981 34391
rect 19015 34388 19027 34391
rect 19242 34388 19248 34400
rect 19015 34360 19248 34388
rect 19015 34357 19027 34360
rect 18969 34351 19027 34357
rect 19242 34348 19248 34360
rect 19300 34348 19306 34400
rect 23014 34348 23020 34400
rect 23072 34388 23078 34400
rect 23382 34388 23388 34400
rect 23072 34360 23388 34388
rect 23072 34348 23078 34360
rect 23382 34348 23388 34360
rect 23440 34388 23446 34400
rect 23477 34391 23535 34397
rect 23477 34388 23489 34391
rect 23440 34360 23489 34388
rect 23440 34348 23446 34360
rect 23477 34357 23489 34360
rect 23523 34357 23535 34391
rect 23477 34351 23535 34357
rect 23566 34348 23572 34400
rect 23624 34388 23630 34400
rect 23661 34391 23719 34397
rect 23661 34388 23673 34391
rect 23624 34360 23673 34388
rect 23624 34348 23630 34360
rect 23661 34357 23673 34360
rect 23707 34357 23719 34391
rect 23661 34351 23719 34357
rect 23842 34348 23848 34400
rect 23900 34388 23906 34400
rect 27540 34397 27568 34428
rect 33318 34416 33324 34428
rect 33376 34416 33382 34468
rect 24470 34391 24528 34397
rect 24470 34388 24482 34391
rect 23900 34360 24482 34388
rect 23900 34348 23906 34360
rect 24470 34357 24482 34360
rect 24516 34357 24528 34391
rect 24470 34351 24528 34357
rect 27525 34391 27583 34397
rect 27525 34357 27537 34391
rect 27571 34357 27583 34391
rect 29914 34388 29920 34400
rect 29875 34360 29920 34388
rect 27525 34351 27583 34357
rect 29914 34348 29920 34360
rect 29972 34348 29978 34400
rect 35710 34388 35716 34400
rect 35671 34360 35716 34388
rect 35710 34348 35716 34360
rect 35768 34348 35774 34400
rect 47946 34388 47952 34400
rect 47907 34360 47952 34388
rect 47946 34348 47952 34360
rect 48004 34348 48010 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 14642 34144 14648 34196
rect 14700 34184 14706 34196
rect 14700 34156 22237 34184
rect 14700 34144 14706 34156
rect 20346 34076 20352 34128
rect 20404 34116 20410 34128
rect 21082 34116 21088 34128
rect 20404 34088 21088 34116
rect 20404 34076 20410 34088
rect 21082 34076 21088 34088
rect 21140 34076 21146 34128
rect 21560 34020 22140 34048
rect 19242 33940 19248 33992
rect 19300 33980 19306 33992
rect 19337 33983 19395 33989
rect 19337 33980 19349 33983
rect 19300 33952 19349 33980
rect 19300 33940 19306 33952
rect 19337 33949 19349 33952
rect 19383 33949 19395 33983
rect 19337 33943 19395 33949
rect 20625 33983 20683 33989
rect 20625 33949 20637 33983
rect 20671 33949 20683 33983
rect 20625 33943 20683 33949
rect 19426 33844 19432 33856
rect 19387 33816 19432 33844
rect 19426 33804 19432 33816
rect 19484 33804 19490 33856
rect 20640 33844 20668 33943
rect 20714 33940 20720 33992
rect 20772 33980 20778 33992
rect 20772 33952 20817 33980
rect 20772 33940 20778 33952
rect 20898 33940 20904 33992
rect 20956 33980 20962 33992
rect 20956 33952 21001 33980
rect 20956 33940 20962 33952
rect 21082 33940 21088 33992
rect 21140 33989 21146 33992
rect 21140 33980 21148 33989
rect 21140 33952 21185 33980
rect 21140 33943 21148 33952
rect 21140 33940 21146 33943
rect 20993 33915 21051 33921
rect 20993 33881 21005 33915
rect 21039 33912 21051 33915
rect 21560 33912 21588 34020
rect 21910 33989 21916 33992
rect 21729 33983 21787 33989
rect 21729 33980 21741 33983
rect 21039 33884 21588 33912
rect 21652 33952 21741 33980
rect 21039 33881 21051 33884
rect 20993 33875 21051 33881
rect 20898 33844 20904 33856
rect 20640 33816 20904 33844
rect 20898 33804 20904 33816
rect 20956 33804 20962 33856
rect 21266 33844 21272 33856
rect 21227 33816 21272 33844
rect 21266 33804 21272 33816
rect 21324 33804 21330 33856
rect 21652 33844 21680 33952
rect 21729 33949 21741 33952
rect 21775 33949 21787 33983
rect 21729 33943 21787 33949
rect 21877 33983 21916 33989
rect 21877 33949 21889 33983
rect 21877 33943 21916 33949
rect 21910 33940 21916 33943
rect 21968 33940 21974 33992
rect 22002 33912 22008 33924
rect 21963 33884 22008 33912
rect 22002 33872 22008 33884
rect 22060 33872 22066 33924
rect 22112 33921 22140 34020
rect 22209 33989 22237 34156
rect 22370 34144 22376 34196
rect 22428 34184 22434 34196
rect 22428 34156 22473 34184
rect 22428 34144 22434 34156
rect 23290 34144 23296 34196
rect 23348 34184 23354 34196
rect 25774 34184 25780 34196
rect 23348 34156 23796 34184
rect 25735 34156 25780 34184
rect 23348 34144 23354 34156
rect 23566 34116 23572 34128
rect 23124 34088 23572 34116
rect 22194 33983 22252 33989
rect 22194 33949 22206 33983
rect 22240 33949 22252 33983
rect 23124 33980 23152 34088
rect 23566 34076 23572 34088
rect 23624 34076 23630 34128
rect 23768 34116 23796 34156
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 35161 34187 35219 34193
rect 25884 34156 31754 34184
rect 25884 34116 25912 34156
rect 23768 34088 25912 34116
rect 27157 34119 27215 34125
rect 27157 34085 27169 34119
rect 27203 34116 27215 34119
rect 27614 34116 27620 34128
rect 27203 34088 27620 34116
rect 27203 34085 27215 34088
rect 27157 34079 27215 34085
rect 27614 34076 27620 34088
rect 27672 34116 27678 34128
rect 28997 34119 29055 34125
rect 27672 34088 28580 34116
rect 27672 34076 27678 34088
rect 24026 34048 24032 34060
rect 23492 34020 24032 34048
rect 23382 33989 23388 33992
rect 23201 33983 23259 33989
rect 23201 33980 23213 33983
rect 23124 33952 23213 33980
rect 22194 33943 22252 33949
rect 23201 33949 23213 33952
rect 23247 33949 23259 33983
rect 23201 33943 23259 33949
rect 23349 33983 23388 33989
rect 23349 33949 23361 33983
rect 23349 33943 23388 33949
rect 23382 33940 23388 33943
rect 23440 33940 23446 33992
rect 23492 33989 23520 34020
rect 24026 34008 24032 34020
rect 24084 34048 24090 34060
rect 24946 34048 24952 34060
rect 24084 34020 24952 34048
rect 24084 34008 24090 34020
rect 24946 34008 24952 34020
rect 25004 34008 25010 34060
rect 27798 34048 27804 34060
rect 26252 34020 27804 34048
rect 26252 33992 26280 34020
rect 27798 34008 27804 34020
rect 27856 34008 27862 34060
rect 28552 34057 28580 34088
rect 28997 34085 29009 34119
rect 29043 34116 29055 34119
rect 29914 34116 29920 34128
rect 29043 34088 29920 34116
rect 29043 34085 29055 34088
rect 28997 34079 29055 34085
rect 29914 34076 29920 34088
rect 29972 34076 29978 34128
rect 31726 34116 31754 34156
rect 35161 34153 35173 34187
rect 35207 34184 35219 34187
rect 35342 34184 35348 34196
rect 35207 34156 35348 34184
rect 35207 34153 35219 34156
rect 35161 34147 35219 34153
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 35526 34144 35532 34196
rect 35584 34184 35590 34196
rect 35713 34187 35771 34193
rect 35713 34184 35725 34187
rect 35584 34156 35725 34184
rect 35584 34144 35590 34156
rect 35713 34153 35725 34156
rect 35759 34153 35771 34187
rect 35713 34147 35771 34153
rect 47854 34116 47860 34128
rect 31726 34088 47860 34116
rect 47854 34076 47860 34088
rect 47912 34076 47918 34128
rect 28537 34051 28595 34057
rect 28537 34017 28549 34051
rect 28583 34017 28595 34051
rect 34790 34048 34796 34060
rect 34751 34020 34796 34048
rect 28537 34011 28595 34017
rect 34790 34008 34796 34020
rect 34848 34008 34854 34060
rect 35710 34048 35716 34060
rect 34900 34020 35716 34048
rect 23477 33983 23535 33989
rect 23477 33949 23489 33983
rect 23523 33949 23535 33983
rect 23477 33943 23535 33949
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23707 33983 23765 33989
rect 23707 33949 23719 33983
rect 23753 33980 23765 33983
rect 24486 33980 24492 33992
rect 23753 33952 24492 33980
rect 23753 33949 23765 33952
rect 23707 33943 23765 33949
rect 22097 33915 22155 33921
rect 22097 33881 22109 33915
rect 22143 33912 22155 33915
rect 23592 33912 23620 33943
rect 24486 33940 24492 33952
rect 24544 33940 24550 33992
rect 25685 33983 25743 33989
rect 25685 33949 25697 33983
rect 25731 33980 25743 33983
rect 26234 33980 26240 33992
rect 25731 33952 26240 33980
rect 25731 33949 25743 33952
rect 25685 33943 25743 33949
rect 26234 33940 26240 33952
rect 26292 33940 26298 33992
rect 26786 33980 26792 33992
rect 26747 33952 26792 33980
rect 26786 33940 26792 33952
rect 26844 33940 26850 33992
rect 28350 33940 28356 33992
rect 28408 33980 28414 33992
rect 28629 33983 28687 33989
rect 28629 33980 28641 33983
rect 28408 33952 28641 33980
rect 28408 33940 28414 33952
rect 28629 33949 28641 33952
rect 28675 33949 28687 33983
rect 28629 33943 28687 33949
rect 34514 33940 34520 33992
rect 34572 33980 34578 33992
rect 34900 33989 34928 34020
rect 35710 34008 35716 34020
rect 35768 34048 35774 34060
rect 36170 34048 36176 34060
rect 35768 34020 36032 34048
rect 36131 34020 36176 34048
rect 35768 34008 35774 34020
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34572 33952 34897 33980
rect 34572 33940 34578 33952
rect 34885 33949 34897 33952
rect 34931 33949 34943 33983
rect 35894 33980 35900 33992
rect 35855 33952 35900 33980
rect 34885 33943 34943 33949
rect 35894 33940 35900 33952
rect 35952 33940 35958 33992
rect 36004 33989 36032 34020
rect 36170 34008 36176 34020
rect 36228 34008 36234 34060
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34048 46351 34051
rect 47946 34048 47952 34060
rect 46339 34020 47952 34048
rect 46339 34017 46351 34020
rect 46293 34011 46351 34017
rect 47946 34008 47952 34020
rect 48004 34008 48010 34060
rect 35989 33983 36047 33989
rect 35989 33949 36001 33983
rect 36035 33949 36047 33983
rect 36262 33980 36268 33992
rect 36223 33952 36268 33980
rect 35989 33943 36047 33949
rect 36262 33940 36268 33952
rect 36320 33940 36326 33992
rect 24302 33912 24308 33924
rect 22143 33884 24308 33912
rect 22143 33881 22155 33884
rect 22097 33875 22155 33881
rect 24302 33872 24308 33884
rect 24360 33872 24366 33924
rect 24854 33872 24860 33924
rect 24912 33912 24918 33924
rect 26973 33915 27031 33921
rect 26973 33912 26985 33915
rect 24912 33884 26985 33912
rect 24912 33872 24918 33884
rect 26973 33881 26985 33884
rect 27019 33881 27031 33915
rect 26973 33875 27031 33881
rect 46477 33915 46535 33921
rect 46477 33881 46489 33915
rect 46523 33912 46535 33915
rect 47486 33912 47492 33924
rect 46523 33884 47492 33912
rect 46523 33881 46535 33884
rect 46477 33875 46535 33881
rect 47486 33872 47492 33884
rect 47544 33872 47550 33924
rect 48133 33915 48191 33921
rect 48133 33881 48145 33915
rect 48179 33881 48191 33915
rect 48133 33875 48191 33881
rect 22646 33844 22652 33856
rect 21652 33816 22652 33844
rect 22646 33804 22652 33816
rect 22704 33804 22710 33856
rect 23842 33844 23848 33856
rect 23803 33816 23848 33844
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 46198 33804 46204 33856
rect 46256 33844 46262 33856
rect 48148 33844 48176 33875
rect 46256 33816 48176 33844
rect 46256 33804 46262 33816
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 19150 33600 19156 33652
rect 19208 33640 19214 33652
rect 22278 33640 22284 33652
rect 19208 33612 22284 33640
rect 19208 33600 19214 33612
rect 19168 33572 19196 33600
rect 18524 33544 19196 33572
rect 18524 33516 18552 33544
rect 19426 33532 19432 33584
rect 19484 33532 19490 33584
rect 20901 33575 20959 33581
rect 20901 33541 20913 33575
rect 20947 33541 20959 33575
rect 20901 33535 20959 33541
rect 21117 33575 21175 33581
rect 21117 33541 21129 33575
rect 21163 33572 21175 33575
rect 21726 33572 21732 33584
rect 21163 33544 21732 33572
rect 21163 33541 21175 33544
rect 21117 33535 21175 33541
rect 18506 33504 18512 33516
rect 18419 33476 18512 33504
rect 18506 33464 18512 33476
rect 18564 33464 18570 33516
rect 20916 33504 20944 33535
rect 21726 33532 21732 33544
rect 21784 33532 21790 33584
rect 21836 33513 21864 33612
rect 22278 33600 22284 33612
rect 22336 33640 22342 33652
rect 24210 33640 24216 33652
rect 22336 33612 24216 33640
rect 22336 33600 22342 33612
rect 24210 33600 24216 33612
rect 24268 33600 24274 33652
rect 24578 33640 24584 33652
rect 24539 33612 24584 33640
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 28626 33640 28632 33652
rect 28587 33612 28632 33640
rect 28626 33600 28632 33612
rect 28684 33600 28690 33652
rect 47854 33600 47860 33652
rect 47912 33640 47918 33652
rect 48041 33643 48099 33649
rect 48041 33640 48053 33643
rect 47912 33612 48053 33640
rect 47912 33600 47918 33612
rect 48041 33609 48053 33612
rect 48087 33609 48099 33643
rect 48041 33603 48099 33609
rect 22097 33575 22155 33581
rect 22097 33541 22109 33575
rect 22143 33572 22155 33575
rect 22370 33572 22376 33584
rect 22143 33544 22376 33572
rect 22143 33541 22155 33544
rect 22097 33535 22155 33541
rect 22370 33532 22376 33544
rect 22428 33532 22434 33584
rect 22738 33532 22744 33584
rect 22796 33532 22802 33584
rect 25869 33575 25927 33581
rect 25869 33541 25881 33575
rect 25915 33572 25927 33575
rect 26142 33572 26148 33584
rect 25915 33544 26148 33572
rect 25915 33541 25927 33544
rect 25869 33535 25927 33541
rect 26142 33532 26148 33544
rect 26200 33532 26206 33584
rect 28350 33572 28356 33584
rect 27540 33544 28356 33572
rect 21821 33507 21879 33513
rect 20916 33476 21404 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1670 33436 1676 33448
rect 1631 33408 1676 33436
rect 1670 33396 1676 33408
rect 1728 33396 1734 33448
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33436 18843 33439
rect 21266 33436 21272 33448
rect 18831 33408 21272 33436
rect 18831 33405 18843 33408
rect 18785 33399 18843 33405
rect 21266 33396 21272 33408
rect 21324 33396 21330 33448
rect 21376 33368 21404 33476
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 24118 33504 24124 33516
rect 24079 33476 24124 33504
rect 21821 33467 21879 33473
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33473 24455 33507
rect 26050 33504 26056 33516
rect 26011 33476 26056 33504
rect 24397 33467 24455 33473
rect 24302 33436 24308 33448
rect 24263 33408 24308 33436
rect 24302 33396 24308 33408
rect 24360 33396 24366 33448
rect 21376 33340 21956 33368
rect 20257 33303 20315 33309
rect 20257 33269 20269 33303
rect 20303 33300 20315 33303
rect 20530 33300 20536 33312
rect 20303 33272 20536 33300
rect 20303 33269 20315 33272
rect 20257 33263 20315 33269
rect 20530 33260 20536 33272
rect 20588 33260 20594 33312
rect 21085 33303 21143 33309
rect 21085 33269 21097 33303
rect 21131 33300 21143 33303
rect 21174 33300 21180 33312
rect 21131 33272 21180 33300
rect 21131 33269 21143 33272
rect 21085 33263 21143 33269
rect 21174 33260 21180 33272
rect 21232 33260 21238 33312
rect 21269 33303 21327 33309
rect 21269 33269 21281 33303
rect 21315 33300 21327 33303
rect 21358 33300 21364 33312
rect 21315 33272 21364 33300
rect 21315 33269 21327 33272
rect 21269 33263 21327 33269
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 21928 33300 21956 33340
rect 23106 33328 23112 33380
rect 23164 33368 23170 33380
rect 24412 33368 24440 33467
rect 26050 33464 26056 33476
rect 26108 33464 26114 33516
rect 27540 33513 27568 33544
rect 28350 33532 28356 33544
rect 28408 33532 28414 33584
rect 27525 33507 27583 33513
rect 27525 33473 27537 33507
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 27614 33464 27620 33516
rect 27672 33504 27678 33516
rect 28261 33507 28319 33513
rect 28261 33504 28273 33507
rect 27672 33476 28273 33504
rect 27672 33464 27678 33476
rect 28261 33473 28273 33476
rect 28307 33473 28319 33507
rect 28261 33467 28319 33473
rect 34514 33464 34520 33516
rect 34572 33504 34578 33516
rect 34701 33507 34759 33513
rect 34701 33504 34713 33507
rect 34572 33476 34713 33504
rect 34572 33464 34578 33476
rect 34701 33473 34713 33476
rect 34747 33473 34759 33507
rect 47854 33504 47860 33516
rect 47815 33476 47860 33504
rect 34701 33467 34759 33473
rect 47854 33464 47860 33476
rect 47912 33464 47918 33516
rect 27706 33396 27712 33448
rect 27764 33436 27770 33448
rect 27801 33439 27859 33445
rect 27801 33436 27813 33439
rect 27764 33408 27813 33436
rect 27764 33396 27770 33408
rect 27801 33405 27813 33408
rect 27847 33436 27859 33439
rect 28353 33439 28411 33445
rect 28353 33436 28365 33439
rect 27847 33408 28365 33436
rect 27847 33405 27859 33408
rect 27801 33399 27859 33405
rect 28353 33405 28365 33408
rect 28399 33405 28411 33439
rect 28353 33399 28411 33405
rect 34606 33396 34612 33448
rect 34664 33436 34670 33448
rect 34977 33439 35035 33445
rect 34977 33436 34989 33439
rect 34664 33408 34989 33436
rect 34664 33396 34670 33408
rect 34977 33405 34989 33408
rect 35023 33405 35035 33439
rect 34977 33399 35035 33405
rect 23164 33340 24440 33368
rect 26237 33371 26295 33377
rect 23164 33328 23170 33340
rect 26237 33337 26249 33371
rect 26283 33368 26295 33371
rect 26326 33368 26332 33380
rect 26283 33340 26332 33368
rect 26283 33337 26295 33340
rect 26237 33331 26295 33337
rect 26326 33328 26332 33340
rect 26384 33328 26390 33380
rect 34790 33368 34796 33380
rect 34703 33340 34796 33368
rect 34790 33328 34796 33340
rect 34848 33368 34854 33380
rect 35342 33368 35348 33380
rect 34848 33340 35348 33368
rect 34848 33328 34854 33340
rect 35342 33328 35348 33340
rect 35400 33328 35406 33380
rect 22462 33300 22468 33312
rect 21928 33272 22468 33300
rect 22462 33260 22468 33272
rect 22520 33300 22526 33312
rect 23290 33300 23296 33312
rect 22520 33272 23296 33300
rect 22520 33260 22526 33272
rect 23290 33260 23296 33272
rect 23348 33260 23354 33312
rect 23566 33300 23572 33312
rect 23527 33272 23572 33300
rect 23566 33260 23572 33272
rect 23624 33260 23630 33312
rect 24397 33303 24455 33309
rect 24397 33269 24409 33303
rect 24443 33300 24455 33303
rect 25038 33300 25044 33312
rect 24443 33272 25044 33300
rect 24443 33269 24455 33272
rect 24397 33263 24455 33269
rect 25038 33260 25044 33272
rect 25096 33260 25102 33312
rect 27709 33303 27767 33309
rect 27709 33269 27721 33303
rect 27755 33300 27767 33303
rect 27982 33300 27988 33312
rect 27755 33272 27988 33300
rect 27755 33269 27767 33272
rect 27709 33263 27767 33269
rect 27982 33260 27988 33272
rect 28040 33260 28046 33312
rect 28350 33300 28356 33312
rect 28311 33272 28356 33300
rect 28350 33260 28356 33272
rect 28408 33300 28414 33312
rect 28810 33300 28816 33312
rect 28408 33272 28816 33300
rect 28408 33260 28414 33272
rect 28810 33260 28816 33272
rect 28868 33260 28874 33312
rect 29822 33260 29828 33312
rect 29880 33300 29886 33312
rect 31754 33300 31760 33312
rect 29880 33272 31760 33300
rect 29880 33260 29886 33272
rect 31754 33260 31760 33272
rect 31812 33300 31818 33312
rect 32766 33300 32772 33312
rect 31812 33272 32772 33300
rect 31812 33260 31818 33272
rect 32766 33260 32772 33272
rect 32824 33260 32830 33312
rect 34885 33303 34943 33309
rect 34885 33269 34897 33303
rect 34931 33300 34943 33303
rect 35526 33300 35532 33312
rect 34931 33272 35532 33300
rect 34931 33269 34943 33272
rect 34885 33263 34943 33269
rect 35526 33260 35532 33272
rect 35584 33260 35590 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 20898 33056 20904 33108
rect 20956 33096 20962 33108
rect 20993 33099 21051 33105
rect 20993 33096 21005 33099
rect 20956 33068 21005 33096
rect 20956 33056 20962 33068
rect 20993 33065 21005 33068
rect 21039 33065 21051 33099
rect 22646 33096 22652 33108
rect 22607 33068 22652 33096
rect 20993 33059 21051 33065
rect 22646 33056 22652 33068
rect 22704 33056 22710 33108
rect 25133 33099 25191 33105
rect 25133 33065 25145 33099
rect 25179 33096 25191 33099
rect 25590 33096 25596 33108
rect 25179 33068 25596 33096
rect 25179 33065 25191 33068
rect 25133 33059 25191 33065
rect 25590 33056 25596 33068
rect 25648 33096 25654 33108
rect 26050 33096 26056 33108
rect 25648 33068 26056 33096
rect 25648 33056 25654 33068
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 26145 33099 26203 33105
rect 26145 33065 26157 33099
rect 26191 33065 26203 33099
rect 28442 33096 28448 33108
rect 28403 33068 28448 33096
rect 26145 33059 26203 33065
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 21358 33028 21364 33040
rect 21284 33000 21364 33028
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 1397 32923 1455 32929
rect 16945 32963 17003 32969
rect 16945 32929 16957 32963
rect 16991 32960 17003 32963
rect 17954 32960 17960 32972
rect 16991 32932 17960 32960
rect 16991 32929 17003 32932
rect 16945 32923 17003 32929
rect 17954 32920 17960 32932
rect 18012 32960 18018 32972
rect 18506 32960 18512 32972
rect 18012 32932 18512 32960
rect 18012 32920 18018 32932
rect 18506 32920 18512 32932
rect 18564 32920 18570 32972
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 19208 32864 19257 32892
rect 19208 32852 19214 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32861 20407 32895
rect 20530 32892 20536 32904
rect 20491 32864 20536 32892
rect 20349 32855 20407 32861
rect 1394 32784 1400 32836
rect 1452 32824 1458 32836
rect 1581 32827 1639 32833
rect 1581 32824 1593 32827
rect 1452 32796 1593 32824
rect 1452 32784 1458 32796
rect 1581 32793 1593 32796
rect 1627 32793 1639 32827
rect 1581 32787 1639 32793
rect 3237 32827 3295 32833
rect 3237 32793 3249 32827
rect 3283 32824 3295 32827
rect 3786 32824 3792 32836
rect 3283 32796 3792 32824
rect 3283 32793 3295 32796
rect 3237 32787 3295 32793
rect 3786 32784 3792 32796
rect 3844 32784 3850 32836
rect 17218 32824 17224 32836
rect 17179 32796 17224 32824
rect 17218 32784 17224 32796
rect 17276 32784 17282 32836
rect 19337 32827 19395 32833
rect 19337 32824 19349 32827
rect 18446 32796 19349 32824
rect 19337 32793 19349 32796
rect 19383 32793 19395 32827
rect 20364 32824 20392 32855
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 21284 32901 21312 33000
rect 21358 32988 21364 33000
rect 21416 32988 21422 33040
rect 21542 32988 21548 33040
rect 21600 33028 21606 33040
rect 21600 33000 21680 33028
rect 21600 32988 21606 33000
rect 21652 32960 21680 33000
rect 22830 32988 22836 33040
rect 22888 33028 22894 33040
rect 23017 33031 23075 33037
rect 23017 33028 23029 33031
rect 22888 33000 23029 33028
rect 22888 32988 22894 33000
rect 23017 32997 23029 33000
rect 23063 33028 23075 33031
rect 25222 33028 25228 33040
rect 23063 33000 25228 33028
rect 23063 32997 23075 33000
rect 23017 32991 23075 32997
rect 25222 32988 25228 33000
rect 25280 33028 25286 33040
rect 25409 33031 25467 33037
rect 25409 33028 25421 33031
rect 25280 33000 25421 33028
rect 25280 32988 25286 33000
rect 25409 32997 25421 33000
rect 25455 32997 25467 33031
rect 25409 32991 25467 32997
rect 25866 32988 25872 33040
rect 25924 33028 25930 33040
rect 26160 33028 26188 33059
rect 28442 33056 28448 33068
rect 28500 33056 28506 33108
rect 30558 33096 30564 33108
rect 28966 33068 30564 33096
rect 25924 33000 26188 33028
rect 25924 32988 25930 33000
rect 27246 32988 27252 33040
rect 27304 33028 27310 33040
rect 27709 33031 27767 33037
rect 27709 33028 27721 33031
rect 27304 33000 27721 33028
rect 27304 32988 27310 33000
rect 27709 32997 27721 33000
rect 27755 32997 27767 33031
rect 28966 33028 28994 33068
rect 30558 33056 30564 33068
rect 30616 33096 30622 33108
rect 31570 33096 31576 33108
rect 30616 33068 31576 33096
rect 30616 33056 30622 33068
rect 31570 33056 31576 33068
rect 31628 33056 31634 33108
rect 33042 33056 33048 33108
rect 33100 33096 33106 33108
rect 35894 33096 35900 33108
rect 33100 33068 35900 33096
rect 33100 33056 33106 33068
rect 35894 33056 35900 33068
rect 35952 33056 35958 33108
rect 27709 32991 27767 32997
rect 28000 33000 28994 33028
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 21652 32932 22937 32960
rect 22925 32929 22937 32932
rect 22971 32960 22983 32963
rect 23658 32960 23664 32972
rect 22971 32932 23664 32960
rect 22971 32929 22983 32932
rect 22925 32923 22983 32929
rect 23658 32920 23664 32932
rect 23716 32960 23722 32972
rect 24394 32960 24400 32972
rect 23716 32932 24400 32960
rect 23716 32920 23722 32932
rect 24394 32920 24400 32932
rect 24452 32920 24458 32972
rect 25130 32960 25136 32972
rect 25043 32932 25136 32960
rect 25130 32920 25136 32932
rect 25188 32960 25194 32972
rect 26142 32960 26148 32972
rect 25188 32932 26148 32960
rect 25188 32920 25194 32932
rect 26142 32920 26148 32932
rect 26200 32920 26206 32972
rect 28000 32960 28028 33000
rect 29822 32988 29828 33040
rect 29880 33028 29886 33040
rect 29880 33000 29925 33028
rect 29880 32988 29886 33000
rect 30006 32988 30012 33040
rect 30064 33028 30070 33040
rect 33410 33028 33416 33040
rect 30064 33000 33416 33028
rect 30064 32988 30070 33000
rect 27632 32932 28028 32960
rect 21269 32895 21327 32901
rect 21269 32861 21281 32895
rect 21315 32861 21327 32895
rect 21269 32855 21327 32861
rect 21358 32892 21416 32898
rect 21358 32858 21370 32892
rect 21404 32858 21416 32892
rect 21358 32852 21416 32858
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32892 21511 32895
rect 21637 32895 21695 32901
rect 21499 32864 21588 32892
rect 21499 32861 21511 32864
rect 21453 32855 21511 32861
rect 20990 32824 20996 32836
rect 20364 32796 20996 32824
rect 19337 32787 19395 32793
rect 20990 32784 20996 32796
rect 21048 32784 21054 32836
rect 18046 32716 18052 32768
rect 18104 32756 18110 32768
rect 18693 32759 18751 32765
rect 18693 32756 18705 32759
rect 18104 32728 18705 32756
rect 18104 32716 18110 32728
rect 18693 32725 18705 32728
rect 18739 32756 18751 32759
rect 20346 32756 20352 32768
rect 18739 32728 20352 32756
rect 18739 32725 18751 32728
rect 18693 32719 18751 32725
rect 20346 32716 20352 32728
rect 20404 32716 20410 32768
rect 20441 32759 20499 32765
rect 20441 32725 20453 32759
rect 20487 32756 20499 32759
rect 20714 32756 20720 32768
rect 20487 32728 20720 32756
rect 20487 32725 20499 32728
rect 20441 32719 20499 32725
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 21008 32756 21036 32784
rect 21376 32756 21404 32852
rect 21560 32836 21588 32864
rect 21637 32861 21649 32895
rect 21683 32861 21695 32895
rect 21637 32855 21695 32861
rect 21542 32784 21548 32836
rect 21600 32784 21606 32836
rect 21008 32728 21404 32756
rect 21652 32756 21680 32855
rect 22646 32852 22652 32904
rect 22704 32892 22710 32904
rect 22833 32895 22891 32901
rect 22833 32892 22845 32895
rect 22704 32864 22845 32892
rect 22704 32852 22710 32864
rect 22833 32861 22845 32864
rect 22879 32861 22891 32895
rect 22833 32855 22891 32861
rect 23014 32852 23020 32904
rect 23072 32892 23078 32904
rect 23109 32895 23167 32901
rect 23109 32892 23121 32895
rect 23072 32864 23121 32892
rect 23072 32852 23078 32864
rect 23109 32861 23121 32864
rect 23155 32861 23167 32895
rect 23109 32855 23167 32861
rect 23293 32895 23351 32901
rect 23293 32861 23305 32895
rect 23339 32892 23351 32895
rect 23566 32892 23572 32904
rect 23339 32864 23572 32892
rect 23339 32861 23351 32864
rect 23293 32855 23351 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 25038 32852 25044 32904
rect 25096 32892 25102 32904
rect 25225 32895 25283 32901
rect 25225 32892 25237 32895
rect 25096 32864 25237 32892
rect 25096 32852 25102 32864
rect 25225 32861 25237 32864
rect 25271 32892 25283 32895
rect 25961 32895 26019 32901
rect 25271 32864 25912 32892
rect 25271 32861 25283 32864
rect 25225 32855 25283 32861
rect 24302 32784 24308 32836
rect 24360 32824 24366 32836
rect 24949 32827 25007 32833
rect 24949 32824 24961 32827
rect 24360 32796 24961 32824
rect 24360 32784 24366 32796
rect 24949 32793 24961 32796
rect 24995 32824 25007 32827
rect 25498 32824 25504 32836
rect 24995 32796 25504 32824
rect 24995 32793 25007 32796
rect 24949 32787 25007 32793
rect 25498 32784 25504 32796
rect 25556 32784 25562 32836
rect 25884 32824 25912 32864
rect 25961 32861 25973 32895
rect 26007 32892 26019 32895
rect 26050 32892 26056 32904
rect 26007 32864 26056 32892
rect 26007 32861 26019 32864
rect 25961 32855 26019 32861
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 27632 32824 27660 32932
rect 28074 32920 28080 32972
rect 28132 32960 28138 32972
rect 28905 32963 28963 32969
rect 28905 32960 28917 32963
rect 28132 32932 28917 32960
rect 28132 32920 28138 32932
rect 28905 32929 28917 32932
rect 28951 32929 28963 32963
rect 28905 32923 28963 32929
rect 30650 32920 30656 32972
rect 30708 32960 30714 32972
rect 30745 32963 30803 32969
rect 30745 32960 30757 32963
rect 30708 32932 30757 32960
rect 30708 32920 30714 32932
rect 30745 32929 30757 32932
rect 30791 32929 30803 32963
rect 30745 32923 30803 32929
rect 27982 32892 27988 32904
rect 27943 32864 27988 32892
rect 27982 32852 27988 32864
rect 28040 32852 28046 32904
rect 28166 32852 28172 32904
rect 28224 32892 28230 32904
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28224 32864 28641 32892
rect 28224 32852 28230 32864
rect 28629 32861 28641 32864
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 28721 32895 28779 32901
rect 28721 32861 28733 32895
rect 28767 32892 28779 32895
rect 28810 32892 28816 32904
rect 28767 32864 28816 32892
rect 28767 32861 28779 32864
rect 28721 32855 28779 32861
rect 28810 32852 28816 32864
rect 28868 32852 28874 32904
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 30006 32892 30012 32904
rect 29052 32864 30012 32892
rect 29052 32852 29058 32864
rect 30006 32852 30012 32864
rect 30064 32852 30070 32904
rect 30466 32892 30472 32904
rect 30427 32864 30472 32892
rect 30466 32852 30472 32864
rect 30524 32852 30530 32904
rect 30558 32852 30564 32904
rect 30616 32892 30622 32904
rect 30852 32901 30880 33000
rect 33410 32988 33416 33000
rect 33468 32988 33474 33040
rect 31754 32960 31760 32972
rect 31715 32932 31760 32960
rect 31754 32920 31760 32932
rect 31812 32920 31818 32972
rect 35253 32963 35311 32969
rect 35253 32929 35265 32963
rect 35299 32960 35311 32963
rect 35710 32960 35716 32972
rect 35299 32932 35716 32960
rect 35299 32929 35311 32932
rect 35253 32923 35311 32929
rect 35710 32920 35716 32932
rect 35768 32920 35774 32972
rect 30837 32895 30895 32901
rect 30616 32864 30661 32892
rect 30616 32852 30622 32864
rect 30837 32861 30849 32895
rect 30883 32861 30895 32895
rect 30837 32855 30895 32861
rect 31481 32895 31539 32901
rect 31481 32861 31493 32895
rect 31527 32861 31539 32895
rect 31662 32892 31668 32904
rect 31623 32864 31668 32892
rect 31481 32855 31539 32861
rect 25884 32796 27660 32824
rect 27709 32827 27767 32833
rect 27709 32793 27721 32827
rect 27755 32824 27767 32827
rect 29546 32824 29552 32836
rect 27755 32796 29552 32824
rect 27755 32793 27767 32796
rect 27709 32787 27767 32793
rect 29546 32784 29552 32796
rect 29604 32824 29610 32836
rect 29641 32827 29699 32833
rect 29641 32824 29653 32827
rect 29604 32796 29653 32824
rect 29604 32784 29610 32796
rect 29641 32793 29653 32796
rect 29687 32793 29699 32827
rect 29641 32787 29699 32793
rect 30285 32827 30343 32833
rect 30285 32793 30297 32827
rect 30331 32824 30343 32827
rect 31496 32824 31524 32855
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 32214 32852 32220 32904
rect 32272 32892 32278 32904
rect 32401 32895 32459 32901
rect 32272 32864 32317 32892
rect 32272 32852 32278 32864
rect 32401 32861 32413 32895
rect 32447 32892 32459 32895
rect 34790 32892 34796 32904
rect 32447 32864 34796 32892
rect 32447 32861 32459 32864
rect 32401 32855 32459 32861
rect 32416 32824 32444 32855
rect 34790 32852 34796 32864
rect 34848 32852 34854 32904
rect 35069 32895 35127 32901
rect 35069 32861 35081 32895
rect 35115 32861 35127 32895
rect 35069 32855 35127 32861
rect 35345 32895 35403 32901
rect 35345 32861 35357 32895
rect 35391 32892 35403 32895
rect 35434 32892 35440 32904
rect 35391 32864 35440 32892
rect 35391 32861 35403 32864
rect 35345 32855 35403 32861
rect 30331 32796 31524 32824
rect 32232 32796 32444 32824
rect 35084 32824 35112 32855
rect 35434 32852 35440 32864
rect 35492 32852 35498 32904
rect 35802 32892 35808 32904
rect 35763 32864 35808 32892
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 35618 32824 35624 32836
rect 35084 32796 35624 32824
rect 30331 32793 30343 32796
rect 30285 32787 30343 32793
rect 23014 32756 23020 32768
rect 21652 32728 23020 32756
rect 23014 32716 23020 32728
rect 23072 32716 23078 32768
rect 25866 32716 25872 32768
rect 25924 32756 25930 32768
rect 26142 32756 26148 32768
rect 25924 32728 26148 32756
rect 25924 32716 25930 32728
rect 26142 32716 26148 32728
rect 26200 32716 26206 32768
rect 27893 32759 27951 32765
rect 27893 32725 27905 32759
rect 27939 32756 27951 32759
rect 28534 32756 28540 32768
rect 27939 32728 28540 32756
rect 27939 32725 27951 32728
rect 27893 32719 27951 32725
rect 28534 32716 28540 32728
rect 28592 32716 28598 32768
rect 30374 32716 30380 32768
rect 30432 32756 30438 32768
rect 31297 32759 31355 32765
rect 31297 32756 31309 32759
rect 30432 32728 31309 32756
rect 30432 32716 30438 32728
rect 31297 32725 31309 32728
rect 31343 32725 31355 32759
rect 31297 32719 31355 32725
rect 31386 32716 31392 32768
rect 31444 32756 31450 32768
rect 32232 32756 32260 32796
rect 35618 32784 35624 32796
rect 35676 32784 35682 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 47670 32824 47676 32836
rect 46523 32796 47676 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 47670 32784 47676 32796
rect 47728 32784 47734 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 31444 32728 32260 32756
rect 32309 32759 32367 32765
rect 31444 32716 31450 32728
rect 32309 32725 32321 32759
rect 32355 32756 32367 32759
rect 32582 32756 32588 32768
rect 32355 32728 32588 32756
rect 32355 32725 32367 32728
rect 32309 32719 32367 32725
rect 32582 32716 32588 32728
rect 32640 32716 32646 32768
rect 34885 32759 34943 32765
rect 34885 32725 34897 32759
rect 34931 32756 34943 32759
rect 35066 32756 35072 32768
rect 34931 32728 35072 32756
rect 34931 32725 34943 32728
rect 34885 32719 34943 32725
rect 35066 32716 35072 32728
rect 35124 32716 35130 32768
rect 35897 32759 35955 32765
rect 35897 32725 35909 32759
rect 35943 32756 35955 32759
rect 36078 32756 36084 32768
rect 35943 32728 36084 32756
rect 35943 32725 35955 32728
rect 35897 32719 35955 32725
rect 36078 32716 36084 32728
rect 36136 32716 36142 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 17218 32512 17224 32564
rect 17276 32552 17282 32564
rect 18509 32555 18567 32561
rect 18509 32552 18521 32555
rect 17276 32524 18521 32552
rect 17276 32512 17282 32524
rect 18509 32521 18521 32524
rect 18555 32521 18567 32555
rect 18509 32515 18567 32521
rect 20530 32512 20536 32564
rect 20588 32552 20594 32564
rect 21542 32552 21548 32564
rect 20588 32524 21548 32552
rect 20588 32512 20594 32524
rect 21542 32512 21548 32524
rect 21600 32512 21606 32564
rect 22278 32552 22284 32564
rect 22239 32524 22284 32552
rect 22278 32512 22284 32524
rect 22336 32512 22342 32564
rect 22370 32512 22376 32564
rect 22428 32552 22434 32564
rect 23201 32555 23259 32561
rect 23201 32552 23213 32555
rect 22428 32524 23213 32552
rect 22428 32512 22434 32524
rect 23201 32521 23213 32524
rect 23247 32552 23259 32555
rect 24118 32552 24124 32564
rect 23247 32524 24124 32552
rect 23247 32521 23259 32524
rect 23201 32515 23259 32521
rect 24118 32512 24124 32524
rect 24176 32512 24182 32564
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 26234 32552 26240 32564
rect 24820 32524 26004 32552
rect 26195 32524 26240 32552
rect 24820 32512 24826 32524
rect 1670 32444 1676 32496
rect 1728 32484 1734 32496
rect 2133 32487 2191 32493
rect 2133 32484 2145 32487
rect 1728 32456 2145 32484
rect 1728 32444 1734 32456
rect 2133 32453 2145 32456
rect 2179 32453 2191 32487
rect 2133 32447 2191 32453
rect 16942 32444 16948 32496
rect 17000 32484 17006 32496
rect 18138 32484 18144 32496
rect 17000 32456 18144 32484
rect 17000 32444 17006 32456
rect 18138 32444 18144 32456
rect 18196 32444 18202 32496
rect 22189 32487 22247 32493
rect 22189 32453 22201 32487
rect 22235 32484 22247 32487
rect 23750 32484 23756 32496
rect 22235 32456 23756 32484
rect 22235 32453 22247 32456
rect 22189 32447 22247 32453
rect 23750 32444 23756 32456
rect 23808 32444 23814 32496
rect 24578 32484 24584 32496
rect 23860 32456 24440 32484
rect 24539 32456 24584 32484
rect 23860 32428 23888 32456
rect 17770 32416 17776 32428
rect 17731 32388 17776 32416
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 17957 32419 18015 32425
rect 17957 32416 17969 32419
rect 17880 32388 17969 32416
rect 1946 32348 1952 32360
rect 1907 32320 1952 32348
rect 1946 32308 1952 32320
rect 2004 32308 2010 32360
rect 3786 32348 3792 32360
rect 3747 32320 3792 32348
rect 3786 32308 3792 32320
rect 3844 32308 3850 32360
rect 17880 32212 17908 32388
rect 17957 32385 17969 32388
rect 18003 32385 18015 32419
rect 17957 32379 18015 32385
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 18380 32388 18425 32416
rect 18380 32376 18386 32388
rect 22646 32376 22652 32428
rect 22704 32416 22710 32428
rect 22833 32419 22891 32425
rect 22833 32416 22845 32419
rect 22704 32388 22845 32416
rect 22704 32376 22710 32388
rect 22833 32385 22845 32388
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32416 23075 32419
rect 23566 32416 23572 32428
rect 23063 32388 23572 32416
rect 23063 32385 23075 32388
rect 23017 32379 23075 32385
rect 18046 32348 18052 32360
rect 18007 32320 18052 32348
rect 18046 32308 18052 32320
rect 18104 32308 18110 32360
rect 18138 32308 18144 32360
rect 18196 32348 18202 32360
rect 22848 32348 22876 32379
rect 23566 32376 23572 32388
rect 23624 32376 23630 32428
rect 23842 32416 23848 32428
rect 23803 32388 23848 32416
rect 23842 32376 23848 32388
rect 23900 32376 23906 32428
rect 24412 32416 24440 32456
rect 24578 32444 24584 32456
rect 24636 32444 24642 32496
rect 25976 32484 26004 32524
rect 26234 32512 26240 32524
rect 26292 32512 26298 32564
rect 28077 32555 28135 32561
rect 28077 32521 28089 32555
rect 28123 32552 28135 32555
rect 28258 32552 28264 32564
rect 28123 32524 28264 32552
rect 28123 32521 28135 32524
rect 28077 32515 28135 32521
rect 28258 32512 28264 32524
rect 28316 32552 28322 32564
rect 31846 32552 31852 32564
rect 28316 32524 28856 32552
rect 28316 32512 28322 32524
rect 28828 32496 28856 32524
rect 29840 32524 31852 32552
rect 27985 32487 28043 32493
rect 25976 32456 27384 32484
rect 24857 32419 24915 32425
rect 24857 32416 24869 32419
rect 24412 32388 24869 32416
rect 24857 32385 24869 32388
rect 24903 32385 24915 32419
rect 24857 32379 24915 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32416 26019 32419
rect 26050 32416 26056 32428
rect 26007 32388 26056 32416
rect 26007 32385 26019 32388
rect 25961 32379 26019 32385
rect 26050 32376 26056 32388
rect 26108 32376 26114 32428
rect 26142 32376 26148 32428
rect 26200 32416 26206 32428
rect 27249 32419 27307 32425
rect 27249 32416 27261 32419
rect 26200 32388 27261 32416
rect 26200 32376 26206 32388
rect 27249 32385 27261 32388
rect 27295 32385 27307 32419
rect 27356 32416 27384 32456
rect 27985 32453 27997 32487
rect 28031 32484 28043 32487
rect 28166 32484 28172 32496
rect 28031 32456 28172 32484
rect 28031 32453 28043 32456
rect 27985 32447 28043 32453
rect 28166 32444 28172 32456
rect 28224 32444 28230 32496
rect 28810 32444 28816 32496
rect 28868 32444 28874 32496
rect 28905 32487 28963 32493
rect 28905 32453 28917 32487
rect 28951 32484 28963 32487
rect 28994 32484 29000 32496
rect 28951 32456 29000 32484
rect 28951 32453 28963 32456
rect 28905 32447 28963 32453
rect 28994 32444 29000 32456
rect 29052 32444 29058 32496
rect 28442 32416 28448 32428
rect 27356 32388 28448 32416
rect 27249 32379 27307 32385
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 28718 32416 28724 32428
rect 28679 32388 28724 32416
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 29840 32360 29868 32524
rect 31846 32512 31852 32524
rect 31904 32552 31910 32564
rect 32674 32552 32680 32564
rect 31904 32524 32680 32552
rect 31904 32512 31910 32524
rect 32674 32512 32680 32524
rect 32732 32512 32738 32564
rect 33781 32555 33839 32561
rect 33781 32552 33793 32555
rect 32784 32524 33793 32552
rect 30101 32487 30159 32493
rect 30101 32453 30113 32487
rect 30147 32484 30159 32487
rect 30374 32484 30380 32496
rect 30147 32456 30380 32484
rect 30147 32453 30159 32456
rect 30101 32447 30159 32453
rect 30374 32444 30380 32456
rect 30432 32444 30438 32496
rect 31202 32376 31208 32428
rect 31260 32376 31266 32428
rect 32398 32416 32404 32428
rect 32359 32388 32404 32416
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 32784 32425 32812 32524
rect 33781 32521 33793 32524
rect 33827 32521 33839 32555
rect 47670 32552 47676 32564
rect 47631 32524 47676 32552
rect 33781 32515 33839 32521
rect 47670 32512 47676 32524
rect 47728 32512 47734 32564
rect 32950 32444 32956 32496
rect 33008 32484 33014 32496
rect 35066 32484 35072 32496
rect 33008 32456 33916 32484
rect 35027 32456 35072 32484
rect 33008 32444 33014 32456
rect 32769 32419 32827 32425
rect 32769 32385 32781 32419
rect 32815 32385 32827 32419
rect 32769 32379 32827 32385
rect 33597 32419 33655 32425
rect 33597 32385 33609 32419
rect 33643 32416 33655 32419
rect 33888 32416 33916 32456
rect 35066 32444 35072 32456
rect 35124 32444 35130 32496
rect 36078 32444 36084 32496
rect 36136 32444 36142 32496
rect 34793 32419 34851 32425
rect 34793 32416 34805 32419
rect 33643 32388 33824 32416
rect 33888 32388 34805 32416
rect 33643 32385 33655 32388
rect 33597 32379 33655 32385
rect 23474 32348 23480 32360
rect 18196 32320 18241 32348
rect 22848 32320 23480 32348
rect 18196 32308 18202 32320
rect 23474 32308 23480 32320
rect 23532 32308 23538 32360
rect 24118 32348 24124 32360
rect 24079 32320 24124 32348
rect 24118 32308 24124 32320
rect 24176 32308 24182 32360
rect 24765 32351 24823 32357
rect 24765 32317 24777 32351
rect 24811 32348 24823 32351
rect 25130 32348 25136 32360
rect 24811 32320 25136 32348
rect 24811 32317 24823 32320
rect 24765 32311 24823 32317
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 25498 32308 25504 32360
rect 25556 32348 25562 32360
rect 28258 32348 28264 32360
rect 25556 32320 28264 32348
rect 25556 32308 25562 32320
rect 28258 32308 28264 32320
rect 28316 32308 28322 32360
rect 29822 32348 29828 32360
rect 29783 32320 29828 32348
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 31386 32348 31392 32360
rect 29932 32320 31392 32348
rect 19334 32280 19340 32292
rect 19306 32240 19340 32280
rect 19392 32240 19398 32292
rect 23290 32240 23296 32292
rect 23348 32280 23354 32292
rect 25041 32283 25099 32289
rect 25041 32280 25053 32283
rect 23348 32252 25053 32280
rect 23348 32240 23354 32252
rect 25041 32249 25053 32252
rect 25087 32249 25099 32283
rect 25041 32243 25099 32249
rect 26326 32240 26332 32292
rect 26384 32280 26390 32292
rect 29932 32280 29960 32320
rect 31386 32308 31392 32320
rect 31444 32308 31450 32360
rect 31570 32348 31576 32360
rect 31531 32320 31576 32348
rect 31570 32308 31576 32320
rect 31628 32308 31634 32360
rect 32214 32348 32220 32360
rect 31726 32320 32220 32348
rect 31726 32280 31754 32320
rect 32214 32308 32220 32320
rect 32272 32348 32278 32360
rect 33410 32348 33416 32360
rect 32272 32320 33088 32348
rect 33371 32320 33416 32348
rect 32272 32308 32278 32320
rect 26384 32252 29960 32280
rect 31128 32252 31754 32280
rect 26384 32240 26390 32252
rect 19306 32212 19334 32240
rect 17880 32184 19334 32212
rect 23382 32172 23388 32224
rect 23440 32212 23446 32224
rect 23661 32215 23719 32221
rect 23661 32212 23673 32215
rect 23440 32184 23673 32212
rect 23440 32172 23446 32184
rect 23661 32181 23673 32184
rect 23707 32181 23719 32215
rect 23661 32175 23719 32181
rect 24029 32215 24087 32221
rect 24029 32181 24041 32215
rect 24075 32212 24087 32215
rect 24578 32212 24584 32224
rect 24075 32184 24584 32212
rect 24075 32181 24087 32184
rect 24029 32175 24087 32181
rect 24578 32172 24584 32184
rect 24636 32172 24642 32224
rect 24765 32215 24823 32221
rect 24765 32181 24777 32215
rect 24811 32212 24823 32215
rect 24854 32212 24860 32224
rect 24811 32184 24860 32212
rect 24811 32181 24823 32184
rect 24765 32175 24823 32181
rect 24854 32172 24860 32184
rect 24912 32172 24918 32224
rect 27341 32215 27399 32221
rect 27341 32181 27353 32215
rect 27387 32212 27399 32215
rect 27982 32212 27988 32224
rect 27387 32184 27988 32212
rect 27387 32181 27399 32184
rect 27341 32175 27399 32181
rect 27982 32172 27988 32184
rect 28040 32172 28046 32224
rect 28258 32172 28264 32224
rect 28316 32212 28322 32224
rect 31128 32212 31156 32252
rect 32030 32240 32036 32292
rect 32088 32280 32094 32292
rect 32953 32283 33011 32289
rect 32953 32280 32965 32283
rect 32088 32252 32965 32280
rect 32088 32240 32094 32252
rect 32953 32249 32965 32252
rect 32999 32249 33011 32283
rect 33060 32280 33088 32320
rect 33410 32308 33416 32320
rect 33468 32308 33474 32360
rect 33796 32348 33824 32388
rect 34793 32385 34805 32388
rect 34839 32385 34851 32419
rect 34793 32379 34851 32385
rect 46842 32376 46848 32428
rect 46900 32416 46906 32428
rect 47029 32419 47087 32425
rect 47029 32416 47041 32419
rect 46900 32388 47041 32416
rect 46900 32376 46906 32388
rect 47029 32385 47041 32388
rect 47075 32385 47087 32419
rect 47578 32416 47584 32428
rect 47539 32388 47584 32416
rect 47029 32379 47087 32385
rect 47578 32376 47584 32388
rect 47636 32376 47642 32428
rect 34698 32348 34704 32360
rect 33796 32320 34704 32348
rect 34698 32308 34704 32320
rect 34756 32308 34762 32360
rect 34790 32280 34796 32292
rect 33060 32252 34796 32280
rect 32953 32243 33011 32249
rect 34790 32240 34796 32252
rect 34848 32240 34854 32292
rect 32490 32212 32496 32224
rect 28316 32184 31156 32212
rect 32451 32184 32496 32212
rect 28316 32172 28322 32184
rect 32490 32172 32496 32184
rect 32548 32172 32554 32224
rect 35802 32172 35808 32224
rect 35860 32212 35866 32224
rect 36541 32215 36599 32221
rect 36541 32212 36553 32215
rect 35860 32184 36553 32212
rect 35860 32172 35866 32184
rect 36541 32181 36553 32184
rect 36587 32181 36599 32215
rect 46842 32212 46848 32224
rect 46803 32184 46848 32212
rect 36541 32175 36599 32181
rect 46842 32172 46848 32184
rect 46900 32172 46906 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1394 32008 1400 32020
rect 1355 31980 1400 32008
rect 1394 31968 1400 31980
rect 1452 31968 1458 32020
rect 21910 31968 21916 32020
rect 21968 32008 21974 32020
rect 22189 32011 22247 32017
rect 22189 32008 22201 32011
rect 21968 31980 22201 32008
rect 21968 31968 21974 31980
rect 22189 31977 22201 31980
rect 22235 31977 22247 32011
rect 23382 32008 23388 32020
rect 23343 31980 23388 32008
rect 22189 31971 22247 31977
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 24118 31968 24124 32020
rect 24176 32008 24182 32020
rect 24762 32008 24768 32020
rect 24176 31980 24768 32008
rect 24176 31968 24182 31980
rect 24762 31968 24768 31980
rect 24820 31968 24826 32020
rect 26513 32011 26571 32017
rect 26513 32008 26525 32011
rect 24872 31980 26525 32008
rect 1762 31900 1768 31952
rect 1820 31940 1826 31952
rect 2038 31940 2044 31952
rect 1820 31912 2044 31940
rect 1820 31900 1826 31912
rect 2038 31900 2044 31912
rect 2096 31900 2102 31952
rect 17770 31900 17776 31952
rect 17828 31940 17834 31952
rect 21450 31940 21456 31952
rect 17828 31912 21456 31940
rect 17828 31900 17834 31912
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 22370 31900 22376 31952
rect 22428 31900 22434 31952
rect 23014 31900 23020 31952
rect 23072 31900 23078 31952
rect 23566 31940 23572 31952
rect 23527 31912 23572 31940
rect 23566 31900 23572 31912
rect 23624 31900 23630 31952
rect 24872 31940 24900 31980
rect 26513 31977 26525 31980
rect 26559 31977 26571 32011
rect 26513 31971 26571 31977
rect 28626 31968 28632 32020
rect 28684 32008 28690 32020
rect 30374 32008 30380 32020
rect 28684 31980 30380 32008
rect 28684 31968 28690 31980
rect 30374 31968 30380 31980
rect 30432 31968 30438 32020
rect 31481 32011 31539 32017
rect 31481 31977 31493 32011
rect 31527 32008 31539 32011
rect 31662 32008 31668 32020
rect 31527 31980 31668 32008
rect 31527 31977 31539 31980
rect 31481 31971 31539 31977
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 32214 31968 32220 32020
rect 32272 32008 32278 32020
rect 32398 32008 32404 32020
rect 32272 31980 32404 32008
rect 32272 31968 32278 31980
rect 32398 31968 32404 31980
rect 32456 32008 32462 32020
rect 33781 32011 33839 32017
rect 33781 32008 33793 32011
rect 32456 31980 33793 32008
rect 32456 31968 32462 31980
rect 33781 31977 33793 31980
rect 33827 31977 33839 32011
rect 33781 31971 33839 31977
rect 34330 31968 34336 32020
rect 34388 32008 34394 32020
rect 34701 32011 34759 32017
rect 34701 32008 34713 32011
rect 34388 31980 34713 32008
rect 34388 31968 34394 31980
rect 34701 31977 34713 31980
rect 34747 31977 34759 32011
rect 34701 31971 34759 31977
rect 34790 31968 34796 32020
rect 34848 32008 34854 32020
rect 35161 32011 35219 32017
rect 35161 32008 35173 32011
rect 34848 31980 35173 32008
rect 34848 31968 34854 31980
rect 35161 31977 35173 31980
rect 35207 31977 35219 32011
rect 35161 31971 35219 31977
rect 35618 31968 35624 32020
rect 35676 32008 35682 32020
rect 35713 32011 35771 32017
rect 35713 32008 35725 32011
rect 35676 31980 35725 32008
rect 35676 31968 35682 31980
rect 35713 31977 35725 31980
rect 35759 31977 35771 32011
rect 35713 31971 35771 31977
rect 46290 31968 46296 32020
rect 46348 32008 46354 32020
rect 47673 32011 47731 32017
rect 47673 32008 47685 32011
rect 46348 31980 47685 32008
rect 46348 31968 46354 31980
rect 47673 31977 47685 31980
rect 47719 31977 47731 32011
rect 47673 31971 47731 31977
rect 24228 31912 24900 31940
rect 9306 31832 9312 31884
rect 9364 31872 9370 31884
rect 22278 31872 22284 31884
rect 9364 31844 22284 31872
rect 9364 31832 9370 31844
rect 22278 31832 22284 31844
rect 22336 31832 22342 31884
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 2038 31764 2044 31816
rect 2096 31804 2102 31816
rect 2317 31807 2375 31813
rect 2317 31804 2329 31807
rect 2096 31776 2329 31804
rect 2096 31764 2102 31776
rect 2317 31773 2329 31776
rect 2363 31773 2375 31807
rect 2958 31804 2964 31816
rect 2919 31776 2964 31804
rect 2317 31767 2375 31773
rect 2958 31764 2964 31776
rect 3016 31764 3022 31816
rect 19978 31764 19984 31816
rect 20036 31804 20042 31816
rect 20254 31804 20260 31816
rect 20036 31776 20260 31804
rect 20036 31764 20042 31776
rect 20254 31764 20260 31776
rect 20312 31804 20318 31816
rect 22388 31813 22416 31900
rect 23032 31872 23060 31900
rect 24228 31872 24256 31912
rect 25222 31900 25228 31952
rect 25280 31900 25286 31952
rect 25593 31943 25651 31949
rect 25593 31909 25605 31943
rect 25639 31940 25651 31943
rect 25866 31940 25872 31952
rect 25639 31912 25872 31940
rect 25639 31909 25651 31912
rect 25593 31903 25651 31909
rect 25866 31900 25872 31912
rect 25924 31900 25930 31952
rect 28902 31900 28908 31952
rect 28960 31940 28966 31952
rect 33410 31940 33416 31952
rect 28960 31912 32628 31940
rect 28960 31900 28966 31912
rect 23032 31844 24256 31872
rect 25133 31875 25191 31881
rect 25133 31841 25145 31875
rect 25179 31872 25191 31875
rect 25240 31872 25268 31900
rect 25179 31844 25268 31872
rect 27249 31875 27307 31881
rect 25179 31841 25191 31844
rect 25133 31835 25191 31841
rect 27249 31841 27261 31875
rect 27295 31872 27307 31875
rect 29822 31872 29828 31884
rect 27295 31844 29828 31872
rect 27295 31841 27307 31844
rect 27249 31835 27307 31841
rect 29822 31832 29828 31844
rect 29880 31832 29886 31884
rect 32600 31881 32628 31912
rect 32692 31912 33416 31940
rect 31205 31875 31263 31881
rect 31205 31841 31217 31875
rect 31251 31872 31263 31875
rect 32493 31875 32551 31881
rect 31251 31844 31892 31872
rect 31251 31841 31263 31844
rect 31205 31835 31263 31841
rect 20533 31807 20591 31813
rect 20533 31804 20545 31807
rect 20312 31776 20545 31804
rect 20312 31764 20318 31776
rect 20533 31773 20545 31776
rect 20579 31773 20591 31807
rect 20533 31767 20591 31773
rect 22189 31807 22247 31813
rect 22189 31773 22201 31807
rect 22235 31773 22247 31807
rect 22189 31767 22247 31773
rect 22373 31807 22431 31813
rect 22373 31773 22385 31807
rect 22419 31773 22431 31807
rect 23014 31804 23020 31816
rect 22975 31776 23020 31804
rect 22373 31767 22431 31773
rect 20901 31739 20959 31745
rect 20901 31705 20913 31739
rect 20947 31736 20959 31739
rect 22094 31736 22100 31748
rect 20947 31708 22100 31736
rect 20947 31705 20959 31708
rect 20901 31699 20959 31705
rect 22094 31696 22100 31708
rect 22152 31696 22158 31748
rect 3050 31668 3056 31680
rect 3011 31640 3056 31668
rect 3050 31628 3056 31640
rect 3108 31628 3114 31680
rect 22204 31668 22232 31767
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 23293 31807 23351 31813
rect 23293 31773 23305 31807
rect 23339 31804 23351 31807
rect 23339 31776 23373 31804
rect 23339 31773 23351 31776
rect 23293 31767 23351 31773
rect 23308 31736 23336 31767
rect 23474 31764 23480 31816
rect 23532 31804 23538 31816
rect 25222 31804 25228 31816
rect 23532 31776 25228 31804
rect 23532 31764 23538 31776
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 26326 31804 26332 31816
rect 26287 31776 26332 31804
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 28810 31764 28816 31816
rect 28868 31804 28874 31816
rect 30282 31804 30288 31816
rect 28868 31776 30288 31804
rect 28868 31764 28874 31776
rect 30282 31764 30288 31776
rect 30340 31764 30346 31816
rect 31113 31807 31171 31813
rect 31113 31773 31125 31807
rect 31159 31804 31171 31807
rect 31570 31804 31576 31816
rect 31159 31776 31576 31804
rect 31159 31773 31171 31776
rect 31113 31767 31171 31773
rect 31570 31764 31576 31776
rect 31628 31764 31634 31816
rect 23658 31736 23664 31748
rect 23308 31708 23664 31736
rect 23658 31696 23664 31708
rect 23716 31696 23722 31748
rect 27525 31739 27583 31745
rect 27525 31705 27537 31739
rect 27571 31736 27583 31739
rect 27798 31736 27804 31748
rect 27571 31708 27804 31736
rect 27571 31705 27583 31708
rect 27525 31699 27583 31705
rect 27798 31696 27804 31708
rect 27856 31696 27862 31748
rect 27982 31696 27988 31748
rect 28040 31696 28046 31748
rect 29641 31739 29699 31745
rect 29641 31705 29653 31739
rect 29687 31736 29699 31739
rect 30374 31736 30380 31748
rect 29687 31708 30380 31736
rect 29687 31705 29699 31708
rect 29641 31699 29699 31705
rect 30374 31696 30380 31708
rect 30432 31696 30438 31748
rect 31864 31736 31892 31844
rect 32493 31841 32505 31875
rect 32539 31841 32551 31875
rect 32493 31835 32551 31841
rect 32585 31875 32643 31881
rect 32585 31841 32597 31875
rect 32631 31841 32643 31875
rect 32585 31835 32643 31841
rect 32030 31764 32036 31816
rect 32088 31804 32094 31816
rect 32217 31807 32275 31813
rect 32217 31804 32229 31807
rect 32088 31776 32229 31804
rect 32088 31764 32094 31776
rect 32217 31773 32229 31776
rect 32263 31773 32275 31807
rect 32398 31804 32404 31816
rect 32359 31776 32404 31804
rect 32217 31767 32275 31773
rect 32398 31764 32404 31776
rect 32456 31764 32462 31816
rect 32508 31804 32536 31835
rect 32692 31804 32720 31912
rect 33410 31900 33416 31912
rect 33468 31940 33474 31952
rect 33594 31940 33600 31952
rect 33468 31912 33600 31940
rect 33468 31900 33474 31912
rect 33594 31900 33600 31912
rect 33652 31900 33658 31952
rect 34606 31900 34612 31952
rect 34664 31940 34670 31952
rect 34664 31912 34836 31940
rect 34664 31900 34670 31912
rect 34698 31872 34704 31884
rect 33336 31844 34704 31872
rect 32508 31776 32720 31804
rect 32769 31807 32827 31813
rect 32769 31773 32781 31807
rect 32815 31804 32827 31807
rect 32858 31804 32864 31816
rect 32815 31776 32864 31804
rect 32815 31773 32827 31776
rect 32769 31767 32827 31773
rect 32858 31764 32864 31776
rect 32916 31764 32922 31816
rect 32582 31736 32588 31748
rect 31864 31708 32588 31736
rect 32582 31696 32588 31708
rect 32640 31696 32646 31748
rect 33336 31736 33364 31844
rect 34698 31832 34704 31844
rect 34756 31832 34762 31884
rect 34808 31881 34836 31912
rect 34793 31875 34851 31881
rect 34793 31841 34805 31875
rect 34839 31872 34851 31875
rect 34882 31872 34888 31884
rect 34839 31844 34888 31872
rect 34839 31841 34851 31844
rect 34793 31835 34851 31841
rect 34882 31832 34888 31844
rect 34940 31872 34946 31884
rect 35802 31872 35808 31884
rect 34940 31844 35808 31872
rect 34940 31832 34946 31844
rect 35802 31832 35808 31844
rect 35860 31872 35866 31884
rect 36173 31875 36231 31881
rect 35860 31844 36032 31872
rect 35860 31832 35866 31844
rect 33594 31804 33600 31816
rect 33555 31776 33600 31804
rect 33594 31764 33600 31776
rect 33652 31804 33658 31816
rect 34330 31804 34336 31816
rect 33652 31776 34336 31804
rect 33652 31764 33658 31776
rect 34330 31764 34336 31776
rect 34388 31764 34394 31816
rect 34422 31764 34428 31816
rect 34480 31804 34486 31816
rect 36004 31813 36032 31844
rect 36173 31841 36185 31875
rect 36219 31872 36231 31875
rect 46842 31872 46848 31884
rect 36219 31844 46848 31872
rect 36219 31841 36231 31844
rect 36173 31835 36231 31841
rect 46842 31832 46848 31844
rect 46900 31832 46906 31884
rect 34977 31807 35035 31813
rect 34977 31804 34989 31807
rect 34480 31776 34989 31804
rect 34480 31764 34486 31776
rect 34977 31773 34989 31776
rect 35023 31773 35035 31807
rect 34977 31767 35035 31773
rect 35897 31807 35955 31813
rect 35897 31773 35909 31807
rect 35943 31773 35955 31807
rect 35897 31767 35955 31773
rect 35989 31807 36047 31813
rect 35989 31773 36001 31807
rect 36035 31773 36047 31807
rect 36262 31804 36268 31816
rect 36223 31776 36268 31804
rect 35989 31767 36047 31773
rect 33413 31739 33471 31745
rect 33413 31736 33425 31739
rect 33336 31708 33425 31736
rect 33413 31705 33425 31708
rect 33459 31705 33471 31739
rect 33413 31699 33471 31705
rect 34514 31696 34520 31748
rect 34572 31736 34578 31748
rect 34701 31739 34759 31745
rect 34701 31736 34713 31739
rect 34572 31708 34713 31736
rect 34572 31696 34578 31708
rect 34701 31705 34713 31708
rect 34747 31736 34759 31739
rect 34790 31736 34796 31748
rect 34747 31708 34796 31736
rect 34747 31705 34759 31708
rect 34701 31699 34759 31705
rect 34790 31696 34796 31708
rect 34848 31696 34854 31748
rect 35912 31680 35940 31767
rect 36262 31764 36268 31776
rect 36320 31764 36326 31816
rect 22830 31668 22836 31680
rect 22204 31640 22836 31668
rect 22830 31628 22836 31640
rect 22888 31628 22894 31680
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 28442 31668 28448 31680
rect 27764 31640 28448 31668
rect 27764 31628 27770 31640
rect 28442 31628 28448 31640
rect 28500 31668 28506 31680
rect 28997 31671 29055 31677
rect 28997 31668 29009 31671
rect 28500 31640 29009 31668
rect 28500 31628 28506 31640
rect 28997 31637 29009 31640
rect 29043 31637 29055 31671
rect 32950 31668 32956 31680
rect 32911 31640 32956 31668
rect 28997 31631 29055 31637
rect 32950 31628 32956 31640
rect 33008 31628 33014 31680
rect 35894 31628 35900 31680
rect 35952 31628 35958 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 17954 31464 17960 31476
rect 17328 31436 17960 31464
rect 2225 31399 2283 31405
rect 2225 31365 2237 31399
rect 2271 31396 2283 31399
rect 3050 31396 3056 31408
rect 2271 31368 3056 31396
rect 2271 31365 2283 31368
rect 2225 31359 2283 31365
rect 3050 31356 3056 31368
rect 3108 31356 3114 31408
rect 2038 31328 2044 31340
rect 1999 31300 2044 31328
rect 2038 31288 2044 31300
rect 2096 31288 2102 31340
rect 17328 31337 17356 31436
rect 17954 31424 17960 31436
rect 18012 31424 18018 31476
rect 20898 31464 20904 31476
rect 20272 31436 20904 31464
rect 18598 31356 18604 31408
rect 18656 31356 18662 31408
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 19150 31288 19156 31340
rect 19208 31328 19214 31340
rect 20272 31337 20300 31436
rect 20898 31424 20904 31436
rect 20956 31464 20962 31476
rect 22554 31464 22560 31476
rect 20956 31436 22560 31464
rect 20956 31424 20962 31436
rect 22554 31424 22560 31436
rect 22612 31424 22618 31476
rect 22649 31467 22707 31473
rect 22649 31433 22661 31467
rect 22695 31464 22707 31467
rect 22738 31464 22744 31476
rect 22695 31436 22744 31464
rect 22695 31433 22707 31436
rect 22649 31427 22707 31433
rect 22738 31424 22744 31436
rect 22796 31424 22802 31476
rect 23658 31424 23664 31476
rect 23716 31464 23722 31476
rect 23934 31464 23940 31476
rect 23716 31436 23940 31464
rect 23716 31424 23722 31436
rect 23934 31424 23940 31436
rect 23992 31424 23998 31476
rect 27798 31424 27804 31476
rect 27856 31464 27862 31476
rect 27893 31467 27951 31473
rect 27893 31464 27905 31467
rect 27856 31436 27905 31464
rect 27856 31424 27862 31436
rect 27893 31433 27905 31436
rect 27939 31433 27951 31467
rect 31202 31464 31208 31476
rect 31163 31436 31208 31464
rect 27893 31427 27951 31433
rect 31202 31424 31208 31436
rect 31260 31424 31266 31476
rect 34330 31464 34336 31476
rect 34291 31436 34336 31464
rect 34330 31424 34336 31436
rect 34388 31424 34394 31476
rect 34698 31424 34704 31476
rect 34756 31464 34762 31476
rect 35161 31467 35219 31473
rect 35161 31464 35173 31467
rect 34756 31436 35173 31464
rect 34756 31424 34762 31436
rect 35161 31433 35173 31436
rect 35207 31464 35219 31467
rect 35710 31464 35716 31476
rect 35207 31436 35572 31464
rect 35671 31436 35716 31464
rect 35207 31433 35219 31436
rect 35161 31427 35219 31433
rect 20990 31356 20996 31408
rect 21048 31396 21054 31408
rect 21821 31399 21879 31405
rect 21048 31368 21312 31396
rect 21048 31356 21054 31368
rect 19521 31331 19579 31337
rect 19521 31328 19533 31331
rect 19208 31300 19533 31328
rect 19208 31288 19214 31300
rect 19521 31297 19533 31300
rect 19567 31297 19579 31331
rect 19521 31291 19579 31297
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20257 31291 20315 31297
rect 20441 31331 20499 31337
rect 20441 31297 20453 31331
rect 20487 31297 20499 31331
rect 20898 31328 20904 31340
rect 20859 31300 20904 31328
rect 20441 31291 20499 31297
rect 2774 31260 2780 31272
rect 2735 31232 2780 31260
rect 2774 31220 2780 31232
rect 2832 31220 2838 31272
rect 17589 31263 17647 31269
rect 17589 31229 17601 31263
rect 17635 31260 17647 31263
rect 19242 31260 19248 31272
rect 17635 31232 19248 31260
rect 17635 31229 17647 31232
rect 17589 31223 17647 31229
rect 19242 31220 19248 31232
rect 19300 31220 19306 31272
rect 20456 31260 20484 31291
rect 20898 31288 20904 31300
rect 20956 31288 20962 31340
rect 21082 31328 21088 31340
rect 21008 31300 21088 31328
rect 21008 31260 21036 31300
rect 21082 31288 21088 31300
rect 21140 31328 21146 31340
rect 21284 31337 21312 31368
rect 21821 31365 21833 31399
rect 21867 31396 21879 31399
rect 22186 31396 22192 31408
rect 21867 31368 22192 31396
rect 21867 31365 21879 31368
rect 21821 31359 21879 31365
rect 22186 31356 22192 31368
rect 22244 31356 22250 31408
rect 22572 31396 22600 31424
rect 23014 31396 23020 31408
rect 22572 31368 23020 31396
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 28166 31356 28172 31408
rect 28224 31396 28230 31408
rect 29270 31396 29276 31408
rect 28224 31368 29276 31396
rect 28224 31356 28230 31368
rect 21269 31331 21327 31337
rect 21140 31300 21233 31328
rect 21140 31288 21146 31300
rect 21269 31297 21281 31331
rect 21315 31328 21327 31331
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21315 31300 22017 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 22112 31260 22140 31291
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22557 31331 22615 31337
rect 22557 31328 22569 31331
rect 22336 31300 22569 31328
rect 22336 31288 22342 31300
rect 22557 31297 22569 31300
rect 22603 31328 22615 31331
rect 23937 31331 23995 31337
rect 23937 31328 23949 31331
rect 22603 31300 23949 31328
rect 22603 31297 22615 31300
rect 22557 31291 22615 31297
rect 23937 31297 23949 31300
rect 23983 31328 23995 31331
rect 23983 31300 24072 31328
rect 23983 31297 23995 31300
rect 23937 31291 23995 31297
rect 20456 31232 21036 31260
rect 21652 31232 22140 31260
rect 20456 31192 20484 31232
rect 19076 31164 20484 31192
rect 19076 31136 19104 31164
rect 19058 31124 19064 31136
rect 19019 31096 19064 31124
rect 19058 31084 19064 31096
rect 19116 31084 19122 31136
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 19613 31127 19671 31133
rect 19613 31124 19625 31127
rect 19484 31096 19625 31124
rect 19484 31084 19490 31096
rect 19613 31093 19625 31096
rect 19659 31093 19671 31127
rect 19613 31087 19671 31093
rect 20349 31127 20407 31133
rect 20349 31093 20361 31127
rect 20395 31124 20407 31127
rect 21652 31124 21680 31232
rect 24044 31192 24072 31300
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 25222 31328 25228 31340
rect 25004 31300 25228 31328
rect 25004 31288 25010 31300
rect 25222 31288 25228 31300
rect 25280 31328 25286 31340
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25280 31300 25421 31328
rect 25280 31288 25286 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 27246 31328 27252 31340
rect 27304 31337 27310 31340
rect 27214 31300 27252 31328
rect 25409 31291 25467 31297
rect 27246 31288 27252 31300
rect 27304 31291 27314 31337
rect 27397 31331 27455 31337
rect 27397 31297 27409 31331
rect 27443 31297 27455 31331
rect 27522 31328 27528 31340
rect 27483 31300 27528 31328
rect 27397 31291 27455 31297
rect 27304 31288 27310 31291
rect 25498 31260 25504 31272
rect 25459 31232 25504 31260
rect 25498 31220 25504 31232
rect 25556 31220 25562 31272
rect 25685 31263 25743 31269
rect 25685 31229 25697 31263
rect 25731 31260 25743 31263
rect 26234 31260 26240 31272
rect 25731 31232 26240 31260
rect 25731 31229 25743 31232
rect 25685 31223 25743 31229
rect 26234 31220 26240 31232
rect 26292 31220 26298 31272
rect 27412 31260 27440 31291
rect 27522 31288 27528 31300
rect 27580 31288 27586 31340
rect 27614 31288 27620 31340
rect 27672 31328 27678 31340
rect 27755 31331 27813 31337
rect 27672 31300 27717 31328
rect 27672 31288 27678 31300
rect 27755 31297 27767 31331
rect 27801 31328 27813 31331
rect 28258 31328 28264 31340
rect 27801 31300 28264 31328
rect 27801 31297 27813 31300
rect 27755 31291 27813 31297
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 28368 31337 28396 31368
rect 29270 31356 29276 31368
rect 29328 31356 29334 31408
rect 32861 31399 32919 31405
rect 32861 31365 32873 31399
rect 32907 31396 32919 31399
rect 32950 31396 32956 31408
rect 32907 31368 32956 31396
rect 32907 31365 32919 31368
rect 32861 31359 32919 31365
rect 32950 31356 32956 31368
rect 33008 31356 33014 31408
rect 33502 31356 33508 31408
rect 33560 31356 33566 31408
rect 35342 31396 35348 31408
rect 34808 31368 35348 31396
rect 28353 31331 28411 31337
rect 28353 31297 28365 31331
rect 28399 31297 28411 31331
rect 29178 31328 29184 31340
rect 29139 31300 29184 31328
rect 28353 31291 28411 31297
rect 29178 31288 29184 31300
rect 29236 31288 29242 31340
rect 31113 31331 31171 31337
rect 31113 31297 31125 31331
rect 31159 31328 31171 31331
rect 31159 31300 31754 31328
rect 31159 31297 31171 31300
rect 31113 31291 31171 31297
rect 28442 31260 28448 31272
rect 27412 31232 28448 31260
rect 28442 31220 28448 31232
rect 28500 31220 28506 31272
rect 31128 31260 31156 31291
rect 28966 31232 31156 31260
rect 31726 31260 31754 31300
rect 31846 31288 31852 31340
rect 31904 31328 31910 31340
rect 34808 31337 34836 31368
rect 35342 31356 35348 31368
rect 35400 31356 35406 31408
rect 35544 31396 35572 31436
rect 35710 31424 35716 31436
rect 35768 31424 35774 31476
rect 35544 31368 35848 31396
rect 32585 31331 32643 31337
rect 32585 31328 32597 31331
rect 31904 31300 32597 31328
rect 31904 31288 31910 31300
rect 32585 31297 32597 31300
rect 32631 31297 32643 31331
rect 32585 31291 32643 31297
rect 34793 31331 34851 31337
rect 34793 31297 34805 31331
rect 34839 31297 34851 31331
rect 34793 31291 34851 31297
rect 34882 31288 34888 31340
rect 34940 31328 34946 31340
rect 34940 31300 34985 31328
rect 34940 31288 34946 31300
rect 35526 31288 35532 31340
rect 35584 31328 35590 31340
rect 35820 31337 35848 31368
rect 35621 31331 35679 31337
rect 35621 31328 35633 31331
rect 35584 31300 35633 31328
rect 35584 31288 35590 31300
rect 35621 31297 35633 31300
rect 35667 31297 35679 31331
rect 35621 31291 35679 31297
rect 35805 31331 35863 31337
rect 35805 31297 35817 31331
rect 35851 31297 35863 31331
rect 35805 31291 35863 31297
rect 33410 31260 33416 31272
rect 31726 31232 33416 31260
rect 28966 31192 28994 31232
rect 33410 31220 33416 31232
rect 33468 31220 33474 31272
rect 24044 31164 28994 31192
rect 29365 31195 29423 31201
rect 29365 31161 29377 31195
rect 29411 31192 29423 31195
rect 30374 31192 30380 31204
rect 29411 31164 30380 31192
rect 29411 31161 29423 31164
rect 29365 31155 29423 31161
rect 30374 31152 30380 31164
rect 30432 31192 30438 31204
rect 30742 31192 30748 31204
rect 30432 31164 30748 31192
rect 30432 31152 30438 31164
rect 30742 31152 30748 31164
rect 30800 31152 30806 31204
rect 21818 31124 21824 31136
rect 20395 31096 21680 31124
rect 21779 31096 21824 31124
rect 20395 31093 20407 31096
rect 20349 31087 20407 31093
rect 21818 31084 21824 31096
rect 21876 31084 21882 31136
rect 24026 31124 24032 31136
rect 23987 31096 24032 31124
rect 24026 31084 24032 31096
rect 24084 31084 24090 31136
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 25041 31127 25099 31133
rect 25041 31124 25053 31127
rect 24636 31096 25053 31124
rect 24636 31084 24642 31096
rect 25041 31093 25053 31096
rect 25087 31093 25099 31127
rect 25041 31087 25099 31093
rect 26786 31084 26792 31136
rect 26844 31124 26850 31136
rect 28537 31127 28595 31133
rect 28537 31124 28549 31127
rect 26844 31096 28549 31124
rect 26844 31084 26850 31096
rect 28537 31093 28549 31096
rect 28583 31093 28595 31127
rect 34790 31124 34796 31136
rect 34751 31096 34796 31124
rect 28537 31087 28595 31093
rect 34790 31084 34796 31096
rect 34848 31084 34854 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 18509 30923 18567 30929
rect 18509 30889 18521 30923
rect 18555 30920 18567 30923
rect 18598 30920 18604 30932
rect 18555 30892 18604 30920
rect 18555 30889 18567 30892
rect 18509 30883 18567 30889
rect 18598 30880 18604 30892
rect 18656 30880 18662 30932
rect 19242 30920 19248 30932
rect 19203 30892 19248 30920
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 20530 30880 20536 30932
rect 20588 30920 20594 30932
rect 21269 30923 21327 30929
rect 21269 30920 21281 30923
rect 20588 30892 21281 30920
rect 20588 30880 20594 30892
rect 21269 30889 21281 30892
rect 21315 30889 21327 30923
rect 21269 30883 21327 30889
rect 27890 30880 27896 30932
rect 27948 30920 27954 30932
rect 28353 30923 28411 30929
rect 28353 30920 28365 30923
rect 27948 30892 28365 30920
rect 27948 30880 27954 30892
rect 28353 30889 28365 30892
rect 28399 30920 28411 30923
rect 28442 30920 28448 30932
rect 28399 30892 28448 30920
rect 28399 30889 28411 30892
rect 28353 30883 28411 30889
rect 28442 30880 28448 30892
rect 28500 30880 28506 30932
rect 33502 30920 33508 30932
rect 33463 30892 33508 30920
rect 33502 30880 33508 30892
rect 33560 30880 33566 30932
rect 19334 30812 19340 30864
rect 19392 30852 19398 30864
rect 19613 30855 19671 30861
rect 19613 30852 19625 30855
rect 19392 30824 19625 30852
rect 19392 30812 19398 30824
rect 19613 30821 19625 30824
rect 19659 30852 19671 30855
rect 20622 30852 20628 30864
rect 19659 30824 20628 30852
rect 19659 30821 19671 30824
rect 19613 30815 19671 30821
rect 20622 30812 20628 30824
rect 20680 30812 20686 30864
rect 20898 30852 20904 30864
rect 20732 30824 20904 30852
rect 19058 30744 19064 30796
rect 19116 30784 19122 30796
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19116 30756 19717 30784
rect 19116 30744 19122 30756
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 18417 30719 18475 30725
rect 18417 30685 18429 30719
rect 18463 30716 18475 30719
rect 19150 30716 19156 30728
rect 18463 30688 19156 30716
rect 18463 30685 18475 30688
rect 18417 30679 18475 30685
rect 19150 30676 19156 30688
rect 19208 30676 19214 30728
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19444 30648 19472 30679
rect 20346 30676 20352 30728
rect 20404 30716 20410 30728
rect 20732 30725 20760 30824
rect 20898 30812 20904 30824
rect 20956 30852 20962 30864
rect 24302 30852 24308 30864
rect 20956 30824 24308 30852
rect 20956 30812 20962 30824
rect 24302 30812 24308 30824
rect 24360 30812 24366 30864
rect 21818 30784 21824 30796
rect 20824 30756 21824 30784
rect 20824 30725 20852 30756
rect 21818 30744 21824 30756
rect 21876 30744 21882 30796
rect 22278 30784 22284 30796
rect 22191 30756 22284 30784
rect 22278 30744 22284 30756
rect 22336 30784 22342 30796
rect 23382 30784 23388 30796
rect 22336 30756 23388 30784
rect 22336 30744 22342 30756
rect 23382 30744 23388 30756
rect 23440 30744 23446 30796
rect 23584 30756 26188 30784
rect 20441 30719 20499 30725
rect 20441 30716 20453 30719
rect 20404 30688 20453 30716
rect 20404 30676 20410 30688
rect 20441 30685 20453 30688
rect 20487 30685 20499 30719
rect 20441 30679 20499 30685
rect 20533 30719 20591 30725
rect 20533 30685 20545 30719
rect 20579 30685 20591 30719
rect 20533 30679 20591 30685
rect 20717 30719 20775 30725
rect 20717 30685 20729 30719
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30685 20867 30719
rect 20809 30679 20867 30685
rect 20257 30651 20315 30657
rect 20257 30648 20269 30651
rect 19444 30620 20269 30648
rect 20257 30617 20269 30620
rect 20303 30617 20315 30651
rect 20548 30648 20576 30679
rect 21082 30676 21088 30728
rect 21140 30716 21146 30728
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 21140 30688 21281 30716
rect 21140 30676 21146 30688
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 21358 30676 21364 30728
rect 21416 30716 21422 30728
rect 22554 30716 22560 30728
rect 21416 30688 21461 30716
rect 22515 30688 22560 30716
rect 21416 30676 21422 30688
rect 22554 30676 22560 30688
rect 22612 30676 22618 30728
rect 20257 30611 20315 30617
rect 20456 30620 20576 30648
rect 20456 30592 20484 30620
rect 20622 30608 20628 30660
rect 20680 30648 20686 30660
rect 23584 30648 23612 30756
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 26160 30716 26188 30756
rect 26234 30744 26240 30796
rect 26292 30784 26298 30796
rect 26292 30756 30052 30784
rect 26292 30744 26298 30756
rect 26786 30716 26792 30728
rect 26160 30688 26792 30716
rect 26786 30676 26792 30688
rect 26844 30676 26850 30728
rect 28169 30719 28227 30725
rect 28169 30685 28181 30719
rect 28215 30716 28227 30719
rect 28718 30716 28724 30728
rect 28215 30688 28724 30716
rect 28215 30685 28227 30688
rect 28169 30679 28227 30685
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 30024 30725 30052 30756
rect 32490 30744 32496 30796
rect 32548 30784 32554 30796
rect 32548 30756 32720 30784
rect 32548 30744 32554 30756
rect 30009 30719 30067 30725
rect 30009 30685 30021 30719
rect 30055 30685 30067 30719
rect 30009 30679 30067 30685
rect 20680 30620 23612 30648
rect 23661 30651 23719 30657
rect 20680 30608 20686 30620
rect 23661 30617 23673 30651
rect 23707 30648 23719 30651
rect 23707 30620 25912 30648
rect 23707 30617 23719 30620
rect 23661 30611 23719 30617
rect 20438 30540 20444 30592
rect 20496 30540 20502 30592
rect 21634 30580 21640 30592
rect 21595 30552 21640 30580
rect 21634 30540 21640 30552
rect 21692 30540 21698 30592
rect 23750 30580 23756 30592
rect 23711 30552 23756 30580
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 23842 30540 23848 30592
rect 23900 30580 23906 30592
rect 24397 30583 24455 30589
rect 24397 30580 24409 30583
rect 23900 30552 24409 30580
rect 23900 30540 23906 30552
rect 24397 30549 24409 30552
rect 24443 30549 24455 30583
rect 25884 30580 25912 30620
rect 25958 30608 25964 30660
rect 26016 30648 26022 30660
rect 29178 30648 29184 30660
rect 26016 30620 26061 30648
rect 27264 30620 29184 30648
rect 26016 30608 26022 30620
rect 27264 30589 27292 30620
rect 29178 30608 29184 30620
rect 29236 30608 29242 30660
rect 30024 30648 30052 30679
rect 30466 30676 30472 30728
rect 30524 30716 30530 30728
rect 32306 30716 32312 30728
rect 30524 30688 30972 30716
rect 32267 30688 32312 30716
rect 30524 30676 30530 30688
rect 30944 30657 30972 30688
rect 32306 30676 32312 30688
rect 32364 30676 32370 30728
rect 32401 30719 32459 30725
rect 32401 30685 32413 30719
rect 32447 30685 32459 30719
rect 32582 30716 32588 30728
rect 32543 30688 32588 30716
rect 32401 30679 32459 30685
rect 30745 30651 30803 30657
rect 30745 30648 30757 30651
rect 30024 30620 30757 30648
rect 30745 30617 30757 30620
rect 30791 30617 30803 30651
rect 30745 30611 30803 30617
rect 30929 30651 30987 30657
rect 30929 30617 30941 30651
rect 30975 30648 30987 30651
rect 31386 30648 31392 30660
rect 30975 30620 31392 30648
rect 30975 30617 30987 30620
rect 30929 30611 30987 30617
rect 31386 30608 31392 30620
rect 31444 30608 31450 30660
rect 32416 30648 32444 30679
rect 32582 30676 32588 30688
rect 32640 30676 32646 30728
rect 32692 30725 32720 30756
rect 32677 30719 32735 30725
rect 32677 30685 32689 30719
rect 32723 30685 32735 30719
rect 33410 30716 33416 30728
rect 33371 30688 33416 30716
rect 32677 30679 32735 30685
rect 33410 30676 33416 30688
rect 33468 30676 33474 30728
rect 32490 30648 32496 30660
rect 32416 30620 32496 30648
rect 32490 30608 32496 30620
rect 32548 30608 32554 30660
rect 27249 30583 27307 30589
rect 27249 30580 27261 30583
rect 25884 30552 27261 30580
rect 24397 30543 24455 30549
rect 27249 30549 27261 30552
rect 27295 30549 27307 30583
rect 27249 30543 27307 30549
rect 29270 30540 29276 30592
rect 29328 30580 29334 30592
rect 30101 30583 30159 30589
rect 30101 30580 30113 30583
rect 29328 30552 30113 30580
rect 29328 30540 29334 30552
rect 30101 30549 30113 30552
rect 30147 30549 30159 30583
rect 30101 30543 30159 30549
rect 32125 30583 32183 30589
rect 32125 30549 32137 30583
rect 32171 30580 32183 30583
rect 32398 30580 32404 30592
rect 32171 30552 32404 30580
rect 32171 30549 32183 30552
rect 32125 30543 32183 30549
rect 32398 30540 32404 30552
rect 32456 30540 32462 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 19613 30379 19671 30385
rect 19613 30345 19625 30379
rect 19659 30345 19671 30379
rect 19613 30339 19671 30345
rect 19426 30308 19432 30320
rect 19366 30280 19432 30308
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 19628 30308 19656 30339
rect 20806 30336 20812 30388
rect 20864 30376 20870 30388
rect 46842 30376 46848 30388
rect 20864 30348 46848 30376
rect 20864 30336 20870 30348
rect 46842 30336 46848 30348
rect 46900 30336 46906 30388
rect 21358 30308 21364 30320
rect 19628 30280 21364 30308
rect 20530 30240 20536 30252
rect 20491 30212 20536 30240
rect 20530 30200 20536 30212
rect 20588 30200 20594 30252
rect 20622 30200 20628 30252
rect 20680 30240 20686 30252
rect 20824 30249 20852 30280
rect 21358 30268 21364 30280
rect 21416 30308 21422 30320
rect 21416 30280 21864 30308
rect 21416 30268 21422 30280
rect 20717 30243 20775 30249
rect 20717 30240 20729 30243
rect 20680 30212 20729 30240
rect 20680 30200 20686 30212
rect 20717 30209 20729 30212
rect 20763 30209 20775 30243
rect 20717 30203 20775 30209
rect 20809 30243 20867 30249
rect 20809 30209 20821 30243
rect 20855 30209 20867 30243
rect 21082 30240 21088 30252
rect 21043 30212 21088 30240
rect 20809 30203 20867 30209
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 21836 30249 21864 30280
rect 24026 30268 24032 30320
rect 24084 30268 24090 30320
rect 25866 30308 25872 30320
rect 25827 30280 25872 30308
rect 25866 30268 25872 30280
rect 25924 30268 25930 30320
rect 28534 30268 28540 30320
rect 28592 30308 28598 30320
rect 28592 30280 28994 30308
rect 28592 30268 28598 30280
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22186 30200 22192 30252
rect 22244 30240 22250 30252
rect 22557 30243 22615 30249
rect 22557 30240 22569 30243
rect 22244 30212 22569 30240
rect 22244 30200 22250 30212
rect 22557 30209 22569 30212
rect 22603 30240 22615 30243
rect 23014 30240 23020 30252
rect 22603 30212 23020 30240
rect 22603 30209 22615 30212
rect 22557 30203 22615 30209
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 25038 30200 25044 30252
rect 25096 30240 25102 30252
rect 25777 30243 25835 30249
rect 25777 30240 25789 30243
rect 25096 30212 25789 30240
rect 25096 30200 25102 30212
rect 25777 30209 25789 30212
rect 25823 30209 25835 30243
rect 25777 30203 25835 30209
rect 26326 30200 26332 30252
rect 26384 30240 26390 30252
rect 26973 30243 27031 30249
rect 26973 30240 26985 30243
rect 26384 30212 26985 30240
rect 26384 30200 26390 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27249 30243 27307 30249
rect 27249 30209 27261 30243
rect 27295 30240 27307 30243
rect 28350 30240 28356 30252
rect 27295 30212 28356 30240
rect 27295 30209 27307 30212
rect 27249 30203 27307 30209
rect 17862 30172 17868 30184
rect 17823 30144 17868 30172
rect 17862 30132 17868 30144
rect 17920 30132 17926 30184
rect 18141 30175 18199 30181
rect 18141 30141 18153 30175
rect 18187 30172 18199 30175
rect 20901 30175 20959 30181
rect 18187 30144 19748 30172
rect 18187 30141 18199 30144
rect 18141 30135 18199 30141
rect 19720 30104 19748 30144
rect 20901 30141 20913 30175
rect 20947 30172 20959 30175
rect 20990 30172 20996 30184
rect 20947 30144 20996 30172
rect 20947 30141 20959 30144
rect 20901 30135 20959 30141
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 23198 30172 23204 30184
rect 23159 30144 23204 30172
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 23477 30175 23535 30181
rect 23477 30141 23489 30175
rect 23523 30172 23535 30175
rect 23842 30172 23848 30184
rect 23523 30144 23848 30172
rect 23523 30141 23535 30144
rect 23477 30135 23535 30141
rect 23842 30132 23848 30144
rect 23900 30132 23906 30184
rect 24946 30172 24952 30184
rect 24907 30144 24952 30172
rect 24946 30132 24952 30144
rect 25004 30132 25010 30184
rect 26053 30175 26111 30181
rect 26053 30141 26065 30175
rect 26099 30172 26111 30175
rect 27264 30172 27292 30203
rect 28350 30200 28356 30212
rect 28408 30240 28414 30252
rect 28629 30243 28687 30249
rect 28629 30240 28641 30243
rect 28408 30212 28641 30240
rect 28408 30200 28414 30212
rect 28629 30209 28641 30212
rect 28675 30240 28687 30243
rect 28718 30240 28724 30252
rect 28675 30212 28724 30240
rect 28675 30209 28687 30212
rect 28629 30203 28687 30209
rect 28718 30200 28724 30212
rect 28776 30200 28782 30252
rect 28966 30240 28994 30280
rect 29546 30268 29552 30320
rect 29604 30308 29610 30320
rect 30282 30308 30288 30320
rect 29604 30280 30288 30308
rect 29604 30268 29610 30280
rect 30282 30268 30288 30280
rect 30340 30308 30346 30320
rect 30377 30311 30435 30317
rect 30377 30308 30389 30311
rect 30340 30280 30389 30308
rect 30340 30268 30346 30280
rect 30377 30277 30389 30280
rect 30423 30277 30435 30311
rect 30377 30271 30435 30277
rect 29365 30243 29423 30249
rect 29365 30240 29377 30243
rect 28966 30212 29377 30240
rect 29365 30209 29377 30212
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 26099 30144 27292 30172
rect 29380 30172 29408 30203
rect 29914 30200 29920 30252
rect 29972 30240 29978 30252
rect 30193 30243 30251 30249
rect 30193 30240 30205 30243
rect 29972 30212 30205 30240
rect 29972 30200 29978 30212
rect 30193 30209 30205 30212
rect 30239 30209 30251 30243
rect 30193 30203 30251 30209
rect 33410 30200 33416 30252
rect 33468 30240 33474 30252
rect 33505 30243 33563 30249
rect 33505 30240 33517 30243
rect 33468 30212 33517 30240
rect 33468 30200 33474 30212
rect 33505 30209 33517 30212
rect 33551 30209 33563 30243
rect 33505 30203 33563 30209
rect 30098 30172 30104 30184
rect 29380 30144 30104 30172
rect 26099 30141 26111 30144
rect 26053 30135 26111 30141
rect 30098 30132 30104 30144
rect 30156 30132 30162 30184
rect 21269 30107 21327 30113
rect 21269 30104 21281 30107
rect 19720 30076 21281 30104
rect 21269 30073 21281 30076
rect 21315 30073 21327 30107
rect 21269 30067 21327 30073
rect 25409 30107 25467 30113
rect 25409 30073 25421 30107
rect 25455 30104 25467 30107
rect 25498 30104 25504 30116
rect 25455 30076 25504 30104
rect 25455 30073 25467 30076
rect 25409 30067 25467 30073
rect 25498 30064 25504 30076
rect 25556 30064 25562 30116
rect 32766 30104 32772 30116
rect 31726 30076 32772 30104
rect 20622 29996 20628 30048
rect 20680 30036 20686 30048
rect 21913 30039 21971 30045
rect 21913 30036 21925 30039
rect 20680 30008 21925 30036
rect 20680 29996 20686 30008
rect 21913 30005 21925 30008
rect 21959 30005 21971 30039
rect 22646 30036 22652 30048
rect 22607 30008 22652 30036
rect 21913 29999 21971 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22830 29996 22836 30048
rect 22888 30036 22894 30048
rect 28534 30036 28540 30048
rect 22888 30008 28540 30036
rect 22888 29996 22894 30008
rect 28534 29996 28540 30008
rect 28592 30036 28598 30048
rect 28813 30039 28871 30045
rect 28813 30036 28825 30039
rect 28592 30008 28825 30036
rect 28592 29996 28598 30008
rect 28813 30005 28825 30008
rect 28859 30005 28871 30039
rect 28813 29999 28871 30005
rect 28902 29996 28908 30048
rect 28960 30036 28966 30048
rect 29549 30039 29607 30045
rect 29549 30036 29561 30039
rect 28960 30008 29561 30036
rect 28960 29996 28966 30008
rect 29549 30005 29561 30008
rect 29595 30036 29607 30039
rect 31726 30036 31754 30076
rect 32766 30064 32772 30076
rect 32824 30064 32830 30116
rect 29595 30008 31754 30036
rect 33597 30039 33655 30045
rect 29595 30005 29607 30008
rect 29549 29999 29607 30005
rect 33597 30005 33609 30039
rect 33643 30036 33655 30039
rect 33686 30036 33692 30048
rect 33643 30008 33692 30036
rect 33643 30005 33655 30008
rect 33597 29999 33655 30005
rect 33686 29996 33692 30008
rect 33744 29996 33750 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 20714 29832 20720 29844
rect 20675 29804 20720 29832
rect 20714 29792 20720 29804
rect 20772 29792 20778 29844
rect 26234 29792 26240 29844
rect 26292 29832 26298 29844
rect 26329 29835 26387 29841
rect 26329 29832 26341 29835
rect 26292 29804 26341 29832
rect 26292 29792 26298 29804
rect 26329 29801 26341 29804
rect 26375 29801 26387 29835
rect 28350 29832 28356 29844
rect 28311 29804 28356 29832
rect 26329 29795 26387 29801
rect 28350 29792 28356 29804
rect 28408 29792 28414 29844
rect 28460 29804 28994 29832
rect 20530 29724 20536 29776
rect 20588 29764 20594 29776
rect 20809 29767 20867 29773
rect 20809 29764 20821 29767
rect 20588 29736 20821 29764
rect 20588 29724 20594 29736
rect 20809 29733 20821 29736
rect 20855 29733 20867 29767
rect 20809 29727 20867 29733
rect 23842 29724 23848 29776
rect 23900 29764 23906 29776
rect 25130 29764 25136 29776
rect 23900 29736 25136 29764
rect 23900 29724 23906 29736
rect 25130 29724 25136 29736
rect 25188 29764 25194 29776
rect 28460 29764 28488 29804
rect 25188 29736 28488 29764
rect 28537 29767 28595 29773
rect 25188 29724 25194 29736
rect 28537 29733 28549 29767
rect 28583 29764 28595 29767
rect 28966 29764 28994 29804
rect 32490 29792 32496 29844
rect 32548 29832 32554 29844
rect 34149 29835 34207 29841
rect 34149 29832 34161 29835
rect 32548 29804 34161 29832
rect 32548 29792 32554 29804
rect 34149 29801 34161 29804
rect 34195 29832 34207 29835
rect 34422 29832 34428 29844
rect 34195 29804 34428 29832
rect 34195 29801 34207 29804
rect 34149 29795 34207 29801
rect 34422 29792 34428 29804
rect 34480 29792 34486 29844
rect 28583 29736 28764 29764
rect 28966 29736 29868 29764
rect 28583 29733 28595 29736
rect 28537 29727 28595 29733
rect 18322 29656 18328 29708
rect 18380 29696 18386 29708
rect 19978 29696 19984 29708
rect 18380 29668 19984 29696
rect 18380 29656 18386 29668
rect 19978 29656 19984 29668
rect 20036 29656 20042 29708
rect 20901 29699 20959 29705
rect 20901 29665 20913 29699
rect 20947 29696 20959 29699
rect 23566 29696 23572 29708
rect 20947 29668 23572 29696
rect 20947 29665 20959 29668
rect 20901 29659 20959 29665
rect 23566 29656 23572 29668
rect 23624 29696 23630 29708
rect 24489 29699 24547 29705
rect 24489 29696 24501 29699
rect 23624 29668 24501 29696
rect 23624 29656 23630 29668
rect 24489 29665 24501 29668
rect 24535 29696 24547 29699
rect 24762 29696 24768 29708
rect 24535 29668 24768 29696
rect 24535 29665 24547 29668
rect 24489 29659 24547 29665
rect 24762 29656 24768 29668
rect 24820 29656 24826 29708
rect 20622 29628 20628 29640
rect 20583 29600 20628 29628
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29628 21051 29631
rect 21082 29628 21088 29640
rect 21039 29600 21088 29628
rect 21039 29597 21051 29600
rect 20993 29591 21051 29597
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 24394 29628 24400 29640
rect 24307 29600 24400 29628
rect 24394 29588 24400 29600
rect 24452 29588 24458 29640
rect 24578 29628 24584 29640
rect 24539 29600 24584 29628
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29628 25191 29631
rect 25406 29628 25412 29640
rect 25179 29600 25412 29628
rect 25179 29597 25191 29600
rect 25133 29591 25191 29597
rect 25406 29588 25412 29600
rect 25464 29628 25470 29640
rect 26237 29631 26295 29637
rect 26237 29628 26249 29631
rect 25464 29600 26249 29628
rect 25464 29588 25470 29600
rect 26237 29597 26249 29600
rect 26283 29597 26295 29631
rect 26237 29591 26295 29597
rect 26326 29588 26332 29640
rect 26384 29628 26390 29640
rect 26421 29631 26479 29637
rect 26421 29628 26433 29631
rect 26384 29600 26433 29628
rect 26384 29588 26390 29600
rect 26421 29597 26433 29600
rect 26467 29597 26479 29631
rect 26421 29591 26479 29597
rect 27614 29588 27620 29640
rect 27672 29628 27678 29640
rect 28736 29628 28764 29736
rect 29549 29631 29607 29637
rect 29549 29628 29561 29631
rect 27672 29600 28304 29628
rect 28736 29600 29561 29628
rect 27672 29588 27678 29600
rect 24412 29560 24440 29588
rect 28166 29560 28172 29572
rect 24412 29532 25268 29560
rect 28127 29532 28172 29560
rect 15378 29452 15384 29504
rect 15436 29492 15442 29504
rect 20530 29492 20536 29504
rect 15436 29464 20536 29492
rect 15436 29452 15442 29464
rect 20530 29452 20536 29464
rect 20588 29452 20594 29504
rect 25240 29501 25268 29532
rect 28166 29520 28172 29532
rect 28224 29520 28230 29572
rect 28276 29560 28304 29600
rect 29549 29597 29561 29600
rect 29595 29597 29607 29631
rect 29549 29591 29607 29597
rect 29639 29588 29645 29640
rect 29697 29628 29703 29640
rect 29697 29600 29742 29628
rect 29697 29588 29703 29600
rect 29840 29569 29868 29736
rect 30006 29724 30012 29776
rect 30064 29764 30070 29776
rect 30064 29736 30972 29764
rect 30064 29724 30070 29736
rect 30055 29631 30113 29637
rect 30055 29597 30067 29631
rect 30101 29628 30113 29631
rect 30742 29628 30748 29640
rect 30101 29600 30604 29628
rect 30703 29600 30748 29628
rect 30101 29597 30113 29600
rect 30055 29591 30113 29597
rect 29825 29563 29883 29569
rect 28276 29532 29776 29560
rect 25225 29495 25283 29501
rect 25225 29461 25237 29495
rect 25271 29492 25283 29495
rect 28369 29495 28427 29501
rect 28369 29492 28381 29495
rect 25271 29464 28381 29492
rect 25271 29461 25283 29464
rect 25225 29455 25283 29461
rect 28369 29461 28381 29464
rect 28415 29461 28427 29495
rect 29748 29492 29776 29532
rect 29825 29529 29837 29563
rect 29871 29529 29883 29563
rect 29825 29523 29883 29529
rect 29917 29563 29975 29569
rect 29917 29529 29929 29563
rect 29963 29529 29975 29563
rect 30576 29560 30604 29600
rect 30742 29588 30748 29600
rect 30800 29588 30806 29640
rect 30944 29637 30972 29736
rect 45370 29656 45376 29708
rect 45428 29696 45434 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 45428 29668 47593 29696
rect 45428 29656 45434 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 30929 29631 30987 29637
rect 30929 29597 30941 29631
rect 30975 29628 30987 29631
rect 32401 29631 32459 29637
rect 32401 29628 32413 29631
rect 30975 29600 32413 29628
rect 30975 29597 30987 29600
rect 30929 29591 30987 29597
rect 32401 29597 32413 29600
rect 32447 29597 32459 29631
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 32401 29591 32459 29597
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 31018 29560 31024 29572
rect 30576 29532 31024 29560
rect 29917 29523 29975 29529
rect 29932 29492 29960 29523
rect 31018 29520 31024 29532
rect 31076 29520 31082 29572
rect 32674 29560 32680 29572
rect 32635 29532 32680 29560
rect 32674 29520 32680 29532
rect 32732 29520 32738 29572
rect 33686 29520 33692 29572
rect 33744 29520 33750 29572
rect 30190 29492 30196 29504
rect 29748 29464 29960 29492
rect 30151 29464 30196 29492
rect 28369 29455 28427 29461
rect 30190 29452 30196 29464
rect 30248 29452 30254 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 17954 29288 17960 29300
rect 17144 29260 17960 29288
rect 17144 29220 17172 29260
rect 17954 29248 17960 29260
rect 18012 29288 18018 29300
rect 18966 29288 18972 29300
rect 18012 29260 18972 29288
rect 18012 29248 18018 29260
rect 18966 29248 18972 29260
rect 19024 29248 19030 29300
rect 20438 29288 20444 29300
rect 20351 29260 20444 29288
rect 17052 29192 17172 29220
rect 17052 29161 17080 29192
rect 18322 29180 18328 29232
rect 18380 29180 18386 29232
rect 20364 29229 20392 29260
rect 20438 29248 20444 29260
rect 20496 29288 20502 29300
rect 22646 29288 22652 29300
rect 20496 29260 22652 29288
rect 20496 29248 20502 29260
rect 22646 29248 22652 29260
rect 22704 29288 22710 29300
rect 24397 29291 24455 29297
rect 22704 29260 24348 29288
rect 22704 29248 22710 29260
rect 20349 29223 20407 29229
rect 20349 29189 20361 29223
rect 20395 29189 20407 29223
rect 20349 29183 20407 29189
rect 21634 29180 21640 29232
rect 21692 29220 21698 29232
rect 21821 29223 21879 29229
rect 21821 29220 21833 29223
rect 21692 29192 21833 29220
rect 21692 29180 21698 29192
rect 21821 29189 21833 29192
rect 21867 29189 21879 29223
rect 21821 29183 21879 29189
rect 22741 29223 22799 29229
rect 22741 29189 22753 29223
rect 22787 29220 22799 29223
rect 23750 29220 23756 29232
rect 22787 29192 23756 29220
rect 22787 29189 22799 29192
rect 22741 29183 22799 29189
rect 23750 29180 23756 29192
rect 23808 29180 23814 29232
rect 24320 29220 24348 29260
rect 24397 29257 24409 29291
rect 24443 29288 24455 29291
rect 25406 29288 25412 29300
rect 24443 29260 25412 29288
rect 24443 29257 24455 29260
rect 24397 29251 24455 29257
rect 25406 29248 25412 29260
rect 25464 29248 25470 29300
rect 25682 29248 25688 29300
rect 25740 29288 25746 29300
rect 26145 29291 26203 29297
rect 26145 29288 26157 29291
rect 25740 29260 26157 29288
rect 25740 29248 25746 29260
rect 26145 29257 26157 29260
rect 26191 29288 26203 29291
rect 26326 29288 26332 29300
rect 26191 29260 26332 29288
rect 26191 29257 26203 29260
rect 26145 29251 26203 29257
rect 26326 29248 26332 29260
rect 26384 29248 26390 29300
rect 29181 29291 29239 29297
rect 29181 29257 29193 29291
rect 29227 29288 29239 29291
rect 29638 29288 29644 29300
rect 29227 29260 29644 29288
rect 29227 29257 29239 29260
rect 29181 29251 29239 29257
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 43990 29288 43996 29300
rect 29748 29260 43996 29288
rect 29748 29220 29776 29260
rect 43990 29248 43996 29260
rect 44048 29248 44054 29300
rect 30006 29220 30012 29232
rect 24320 29192 26188 29220
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 19886 29112 19892 29164
rect 19944 29152 19950 29164
rect 20073 29155 20131 29161
rect 20073 29152 20085 29155
rect 19944 29124 20085 29152
rect 19944 29112 19950 29124
rect 20073 29121 20085 29124
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29152 20499 29155
rect 20530 29152 20536 29164
rect 20487 29124 20536 29152
rect 20487 29121 20499 29124
rect 20441 29115 20499 29121
rect 14274 29084 14280 29096
rect 14235 29056 14280 29084
rect 14274 29044 14280 29056
rect 14332 29044 14338 29096
rect 14458 29084 14464 29096
rect 14419 29056 14464 29084
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 14737 29087 14795 29093
rect 14737 29053 14749 29087
rect 14783 29053 14795 29087
rect 17310 29084 17316 29096
rect 17271 29056 17316 29084
rect 14737 29047 14795 29053
rect 8294 28976 8300 29028
rect 8352 29016 8358 29028
rect 14752 29016 14780 29047
rect 17310 29044 17316 29056
rect 17368 29044 17374 29096
rect 20272 29084 20300 29115
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29152 22063 29155
rect 22554 29152 22560 29164
rect 22051 29124 22560 29152
rect 22051 29121 22063 29124
rect 22005 29115 22063 29121
rect 22554 29112 22560 29124
rect 22612 29152 22618 29164
rect 22922 29152 22928 29164
rect 22612 29124 22928 29152
rect 22612 29112 22618 29124
rect 22922 29112 22928 29124
rect 22980 29112 22986 29164
rect 23566 29152 23572 29164
rect 23527 29124 23572 29152
rect 23566 29112 23572 29124
rect 23624 29112 23630 29164
rect 23934 29112 23940 29164
rect 23992 29152 23998 29164
rect 24305 29155 24363 29161
rect 24305 29152 24317 29155
rect 23992 29124 24317 29152
rect 23992 29112 23998 29124
rect 24305 29121 24317 29124
rect 24351 29121 24363 29155
rect 24305 29115 24363 29121
rect 24854 29112 24860 29164
rect 24912 29152 24918 29164
rect 25409 29155 25467 29161
rect 25409 29152 25421 29155
rect 24912 29124 25421 29152
rect 24912 29112 24918 29124
rect 25409 29121 25421 29124
rect 25455 29152 25467 29155
rect 25498 29152 25504 29164
rect 25455 29124 25504 29152
rect 25455 29121 25467 29124
rect 25409 29115 25467 29121
rect 25498 29112 25504 29124
rect 25556 29112 25562 29164
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29121 26111 29155
rect 26053 29115 26111 29121
rect 20898 29084 20904 29096
rect 20272 29056 20904 29084
rect 20898 29044 20904 29056
rect 20956 29044 20962 29096
rect 21082 29044 21088 29096
rect 21140 29084 21146 29096
rect 22189 29087 22247 29093
rect 22189 29084 22201 29087
rect 21140 29056 22201 29084
rect 21140 29044 21146 29056
rect 22189 29053 22201 29056
rect 22235 29053 22247 29087
rect 22189 29047 22247 29053
rect 24578 29044 24584 29096
rect 24636 29084 24642 29096
rect 26068 29084 26096 29115
rect 24636 29056 26096 29084
rect 26160 29084 26188 29192
rect 27172 29192 29776 29220
rect 29840 29192 30012 29220
rect 27172 29161 27200 29192
rect 29840 29164 29868 29192
rect 30006 29180 30012 29192
rect 30064 29180 30070 29232
rect 30101 29223 30159 29229
rect 30101 29189 30113 29223
rect 30147 29220 30159 29223
rect 30190 29220 30196 29232
rect 30147 29192 30196 29220
rect 30147 29189 30159 29192
rect 30101 29183 30159 29189
rect 30190 29180 30196 29192
rect 30248 29180 30254 29232
rect 32674 29180 32680 29232
rect 32732 29220 32738 29232
rect 33137 29223 33195 29229
rect 33137 29220 33149 29223
rect 32732 29192 33149 29220
rect 32732 29180 32738 29192
rect 33137 29189 33149 29192
rect 33183 29189 33195 29223
rect 33137 29183 33195 29189
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 27249 29155 27307 29161
rect 27249 29121 27261 29155
rect 27295 29121 27307 29155
rect 27430 29152 27436 29164
rect 27391 29124 27436 29152
rect 27249 29115 27307 29121
rect 27264 29084 27292 29115
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 27522 29112 27528 29164
rect 27580 29152 27586 29164
rect 27580 29124 27625 29152
rect 27580 29112 27586 29124
rect 28166 29112 28172 29164
rect 28224 29152 28230 29164
rect 28534 29152 28540 29164
rect 28224 29124 28540 29152
rect 28224 29112 28230 29124
rect 28534 29112 28540 29124
rect 28592 29152 28598 29164
rect 28813 29155 28871 29161
rect 28813 29152 28825 29155
rect 28592 29124 28825 29152
rect 28592 29112 28598 29124
rect 28813 29121 28825 29124
rect 28859 29121 28871 29155
rect 29822 29152 29828 29164
rect 29735 29124 29828 29152
rect 28813 29115 28871 29121
rect 27614 29084 27620 29096
rect 26160 29056 27620 29084
rect 24636 29044 24642 29056
rect 27614 29044 27620 29056
rect 27672 29044 27678 29096
rect 28718 29084 28724 29096
rect 28679 29056 28724 29084
rect 28718 29044 28724 29056
rect 28776 29044 28782 29096
rect 8352 28988 14780 29016
rect 8352 28976 8358 28988
rect 18966 28976 18972 29028
rect 19024 29016 19030 29028
rect 22925 29019 22983 29025
rect 22925 29016 22937 29019
rect 19024 28988 22937 29016
rect 19024 28976 19030 28988
rect 22925 28985 22937 28988
rect 22971 29016 22983 29019
rect 23290 29016 23296 29028
rect 22971 28988 23296 29016
rect 22971 28985 22983 28988
rect 22925 28979 22983 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23474 28976 23480 29028
rect 23532 29016 23538 29028
rect 23753 29019 23811 29025
rect 23753 29016 23765 29019
rect 23532 28988 23765 29016
rect 23532 28976 23538 28988
rect 23753 28985 23765 28988
rect 23799 29016 23811 29019
rect 23842 29016 23848 29028
rect 23799 28988 23848 29016
rect 23799 28985 23811 28988
rect 23753 28979 23811 28985
rect 23842 28976 23848 28988
rect 23900 28976 23906 29028
rect 25590 29016 25596 29028
rect 25503 28988 25596 29016
rect 25590 28976 25596 28988
rect 25648 29016 25654 29028
rect 28828 29016 28856 29115
rect 29822 29112 29828 29124
rect 29880 29112 29886 29164
rect 31202 29112 31208 29164
rect 31260 29112 31266 29164
rect 32398 29152 32404 29164
rect 32359 29124 32404 29152
rect 32398 29112 32404 29124
rect 32456 29112 32462 29164
rect 32582 29152 32588 29164
rect 32543 29124 32588 29152
rect 32582 29112 32588 29124
rect 32640 29112 32646 29164
rect 32858 29112 32864 29164
rect 32916 29152 32922 29164
rect 32953 29155 33011 29161
rect 32953 29152 32965 29155
rect 32916 29124 32965 29152
rect 32916 29112 32922 29124
rect 32953 29121 32965 29124
rect 32999 29121 33011 29155
rect 32953 29115 33011 29121
rect 31573 29087 31631 29093
rect 31573 29084 31585 29087
rect 29932 29056 31585 29084
rect 29932 29016 29960 29056
rect 31573 29053 31585 29056
rect 31619 29053 31631 29087
rect 31573 29047 31631 29053
rect 32490 29044 32496 29096
rect 32548 29084 32554 29096
rect 32677 29087 32735 29093
rect 32677 29084 32689 29087
rect 32548 29056 32689 29084
rect 32548 29044 32554 29056
rect 32677 29053 32689 29056
rect 32723 29053 32735 29087
rect 32677 29047 32735 29053
rect 32766 29044 32772 29096
rect 32824 29084 32830 29096
rect 32824 29056 32869 29084
rect 32824 29044 32830 29056
rect 25648 28988 27108 29016
rect 28828 28988 29960 29016
rect 25648 28976 25654 28988
rect 18782 28948 18788 28960
rect 18743 28920 18788 28948
rect 18782 28908 18788 28920
rect 18840 28948 18846 28960
rect 20530 28948 20536 28960
rect 18840 28920 20536 28948
rect 18840 28908 18846 28920
rect 20530 28908 20536 28920
rect 20588 28908 20594 28960
rect 20625 28951 20683 28957
rect 20625 28917 20637 28951
rect 20671 28948 20683 28951
rect 22002 28948 22008 28960
rect 20671 28920 22008 28948
rect 20671 28917 20683 28920
rect 20625 28911 20683 28917
rect 22002 28908 22008 28920
rect 22060 28908 22066 28960
rect 26602 28908 26608 28960
rect 26660 28948 26666 28960
rect 26973 28951 27031 28957
rect 26973 28948 26985 28951
rect 26660 28920 26985 28948
rect 26660 28908 26666 28920
rect 26973 28917 26985 28920
rect 27019 28917 27031 28951
rect 27080 28948 27108 28988
rect 29086 28948 29092 28960
rect 27080 28920 29092 28948
rect 26973 28911 27031 28917
rect 29086 28908 29092 28920
rect 29144 28908 29150 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1854 28704 1860 28756
rect 1912 28744 1918 28756
rect 1912 28716 6914 28744
rect 1912 28704 1918 28716
rect 6886 28676 6914 28716
rect 14458 28704 14464 28756
rect 14516 28744 14522 28756
rect 14737 28747 14795 28753
rect 14737 28744 14749 28747
rect 14516 28716 14749 28744
rect 14516 28704 14522 28716
rect 14737 28713 14749 28716
rect 14783 28713 14795 28747
rect 14737 28707 14795 28713
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 18417 28747 18475 28753
rect 18417 28744 18429 28747
rect 17368 28716 18429 28744
rect 17368 28704 17374 28716
rect 18417 28713 18429 28716
rect 18463 28713 18475 28747
rect 18417 28707 18475 28713
rect 20438 28704 20444 28756
rect 20496 28744 20502 28756
rect 21082 28744 21088 28756
rect 20496 28716 21088 28744
rect 20496 28704 20502 28716
rect 21082 28704 21088 28716
rect 21140 28744 21146 28756
rect 21269 28747 21327 28753
rect 21269 28744 21281 28747
rect 21140 28716 21281 28744
rect 21140 28704 21146 28716
rect 21269 28713 21281 28716
rect 21315 28713 21327 28747
rect 21269 28707 21327 28713
rect 25498 28704 25504 28756
rect 25556 28744 25562 28756
rect 28537 28747 28595 28753
rect 28537 28744 28549 28747
rect 25556 28716 28549 28744
rect 25556 28704 25562 28716
rect 28537 28713 28549 28716
rect 28583 28713 28595 28747
rect 28537 28707 28595 28713
rect 31202 28704 31208 28756
rect 31260 28744 31266 28756
rect 31297 28747 31355 28753
rect 31297 28744 31309 28747
rect 31260 28716 31309 28744
rect 31260 28704 31266 28716
rect 31297 28713 31309 28716
rect 31343 28713 31355 28747
rect 31297 28707 31355 28713
rect 19978 28676 19984 28688
rect 6886 28648 19984 28676
rect 19978 28636 19984 28648
rect 20036 28636 20042 28688
rect 26234 28676 26240 28688
rect 25056 28648 26240 28676
rect 15841 28611 15899 28617
rect 15841 28608 15853 28611
rect 6886 28580 15853 28608
rect 3142 28432 3148 28484
rect 3200 28472 3206 28484
rect 6886 28472 6914 28580
rect 15841 28577 15853 28580
rect 15887 28577 15899 28611
rect 15841 28571 15899 28577
rect 17957 28611 18015 28617
rect 17957 28577 17969 28611
rect 18003 28608 18015 28611
rect 18782 28608 18788 28620
rect 18003 28580 18788 28608
rect 18003 28577 18015 28580
rect 17957 28571 18015 28577
rect 18782 28568 18788 28580
rect 18840 28568 18846 28620
rect 20165 28611 20223 28617
rect 20165 28577 20177 28611
rect 20211 28608 20223 28611
rect 20438 28608 20444 28620
rect 20211 28580 20444 28608
rect 20211 28577 20223 28580
rect 20165 28571 20223 28577
rect 20438 28568 20444 28580
rect 20496 28568 20502 28620
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 20640 28580 21373 28608
rect 20640 28552 20668 28580
rect 21361 28577 21373 28580
rect 21407 28577 21419 28611
rect 23474 28608 23480 28620
rect 21361 28571 21419 28577
rect 22204 28580 23480 28608
rect 14642 28540 14648 28552
rect 14603 28512 14648 28540
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 15378 28540 15384 28552
rect 15339 28512 15384 28540
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 17678 28540 17684 28552
rect 17639 28512 17684 28540
rect 17678 28500 17684 28512
rect 17736 28500 17742 28552
rect 17862 28540 17868 28552
rect 17823 28512 17868 28540
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 18049 28543 18107 28549
rect 18049 28518 18061 28543
rect 17972 28509 18061 28518
rect 18095 28509 18107 28543
rect 18230 28540 18236 28552
rect 18191 28512 18236 28540
rect 17972 28503 18107 28509
rect 17972 28490 18092 28503
rect 18230 28500 18236 28512
rect 18288 28500 18294 28552
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 20073 28543 20131 28549
rect 20073 28540 20085 28543
rect 19944 28512 20085 28540
rect 19944 28500 19950 28512
rect 20073 28509 20085 28512
rect 20119 28540 20131 28543
rect 20622 28540 20628 28552
rect 20119 28512 20628 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20714 28500 20720 28552
rect 20772 28540 20778 28552
rect 21085 28543 21143 28549
rect 21085 28540 21097 28543
rect 20772 28512 21097 28540
rect 20772 28500 20778 28512
rect 21085 28509 21097 28512
rect 21131 28509 21143 28543
rect 22002 28540 22008 28552
rect 21963 28512 22008 28540
rect 21085 28503 21143 28509
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 22204 28549 22232 28580
rect 23474 28568 23480 28580
rect 23532 28568 23538 28620
rect 24302 28568 24308 28620
rect 24360 28608 24366 28620
rect 25056 28617 25084 28648
rect 26234 28636 26240 28648
rect 26292 28636 26298 28688
rect 26786 28676 26792 28688
rect 26747 28648 26792 28676
rect 26786 28636 26792 28648
rect 26844 28636 26850 28688
rect 24857 28611 24915 28617
rect 24857 28608 24869 28611
rect 24360 28580 24869 28608
rect 24360 28568 24366 28580
rect 24857 28577 24869 28580
rect 24903 28577 24915 28611
rect 24857 28571 24915 28577
rect 25041 28611 25099 28617
rect 25041 28577 25053 28611
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28509 22247 28543
rect 22189 28503 22247 28509
rect 22281 28543 22339 28549
rect 22281 28509 22293 28543
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28509 23443 28543
rect 23385 28503 23443 28509
rect 15562 28472 15568 28484
rect 3200 28444 6914 28472
rect 15523 28444 15568 28472
rect 3200 28432 3206 28444
rect 15562 28432 15568 28444
rect 15620 28432 15626 28484
rect 7834 28364 7840 28416
rect 7892 28404 7898 28416
rect 17972 28404 18000 28490
rect 18138 28432 18144 28484
rect 18196 28472 18202 28484
rect 19334 28472 19340 28484
rect 18196 28444 19340 28472
rect 18196 28432 18202 28444
rect 19334 28432 19340 28444
rect 19392 28432 19398 28484
rect 22296 28472 22324 28503
rect 20456 28444 22324 28472
rect 23400 28472 23428 28503
rect 23566 28500 23572 28552
rect 23624 28540 23630 28552
rect 23661 28543 23719 28549
rect 23661 28540 23673 28543
rect 23624 28512 23673 28540
rect 23624 28500 23630 28512
rect 23661 28509 23673 28512
rect 23707 28509 23719 28543
rect 24762 28540 24768 28552
rect 24723 28512 24768 28540
rect 23661 28503 23719 28509
rect 24762 28500 24768 28512
rect 24820 28500 24826 28552
rect 24872 28472 24900 28571
rect 25406 28568 25412 28620
rect 25464 28608 25470 28620
rect 27430 28608 27436 28620
rect 25464 28580 25820 28608
rect 25464 28568 25470 28580
rect 25682 28540 25688 28552
rect 25643 28512 25688 28540
rect 25682 28500 25688 28512
rect 25740 28500 25746 28552
rect 25792 28549 25820 28580
rect 25884 28580 27436 28608
rect 25777 28543 25835 28549
rect 25777 28509 25789 28543
rect 25823 28509 25835 28543
rect 25777 28503 25835 28509
rect 25884 28472 25912 28580
rect 27430 28568 27436 28580
rect 27488 28608 27494 28620
rect 27617 28611 27675 28617
rect 27617 28608 27629 28611
rect 27488 28580 27629 28608
rect 27488 28568 27494 28580
rect 27617 28577 27629 28580
rect 27663 28577 27675 28611
rect 27617 28571 27675 28577
rect 26602 28540 26608 28552
rect 26563 28512 26608 28540
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 26878 28500 26884 28552
rect 26936 28540 26942 28552
rect 26936 28512 26981 28540
rect 26936 28500 26942 28512
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 28353 28543 28411 28549
rect 28353 28540 28365 28543
rect 27764 28512 28365 28540
rect 27764 28500 27770 28512
rect 28353 28509 28365 28512
rect 28399 28540 28411 28543
rect 28718 28540 28724 28552
rect 28399 28512 28724 28540
rect 28399 28509 28411 28512
rect 28353 28503 28411 28509
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 30926 28500 30932 28552
rect 30984 28540 30990 28552
rect 31205 28543 31263 28549
rect 31205 28540 31217 28543
rect 30984 28512 31217 28540
rect 30984 28500 30990 28512
rect 31205 28509 31217 28512
rect 31251 28509 31263 28543
rect 31205 28503 31263 28509
rect 23400 28444 24440 28472
rect 24872 28444 25912 28472
rect 25961 28475 26019 28481
rect 20456 28413 20484 28444
rect 7892 28376 18000 28404
rect 20441 28407 20499 28413
rect 7892 28364 7898 28376
rect 20441 28373 20453 28407
rect 20487 28373 20499 28407
rect 20898 28404 20904 28416
rect 20859 28376 20904 28404
rect 20441 28367 20499 28373
rect 20898 28364 20904 28376
rect 20956 28364 20962 28416
rect 21818 28404 21824 28416
rect 21779 28376 21824 28404
rect 21818 28364 21824 28376
rect 21876 28364 21882 28416
rect 23201 28407 23259 28413
rect 23201 28373 23213 28407
rect 23247 28404 23259 28407
rect 23474 28404 23480 28416
rect 23247 28376 23480 28404
rect 23247 28373 23259 28376
rect 23201 28367 23259 28373
rect 23474 28364 23480 28376
rect 23532 28364 23538 28416
rect 23566 28364 23572 28416
rect 23624 28404 23630 28416
rect 24210 28404 24216 28416
rect 23624 28376 24216 28404
rect 23624 28364 23630 28376
rect 24210 28364 24216 28376
rect 24268 28364 24274 28416
rect 24412 28413 24440 28444
rect 25961 28441 25973 28475
rect 26007 28472 26019 28475
rect 27154 28472 27160 28484
rect 26007 28444 27160 28472
rect 26007 28441 26019 28444
rect 25961 28435 26019 28441
rect 27154 28432 27160 28444
rect 27212 28472 27218 28484
rect 27433 28475 27491 28481
rect 27433 28472 27445 28475
rect 27212 28444 27445 28472
rect 27212 28432 27218 28444
rect 27433 28441 27445 28444
rect 27479 28441 27491 28475
rect 28166 28472 28172 28484
rect 28127 28444 28172 28472
rect 27433 28435 27491 28441
rect 28166 28432 28172 28444
rect 28224 28432 28230 28484
rect 24397 28407 24455 28413
rect 24397 28373 24409 28407
rect 24443 28373 24455 28407
rect 26418 28404 26424 28416
rect 26379 28376 26424 28404
rect 24397 28367 24455 28373
rect 26418 28364 26424 28376
rect 26476 28364 26482 28416
rect 28442 28364 28448 28416
rect 28500 28404 28506 28416
rect 32490 28404 32496 28416
rect 28500 28376 32496 28404
rect 28500 28364 28506 28376
rect 32490 28364 32496 28376
rect 32548 28364 32554 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 15562 28200 15568 28212
rect 15523 28172 15568 28200
rect 15562 28160 15568 28172
rect 15620 28160 15626 28212
rect 21818 28200 21824 28212
rect 19260 28172 21824 28200
rect 14182 28132 14188 28144
rect 13754 28104 14188 28132
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 18138 28132 18144 28144
rect 14700 28104 18144 28132
rect 14700 28092 14706 28104
rect 15488 28073 15516 28104
rect 18138 28092 18144 28104
rect 18196 28092 18202 28144
rect 19260 28141 19288 28172
rect 21818 28160 21824 28172
rect 21876 28160 21882 28212
rect 27157 28203 27215 28209
rect 27157 28169 27169 28203
rect 27203 28200 27215 28203
rect 28077 28203 28135 28209
rect 28077 28200 28089 28203
rect 27203 28172 28089 28200
rect 27203 28169 27215 28172
rect 27157 28163 27215 28169
rect 28077 28169 28089 28172
rect 28123 28169 28135 28203
rect 28077 28163 28135 28169
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28101 19303 28135
rect 19245 28095 19303 28101
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 22922 28132 22928 28144
rect 19392 28104 19734 28132
rect 22066 28104 22784 28132
rect 22883 28104 22928 28132
rect 19392 28092 19398 28104
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28033 15531 28067
rect 18966 28064 18972 28076
rect 18927 28036 18972 28064
rect 15473 28027 15531 28033
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 21821 28067 21879 28073
rect 21821 28033 21833 28067
rect 21867 28064 21879 28067
rect 22066 28064 22094 28104
rect 22646 28064 22652 28076
rect 21867 28036 22094 28064
rect 22607 28036 22652 28064
rect 21867 28033 21879 28036
rect 21821 28027 21879 28033
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 22756 28064 22784 28104
rect 22922 28092 22928 28104
rect 22980 28092 22986 28144
rect 24026 28132 24032 28144
rect 23768 28104 24032 28132
rect 23768 28076 23796 28104
rect 24026 28092 24032 28104
rect 24084 28092 24090 28144
rect 28092 28132 28120 28163
rect 28166 28160 28172 28212
rect 28224 28200 28230 28212
rect 28997 28203 29055 28209
rect 28997 28200 29009 28203
rect 28224 28172 29009 28200
rect 28224 28160 28230 28172
rect 28997 28169 29009 28172
rect 29043 28169 29055 28203
rect 28997 28163 29055 28169
rect 29086 28160 29092 28212
rect 29144 28200 29150 28212
rect 31205 28203 31263 28209
rect 31205 28200 31217 28203
rect 29144 28172 31217 28200
rect 29144 28160 29150 28172
rect 31205 28169 31217 28172
rect 31251 28169 31263 28203
rect 31205 28163 31263 28169
rect 28626 28132 28632 28144
rect 28092 28104 28632 28132
rect 28626 28092 28632 28104
rect 28684 28132 28690 28144
rect 30282 28132 30288 28144
rect 28684 28104 29684 28132
rect 30243 28104 30288 28132
rect 28684 28092 28690 28104
rect 23750 28064 23756 28076
rect 22756 28036 23756 28064
rect 23750 28024 23756 28036
rect 23808 28024 23814 28076
rect 23934 28064 23940 28076
rect 23895 28036 23940 28064
rect 23934 28024 23940 28036
rect 23992 28024 23998 28076
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28064 24179 28067
rect 24578 28064 24584 28076
rect 24167 28036 24584 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 24578 28024 24584 28036
rect 24636 28064 24642 28076
rect 24762 28064 24768 28076
rect 24636 28036 24768 28064
rect 24636 28024 24642 28036
rect 24762 28024 24768 28036
rect 24820 28024 24826 28076
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 26510 28064 26516 28076
rect 26283 28036 26516 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 26510 28024 26516 28036
rect 26568 28024 26574 28076
rect 26970 28064 26976 28076
rect 26931 28036 26976 28064
rect 26970 28024 26976 28036
rect 27028 28024 27034 28076
rect 27249 28067 27307 28073
rect 27249 28033 27261 28067
rect 27295 28064 27307 28067
rect 27614 28064 27620 28076
rect 27295 28036 27620 28064
rect 27295 28033 27307 28036
rect 27249 28027 27307 28033
rect 27614 28024 27620 28036
rect 27672 28024 27678 28076
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 28534 28064 28540 28076
rect 27764 28036 27809 28064
rect 28495 28036 28540 28064
rect 27764 28024 27770 28036
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 29656 28073 29684 28104
rect 30282 28092 30288 28104
rect 30340 28092 30346 28144
rect 30469 28135 30527 28141
rect 30469 28132 30481 28135
rect 30392 28104 30481 28132
rect 28813 28067 28871 28073
rect 28813 28033 28825 28067
rect 28859 28064 28871 28067
rect 29641 28067 29699 28073
rect 28859 28036 29592 28064
rect 28859 28033 28871 28036
rect 28813 28027 28871 28033
rect 12250 27996 12256 28008
rect 12211 27968 12256 27996
rect 12250 27956 12256 27968
rect 12308 27956 12314 28008
rect 12526 27996 12532 28008
rect 12487 27968 12532 27996
rect 12526 27956 12532 27968
rect 12584 27956 12590 28008
rect 14001 27999 14059 28005
rect 14001 27965 14013 27999
rect 14047 27996 14059 27999
rect 14550 27996 14556 28008
rect 14047 27968 14556 27996
rect 14047 27965 14059 27968
rect 14001 27959 14059 27965
rect 14550 27956 14556 27968
rect 14608 27996 14614 28008
rect 16669 27999 16727 28005
rect 16669 27996 16681 27999
rect 14608 27968 16681 27996
rect 14608 27956 14614 27968
rect 16669 27965 16681 27968
rect 16715 27965 16727 27999
rect 16850 27996 16856 28008
rect 16811 27968 16856 27996
rect 16669 27959 16727 27965
rect 16850 27956 16856 27968
rect 16908 27956 16914 28008
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27965 17187 27999
rect 17129 27959 17187 27965
rect 16574 27888 16580 27940
rect 16632 27928 16638 27940
rect 17144 27928 17172 27959
rect 17678 27956 17684 28008
rect 17736 27996 17742 28008
rect 17736 27968 20300 27996
rect 17736 27956 17742 27968
rect 16632 27900 17172 27928
rect 20272 27928 20300 27968
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 20717 27999 20775 28005
rect 20717 27996 20729 27999
rect 20680 27968 20729 27996
rect 20680 27956 20686 27968
rect 20717 27965 20729 27968
rect 20763 27965 20775 27999
rect 20717 27959 20775 27965
rect 21913 27999 21971 28005
rect 21913 27965 21925 27999
rect 21959 27996 21971 27999
rect 21959 27968 22876 27996
rect 21959 27965 21971 27968
rect 21913 27959 21971 27965
rect 22189 27931 22247 27937
rect 22189 27928 22201 27931
rect 20272 27900 22201 27928
rect 16632 27888 16638 27900
rect 22189 27897 22201 27900
rect 22235 27897 22247 27931
rect 22738 27928 22744 27940
rect 22699 27900 22744 27928
rect 22189 27891 22247 27897
rect 22738 27888 22744 27900
rect 22796 27888 22802 27940
rect 22848 27872 22876 27968
rect 26878 27956 26884 28008
rect 26936 27996 26942 28008
rect 27801 27999 27859 28005
rect 27801 27996 27813 27999
rect 26936 27968 27813 27996
rect 26936 27956 26942 27968
rect 27801 27965 27813 27968
rect 27847 27996 27859 27999
rect 28629 27999 28687 28005
rect 28629 27996 28641 27999
rect 27847 27968 28641 27996
rect 27847 27965 27859 27968
rect 27801 27959 27859 27965
rect 28629 27965 28641 27968
rect 28675 27965 28687 27999
rect 28629 27959 28687 27965
rect 28902 27956 28908 28008
rect 28960 27996 28966 28008
rect 29457 27999 29515 28005
rect 29457 27996 29469 27999
rect 28960 27968 29469 27996
rect 28960 27956 28966 27968
rect 29457 27965 29469 27968
rect 29503 27965 29515 27999
rect 29564 27996 29592 28036
rect 29641 28033 29653 28067
rect 29687 28033 29699 28067
rect 29641 28027 29699 28033
rect 30392 28008 30420 28104
rect 30469 28101 30481 28104
rect 30515 28101 30527 28135
rect 30469 28095 30527 28101
rect 31021 28135 31079 28141
rect 31021 28101 31033 28135
rect 31067 28132 31079 28135
rect 32195 28135 32253 28141
rect 32195 28132 32207 28135
rect 31067 28104 32207 28132
rect 31067 28101 31079 28104
rect 31021 28095 31079 28101
rect 32195 28101 32207 28104
rect 32241 28101 32253 28135
rect 32195 28095 32253 28101
rect 30558 28024 30564 28076
rect 30616 28064 30622 28076
rect 31297 28067 31355 28073
rect 31297 28064 31309 28067
rect 30616 28036 30661 28064
rect 30944 28036 31309 28064
rect 30616 28024 30622 28036
rect 30374 27996 30380 28008
rect 29564 27968 30380 27996
rect 29457 27959 29515 27965
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 30944 27996 30972 28036
rect 31297 28033 31309 28036
rect 31343 28033 31355 28067
rect 32490 28064 32496 28076
rect 32451 28036 32496 28064
rect 31297 28027 31355 28033
rect 32490 28024 32496 28036
rect 32548 28024 32554 28076
rect 45922 28024 45928 28076
rect 45980 28064 45986 28076
rect 46753 28067 46811 28073
rect 46753 28064 46765 28067
rect 45980 28036 46765 28064
rect 45980 28024 45986 28036
rect 46753 28033 46765 28036
rect 46799 28033 46811 28067
rect 46753 28027 46811 28033
rect 30760 27968 30972 27996
rect 23658 27888 23664 27940
rect 23716 27928 23722 27940
rect 24305 27931 24363 27937
rect 24305 27928 24317 27931
rect 23716 27900 24317 27928
rect 23716 27888 23722 27900
rect 24305 27897 24317 27900
rect 24351 27928 24363 27931
rect 26973 27931 27031 27937
rect 24351 27900 26464 27928
rect 24351 27897 24363 27900
rect 24305 27891 24363 27897
rect 20898 27820 20904 27872
rect 20956 27860 20962 27872
rect 21821 27863 21879 27869
rect 21821 27860 21833 27863
rect 20956 27832 21833 27860
rect 20956 27820 20962 27832
rect 21821 27829 21833 27832
rect 21867 27829 21879 27863
rect 22830 27860 22836 27872
rect 22791 27832 22836 27860
rect 21821 27823 21879 27829
rect 22830 27820 22836 27832
rect 22888 27820 22894 27872
rect 26326 27860 26332 27872
rect 26287 27832 26332 27860
rect 26326 27820 26332 27832
rect 26384 27820 26390 27872
rect 26436 27860 26464 27900
rect 26973 27897 26985 27931
rect 27019 27928 27031 27931
rect 27522 27928 27528 27940
rect 27019 27900 27528 27928
rect 27019 27897 27031 27900
rect 26973 27891 27031 27897
rect 27522 27888 27528 27900
rect 27580 27888 27586 27940
rect 29914 27928 29920 27940
rect 27632 27900 29920 27928
rect 27632 27860 27660 27900
rect 29914 27888 29920 27900
rect 29972 27888 29978 27940
rect 30285 27931 30343 27937
rect 30285 27897 30297 27931
rect 30331 27928 30343 27931
rect 30760 27928 30788 27968
rect 31386 27956 31392 28008
rect 31444 27996 31450 28008
rect 32125 27999 32183 28005
rect 32125 27996 32137 27999
rect 31444 27968 32137 27996
rect 31444 27956 31450 27968
rect 32125 27965 32137 27968
rect 32171 27965 32183 27999
rect 32125 27959 32183 27965
rect 32214 27956 32220 28008
rect 32272 27996 32278 28008
rect 32309 27999 32367 28005
rect 32309 27996 32321 27999
rect 32272 27968 32321 27996
rect 32272 27956 32278 27968
rect 32309 27965 32321 27968
rect 32355 27965 32367 27999
rect 32309 27959 32367 27965
rect 30331 27900 30788 27928
rect 30331 27897 30343 27900
rect 30285 27891 30343 27897
rect 27890 27860 27896 27872
rect 26436 27832 27660 27860
rect 27803 27832 27896 27860
rect 27890 27820 27896 27832
rect 27948 27860 27954 27872
rect 28534 27860 28540 27872
rect 27948 27832 28540 27860
rect 27948 27820 27954 27832
rect 28534 27820 28540 27832
rect 28592 27820 28598 27872
rect 28813 27863 28871 27869
rect 28813 27829 28825 27863
rect 28859 27860 28871 27863
rect 28902 27860 28908 27872
rect 28859 27832 28908 27860
rect 28859 27829 28871 27832
rect 28813 27823 28871 27829
rect 28902 27820 28908 27832
rect 28960 27820 28966 27872
rect 29730 27820 29736 27872
rect 29788 27860 29794 27872
rect 29825 27863 29883 27869
rect 29825 27860 29837 27863
rect 29788 27832 29837 27860
rect 29788 27820 29794 27832
rect 29825 27829 29837 27832
rect 29871 27829 29883 27863
rect 31018 27860 31024 27872
rect 30979 27832 31024 27860
rect 29825 27823 29883 27829
rect 31018 27820 31024 27832
rect 31076 27820 31082 27872
rect 32398 27820 32404 27872
rect 32456 27860 32462 27872
rect 32456 27832 32501 27860
rect 32456 27820 32462 27832
rect 46474 27820 46480 27872
rect 46532 27860 46538 27872
rect 46845 27863 46903 27869
rect 46845 27860 46857 27863
rect 46532 27832 46857 27860
rect 46532 27820 46538 27832
rect 46845 27829 46857 27832
rect 46891 27829 46903 27863
rect 46845 27823 46903 27829
rect 47026 27820 47032 27872
rect 47084 27860 47090 27872
rect 47765 27863 47823 27869
rect 47765 27860 47777 27863
rect 47084 27832 47777 27860
rect 47084 27820 47090 27832
rect 47765 27829 47777 27832
rect 47811 27829 47823 27863
rect 47765 27823 47823 27829
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 11517 27659 11575 27665
rect 11517 27625 11529 27659
rect 11563 27656 11575 27659
rect 12250 27656 12256 27668
rect 11563 27628 12256 27656
rect 11563 27625 11575 27628
rect 11517 27619 11575 27625
rect 12250 27616 12256 27628
rect 12308 27616 12314 27668
rect 12526 27656 12532 27668
rect 12487 27628 12532 27656
rect 12526 27616 12532 27628
rect 12584 27616 12590 27668
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 17221 27659 17279 27665
rect 17221 27656 17233 27659
rect 16908 27628 17233 27656
rect 16908 27616 16914 27628
rect 17221 27625 17233 27628
rect 17267 27625 17279 27659
rect 17221 27619 17279 27625
rect 25764 27659 25822 27665
rect 25764 27625 25776 27659
rect 25810 27656 25822 27659
rect 26418 27656 26424 27668
rect 25810 27628 26424 27656
rect 25810 27625 25822 27628
rect 25764 27619 25822 27625
rect 26418 27616 26424 27628
rect 26476 27616 26482 27668
rect 26878 27616 26884 27668
rect 26936 27656 26942 27668
rect 27249 27659 27307 27665
rect 27249 27656 27261 27659
rect 26936 27628 27261 27656
rect 26936 27616 26942 27628
rect 27249 27625 27261 27628
rect 27295 27656 27307 27659
rect 29914 27656 29920 27668
rect 27295 27628 28028 27656
rect 29875 27628 29920 27656
rect 27295 27625 27307 27628
rect 27249 27619 27307 27625
rect 14182 27588 14188 27600
rect 14143 27560 14188 27588
rect 14182 27548 14188 27560
rect 14240 27548 14246 27600
rect 18233 27591 18291 27597
rect 18233 27557 18245 27591
rect 18279 27588 18291 27591
rect 18322 27588 18328 27600
rect 18279 27560 18328 27588
rect 18279 27557 18291 27560
rect 18233 27551 18291 27557
rect 18322 27548 18328 27560
rect 18380 27548 18386 27600
rect 19334 27588 19340 27600
rect 19295 27560 19340 27588
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 21634 27548 21640 27600
rect 21692 27588 21698 27600
rect 21910 27588 21916 27600
rect 21692 27560 21916 27588
rect 21692 27548 21698 27560
rect 21910 27548 21916 27560
rect 21968 27588 21974 27600
rect 22738 27588 22744 27600
rect 21968 27560 22744 27588
rect 21968 27548 21974 27560
rect 22738 27548 22744 27560
rect 22796 27548 22802 27600
rect 27614 27548 27620 27600
rect 27672 27588 27678 27600
rect 27893 27591 27951 27597
rect 27893 27588 27905 27591
rect 27672 27560 27905 27588
rect 27672 27548 27678 27560
rect 27893 27557 27905 27560
rect 27939 27557 27951 27591
rect 27893 27551 27951 27557
rect 12345 27523 12403 27529
rect 12345 27489 12357 27523
rect 12391 27520 12403 27523
rect 13173 27523 13231 27529
rect 13173 27520 13185 27523
rect 12391 27492 13185 27520
rect 12391 27489 12403 27492
rect 12345 27483 12403 27489
rect 13173 27489 13185 27492
rect 13219 27489 13231 27523
rect 16482 27520 16488 27532
rect 13173 27483 13231 27489
rect 13280 27492 14688 27520
rect 16443 27492 16488 27520
rect 13280 27464 13308 27492
rect 14660 27464 14688 27492
rect 16482 27480 16488 27492
rect 16540 27480 16546 27532
rect 20622 27520 20628 27532
rect 20456 27492 20628 27520
rect 11422 27452 11428 27464
rect 11383 27424 11428 27452
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 12253 27455 12311 27461
rect 12253 27421 12265 27455
rect 12299 27421 12311 27455
rect 12253 27415 12311 27421
rect 13081 27455 13139 27461
rect 13081 27421 13093 27455
rect 13127 27421 13139 27455
rect 13081 27415 13139 27421
rect 12268 27384 12296 27415
rect 12342 27384 12348 27396
rect 12268 27356 12348 27384
rect 12342 27344 12348 27356
rect 12400 27344 12406 27396
rect 13096 27384 13124 27415
rect 13262 27412 13268 27464
rect 13320 27452 13326 27464
rect 14090 27452 14096 27464
rect 13320 27424 13413 27452
rect 14051 27424 14096 27452
rect 13320 27412 13326 27424
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14642 27412 14648 27464
rect 14700 27452 14706 27464
rect 14829 27455 14887 27461
rect 14829 27452 14841 27455
rect 14700 27424 14841 27452
rect 14700 27412 14706 27424
rect 14829 27421 14841 27424
rect 14875 27421 14887 27455
rect 14829 27415 14887 27421
rect 16942 27412 16948 27464
rect 17000 27452 17006 27464
rect 17129 27455 17187 27461
rect 17129 27452 17141 27455
rect 17000 27424 17141 27452
rect 17000 27412 17006 27424
rect 17129 27421 17141 27424
rect 17175 27421 17187 27455
rect 17129 27415 17187 27421
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 18187 27424 19257 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 19245 27421 19257 27424
rect 19291 27452 19303 27455
rect 19426 27452 19432 27464
rect 19291 27424 19432 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 20456 27461 20484 27492
rect 20622 27480 20628 27492
rect 20680 27480 20686 27532
rect 22005 27523 22063 27529
rect 22005 27489 22017 27523
rect 22051 27520 22063 27523
rect 22278 27520 22284 27532
rect 22051 27492 22284 27520
rect 22051 27489 22063 27492
rect 22005 27483 22063 27489
rect 22278 27480 22284 27492
rect 22336 27480 22342 27532
rect 28000 27529 28028 27628
rect 29914 27616 29920 27628
rect 29972 27616 29978 27668
rect 31018 27616 31024 27668
rect 31076 27656 31082 27668
rect 31278 27659 31336 27665
rect 31278 27656 31290 27659
rect 31076 27628 31290 27656
rect 31076 27616 31082 27628
rect 31278 27625 31290 27628
rect 31324 27625 31336 27659
rect 31278 27619 31336 27625
rect 30926 27588 30932 27600
rect 28736 27560 30932 27588
rect 27985 27523 28043 27529
rect 27985 27489 27997 27523
rect 28031 27489 28043 27523
rect 27985 27483 28043 27489
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21082 27452 21088 27464
rect 20855 27424 21088 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21082 27412 21088 27424
rect 21140 27452 21146 27464
rect 21784 27455 21842 27461
rect 21784 27452 21796 27455
rect 21140 27424 21796 27452
rect 21140 27412 21146 27424
rect 21784 27421 21796 27424
rect 21830 27452 21842 27455
rect 22186 27452 22192 27464
rect 21830 27424 22192 27452
rect 21830 27421 21842 27424
rect 21784 27415 21842 27421
rect 22186 27412 22192 27424
rect 22244 27452 22250 27464
rect 22646 27452 22652 27464
rect 22244 27424 22652 27452
rect 22244 27412 22250 27424
rect 22646 27412 22652 27424
rect 22704 27412 22710 27464
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 25501 27455 25559 27461
rect 25501 27452 25513 27455
rect 23348 27424 25513 27452
rect 23348 27412 23354 27424
rect 25501 27421 25513 27424
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 27709 27455 27767 27461
rect 27709 27421 27721 27455
rect 27755 27421 27767 27455
rect 27709 27415 27767 27421
rect 13354 27384 13360 27396
rect 13096 27356 13360 27384
rect 13354 27344 13360 27356
rect 13412 27344 13418 27396
rect 15010 27384 15016 27396
rect 14971 27356 15016 27384
rect 15010 27344 15016 27356
rect 15068 27344 15074 27396
rect 20530 27344 20536 27396
rect 20588 27384 20594 27396
rect 20625 27387 20683 27393
rect 20625 27384 20637 27387
rect 20588 27356 20637 27384
rect 20588 27344 20594 27356
rect 20625 27353 20637 27356
rect 20671 27353 20683 27387
rect 20625 27347 20683 27353
rect 21637 27387 21695 27393
rect 21637 27353 21649 27387
rect 21683 27384 21695 27387
rect 22002 27384 22008 27396
rect 21683 27356 22008 27384
rect 21683 27353 21695 27356
rect 21637 27347 21695 27353
rect 22002 27344 22008 27356
rect 22060 27344 22066 27396
rect 26326 27344 26332 27396
rect 26384 27344 26390 27396
rect 27724 27384 27752 27415
rect 27798 27412 27804 27464
rect 27856 27452 27862 27464
rect 28626 27452 28632 27464
rect 27856 27424 27901 27452
rect 28587 27424 28632 27452
rect 27856 27412 27862 27424
rect 28626 27412 28632 27424
rect 28684 27412 28690 27464
rect 27890 27384 27896 27396
rect 27724 27356 27896 27384
rect 27890 27344 27896 27356
rect 27948 27344 27954 27396
rect 7558 27276 7564 27328
rect 7616 27316 7622 27328
rect 8202 27316 8208 27328
rect 7616 27288 8208 27316
rect 7616 27276 7622 27288
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 21174 27276 21180 27328
rect 21232 27316 21238 27328
rect 22281 27319 22339 27325
rect 22281 27316 22293 27319
rect 21232 27288 22293 27316
rect 21232 27276 21238 27288
rect 22281 27285 22293 27288
rect 22327 27285 22339 27319
rect 22281 27279 22339 27285
rect 26510 27276 26516 27328
rect 26568 27316 26574 27328
rect 28736 27316 28764 27560
rect 30926 27548 30932 27560
rect 30984 27548 30990 27600
rect 47026 27588 47032 27600
rect 46308 27560 47032 27588
rect 29730 27480 29736 27532
rect 29788 27520 29794 27532
rect 29825 27523 29883 27529
rect 29825 27520 29837 27523
rect 29788 27492 29837 27520
rect 29788 27480 29794 27492
rect 29825 27489 29837 27492
rect 29871 27489 29883 27523
rect 30944 27520 30972 27548
rect 31386 27520 31392 27532
rect 30944 27492 31392 27520
rect 29825 27483 29883 27489
rect 31386 27480 31392 27492
rect 31444 27480 31450 27532
rect 46308 27529 46336 27560
rect 47026 27548 47032 27560
rect 47084 27548 47090 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46474 27520 46480 27532
rect 46435 27492 46480 27520
rect 46293 27483 46351 27489
rect 46474 27480 46480 27492
rect 46532 27480 46538 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 28997 27455 29055 27461
rect 28997 27421 29009 27455
rect 29043 27452 29055 27455
rect 29549 27455 29607 27461
rect 29549 27452 29561 27455
rect 29043 27424 29561 27452
rect 29043 27421 29055 27424
rect 28997 27415 29055 27421
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 28813 27387 28871 27393
rect 28813 27353 28825 27387
rect 28859 27384 28871 27387
rect 28902 27384 28908 27396
rect 28859 27356 28908 27384
rect 28859 27353 28871 27356
rect 28813 27347 28871 27353
rect 28902 27344 28908 27356
rect 28960 27384 28966 27396
rect 29454 27384 29460 27396
rect 28960 27356 29460 27384
rect 28960 27344 28966 27356
rect 29454 27344 29460 27356
rect 29512 27344 29518 27396
rect 29564 27384 29592 27415
rect 30190 27412 30196 27464
rect 30248 27452 30254 27464
rect 31021 27455 31079 27461
rect 31021 27452 31033 27455
rect 30248 27424 31033 27452
rect 30248 27412 30254 27424
rect 31021 27421 31033 27424
rect 31067 27421 31079 27455
rect 31021 27415 31079 27421
rect 30558 27384 30564 27396
rect 29564 27356 30564 27384
rect 30558 27344 30564 27356
rect 30616 27344 30622 27396
rect 32306 27344 32312 27396
rect 32364 27344 32370 27396
rect 26568 27288 28764 27316
rect 26568 27276 26574 27288
rect 28994 27276 29000 27328
rect 29052 27316 29058 27328
rect 30101 27319 30159 27325
rect 30101 27316 30113 27319
rect 29052 27288 30113 27316
rect 29052 27276 29058 27288
rect 30101 27285 30113 27288
rect 30147 27285 30159 27319
rect 30101 27279 30159 27285
rect 30374 27276 30380 27328
rect 30432 27316 30438 27328
rect 32214 27316 32220 27328
rect 30432 27288 32220 27316
rect 30432 27276 30438 27288
rect 32214 27276 32220 27288
rect 32272 27316 32278 27328
rect 32769 27319 32827 27325
rect 32769 27316 32781 27319
rect 32272 27288 32781 27316
rect 32272 27276 32278 27288
rect 32769 27285 32781 27288
rect 32815 27285 32827 27319
rect 32769 27279 32827 27285
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 15010 27112 15016 27124
rect 14971 27084 15016 27112
rect 15010 27072 15016 27084
rect 15068 27072 15074 27124
rect 22278 27112 22284 27124
rect 21284 27084 22284 27112
rect 12894 27004 12900 27056
rect 12952 27044 12958 27056
rect 21174 27044 21180 27056
rect 12952 27016 21180 27044
rect 12952 27004 12958 27016
rect 21174 27004 21180 27016
rect 21232 27004 21238 27056
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26976 10379 26979
rect 11146 26976 11152 26988
rect 10367 26948 11152 26976
rect 10367 26945 10379 26948
rect 10321 26939 10379 26945
rect 11146 26936 11152 26948
rect 11204 26936 11210 26988
rect 12526 26976 12532 26988
rect 12487 26948 12532 26976
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 12713 26979 12771 26985
rect 12713 26945 12725 26979
rect 12759 26976 12771 26979
rect 13814 26976 13820 26988
rect 12759 26948 13820 26976
rect 12759 26945 12771 26948
rect 12713 26939 12771 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26976 14979 26979
rect 15010 26976 15016 26988
rect 14967 26948 15016 26976
rect 14967 26945 14979 26948
rect 14921 26939 14979 26945
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20496 26948 20821 26976
rect 20496 26936 20502 26948
rect 20809 26945 20821 26948
rect 20855 26945 20867 26979
rect 20809 26939 20867 26945
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26976 21051 26979
rect 21082 26976 21088 26988
rect 21039 26948 21088 26976
rect 21039 26945 21051 26948
rect 20993 26939 21051 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 21284 26985 21312 27084
rect 22278 27072 22284 27084
rect 22336 27112 22342 27124
rect 22462 27112 22468 27124
rect 22336 27084 22468 27112
rect 22336 27072 22342 27084
rect 22462 27072 22468 27084
rect 22520 27072 22526 27124
rect 23934 27112 23940 27124
rect 23400 27084 23940 27112
rect 22005 27047 22063 27053
rect 22005 27013 22017 27047
rect 22051 27044 22063 27047
rect 23400 27044 23428 27084
rect 23934 27072 23940 27084
rect 23992 27072 23998 27124
rect 26237 27115 26295 27121
rect 26237 27081 26249 27115
rect 26283 27112 26295 27115
rect 26510 27112 26516 27124
rect 26283 27084 26516 27112
rect 26283 27081 26295 27084
rect 26237 27075 26295 27081
rect 26510 27072 26516 27084
rect 26568 27072 26574 27124
rect 28994 27072 29000 27124
rect 29052 27072 29058 27124
rect 30006 27072 30012 27124
rect 30064 27112 30070 27124
rect 46842 27112 46848 27124
rect 30064 27084 46848 27112
rect 30064 27072 30070 27084
rect 46842 27072 46848 27084
rect 46900 27072 46906 27124
rect 22051 27016 23428 27044
rect 23477 27047 23535 27053
rect 22051 27013 22063 27016
rect 22005 27007 22063 27013
rect 23477 27013 23489 27047
rect 23523 27044 23535 27047
rect 23566 27044 23572 27056
rect 23523 27016 23572 27044
rect 23523 27013 23535 27016
rect 23477 27007 23535 27013
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 24949 27047 25007 27053
rect 24949 27044 24961 27047
rect 24504 27016 24961 27044
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 21818 26936 21824 26988
rect 21876 26976 21882 26988
rect 21913 26979 21971 26985
rect 21913 26976 21925 26979
rect 21876 26948 21925 26976
rect 21876 26936 21882 26948
rect 21913 26945 21925 26948
rect 21959 26945 21971 26979
rect 21913 26939 21971 26945
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26976 22247 26979
rect 22278 26976 22284 26988
rect 22235 26948 22284 26976
rect 22235 26945 22247 26948
rect 22189 26939 22247 26945
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 22462 26976 22468 26988
rect 22423 26948 22468 26976
rect 22462 26936 22468 26948
rect 22520 26936 22526 26988
rect 23014 26936 23020 26988
rect 23072 26976 23078 26988
rect 23293 26979 23351 26985
rect 23293 26976 23305 26979
rect 23072 26948 23305 26976
rect 23072 26936 23078 26948
rect 23293 26945 23305 26948
rect 23339 26976 23351 26979
rect 24504 26976 24532 27016
rect 24949 27013 24961 27016
rect 24995 27044 25007 27047
rect 26970 27044 26976 27056
rect 24995 27016 26976 27044
rect 24995 27013 25007 27016
rect 24949 27007 25007 27013
rect 26970 27004 26976 27016
rect 27028 27004 27034 27056
rect 29012 27044 29040 27072
rect 28644 27016 29040 27044
rect 29365 27047 29423 27053
rect 24762 26976 24768 26988
rect 23339 26948 24532 26976
rect 24723 26948 24768 26976
rect 23339 26945 23351 26948
rect 23293 26939 23351 26945
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 26050 26976 26056 26988
rect 26011 26948 26056 26976
rect 26050 26936 26056 26948
rect 26108 26936 26114 26988
rect 28644 26985 28672 27016
rect 29365 27013 29377 27047
rect 29411 27044 29423 27047
rect 30101 27047 30159 27053
rect 30101 27044 30113 27047
rect 29411 27016 30113 27044
rect 29411 27013 29423 27016
rect 29365 27007 29423 27013
rect 30101 27013 30113 27016
rect 30147 27013 30159 27047
rect 30101 27007 30159 27013
rect 31110 27004 31116 27056
rect 31168 27004 31174 27056
rect 32217 27047 32275 27053
rect 32217 27013 32229 27047
rect 32263 27044 32275 27047
rect 32306 27044 32312 27056
rect 32263 27016 32312 27044
rect 32263 27013 32275 27016
rect 32217 27007 32275 27013
rect 32306 27004 32312 27016
rect 32364 27004 32370 27056
rect 28629 26979 28687 26985
rect 28629 26945 28641 26979
rect 28675 26945 28687 26979
rect 28629 26939 28687 26945
rect 28817 26977 28875 26983
rect 28817 26943 28829 26977
rect 28863 26943 28875 26977
rect 28817 26937 28875 26943
rect 28905 26979 28963 26985
rect 28905 26945 28917 26979
rect 28951 26945 28963 26979
rect 28905 26939 28963 26945
rect 29043 26979 29101 26985
rect 29043 26945 29055 26979
rect 29089 26945 29101 26979
rect 29043 26939 29101 26945
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26877 7895 26911
rect 7837 26871 7895 26877
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 8110 26908 8116 26920
rect 8067 26880 8116 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 7852 26840 7880 26871
rect 8110 26868 8116 26880
rect 8168 26868 8174 26920
rect 8202 26868 8208 26920
rect 8260 26908 8266 26920
rect 8297 26911 8355 26917
rect 8297 26908 8309 26911
rect 8260 26880 8309 26908
rect 8260 26868 8266 26880
rect 8297 26877 8309 26880
rect 8343 26877 8355 26911
rect 10413 26911 10471 26917
rect 10413 26908 10425 26911
rect 8297 26871 8355 26877
rect 10336 26880 10425 26908
rect 10336 26852 10364 26880
rect 10413 26877 10425 26880
rect 10459 26877 10471 26911
rect 10413 26871 10471 26877
rect 20901 26911 20959 26917
rect 20901 26877 20913 26911
rect 20947 26908 20959 26911
rect 22002 26908 22008 26920
rect 20947 26880 22008 26908
rect 20947 26877 20959 26880
rect 20901 26871 20959 26877
rect 22002 26868 22008 26880
rect 22060 26908 22066 26920
rect 22097 26911 22155 26917
rect 22097 26908 22109 26911
rect 22060 26880 22109 26908
rect 22060 26868 22066 26880
rect 22097 26877 22109 26880
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 23106 26868 23112 26920
rect 23164 26908 23170 26920
rect 26068 26908 26096 26936
rect 23164 26880 26096 26908
rect 23164 26868 23170 26880
rect 28828 26852 28856 26937
rect 9306 26840 9312 26852
rect 7852 26812 9312 26840
rect 9306 26800 9312 26812
rect 9364 26800 9370 26852
rect 10318 26800 10324 26852
rect 10376 26800 10382 26852
rect 28810 26800 28816 26852
rect 28868 26800 28874 26852
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 10689 26775 10747 26781
rect 10689 26772 10701 26775
rect 9732 26744 10701 26772
rect 9732 26732 9738 26744
rect 10689 26741 10701 26744
rect 10735 26741 10747 26775
rect 10689 26735 10747 26741
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 12492 26744 12541 26772
rect 12492 26732 12498 26744
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 12529 26735 12587 26741
rect 12618 26732 12624 26784
rect 12676 26772 12682 26784
rect 15010 26772 15016 26784
rect 12676 26744 15016 26772
rect 12676 26732 12682 26744
rect 15010 26732 15016 26744
rect 15068 26732 15074 26784
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 20533 26775 20591 26781
rect 20533 26772 20545 26775
rect 18012 26744 20545 26772
rect 18012 26732 18018 26744
rect 20533 26741 20545 26744
rect 20579 26741 20591 26775
rect 20533 26735 20591 26741
rect 21085 26775 21143 26781
rect 21085 26741 21097 26775
rect 21131 26772 21143 26775
rect 21910 26772 21916 26784
rect 21131 26744 21916 26772
rect 21131 26741 21143 26744
rect 21085 26735 21143 26741
rect 21910 26732 21916 26744
rect 21968 26772 21974 26784
rect 22299 26775 22357 26781
rect 22299 26772 22311 26775
rect 21968 26744 22311 26772
rect 21968 26732 21974 26744
rect 22299 26741 22311 26744
rect 22345 26741 22357 26775
rect 28929 26772 28957 26939
rect 29058 26852 29086 26939
rect 29178 26936 29184 26988
rect 29236 26976 29242 26988
rect 29236 26948 29281 26976
rect 29236 26936 29242 26948
rect 31386 26936 31392 26988
rect 31444 26976 31450 26988
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 31444 26948 32137 26976
rect 31444 26936 31450 26948
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 29822 26908 29828 26920
rect 29735 26880 29828 26908
rect 29822 26868 29828 26880
rect 29880 26908 29886 26920
rect 30190 26908 30196 26920
rect 29880 26880 30196 26908
rect 29880 26868 29886 26880
rect 30190 26868 30196 26880
rect 30248 26868 30254 26920
rect 29058 26812 29092 26852
rect 29086 26800 29092 26812
rect 29144 26800 29150 26852
rect 29178 26800 29184 26852
rect 29236 26840 29242 26852
rect 29840 26840 29868 26868
rect 29236 26812 29868 26840
rect 29236 26800 29242 26812
rect 29454 26772 29460 26784
rect 28929 26744 29460 26772
rect 22299 26735 22357 26741
rect 29454 26732 29460 26744
rect 29512 26772 29518 26784
rect 31573 26775 31631 26781
rect 31573 26772 31585 26775
rect 29512 26744 31585 26772
rect 29512 26732 29518 26744
rect 31573 26741 31585 26744
rect 31619 26741 31631 26775
rect 31573 26735 31631 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 8110 26568 8116 26580
rect 8071 26540 8116 26568
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 12526 26568 12532 26580
rect 12487 26540 12532 26568
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 19426 26568 19432 26580
rect 19387 26540 19432 26568
rect 19426 26528 19432 26540
rect 19484 26528 19490 26580
rect 22002 26568 22008 26580
rect 21963 26540 22008 26568
rect 22002 26528 22008 26540
rect 22060 26528 22066 26580
rect 23106 26568 23112 26580
rect 22480 26540 23112 26568
rect 13262 26500 13268 26512
rect 12268 26472 13268 26500
rect 9674 26432 9680 26444
rect 9635 26404 9680 26432
rect 9674 26392 9680 26404
rect 9732 26392 9738 26444
rect 11146 26432 11152 26444
rect 11059 26404 11152 26432
rect 11146 26392 11152 26404
rect 11204 26432 11210 26444
rect 12268 26432 12296 26472
rect 13262 26460 13268 26472
rect 13320 26460 13326 26512
rect 14274 26500 14280 26512
rect 14235 26472 14280 26500
rect 14274 26460 14280 26472
rect 14332 26460 14338 26512
rect 20622 26460 20628 26512
rect 20680 26500 20686 26512
rect 22480 26500 22508 26540
rect 23106 26528 23112 26540
rect 23164 26528 23170 26580
rect 23198 26528 23204 26580
rect 23256 26568 23262 26580
rect 31110 26568 31116 26580
rect 23256 26540 26648 26568
rect 31071 26540 31116 26568
rect 23256 26528 23262 26540
rect 26510 26500 26516 26512
rect 20680 26472 22508 26500
rect 22572 26472 23612 26500
rect 26471 26472 26516 26500
rect 20680 26460 20686 26472
rect 22572 26444 22600 26472
rect 11204 26404 12296 26432
rect 11204 26392 11210 26404
rect 7377 26367 7435 26373
rect 7377 26333 7389 26367
rect 7423 26364 7435 26367
rect 8018 26364 8024 26376
rect 7423 26336 8024 26364
rect 7423 26333 7435 26336
rect 7377 26327 7435 26333
rect 8018 26324 8024 26336
rect 8076 26324 8082 26376
rect 9398 26364 9404 26376
rect 9359 26336 9404 26364
rect 9398 26324 9404 26336
rect 9456 26324 9462 26376
rect 12158 26364 12164 26376
rect 12119 26336 12164 26364
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12268 26373 12296 26404
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12989 26435 13047 26441
rect 12989 26432 13001 26435
rect 12400 26404 12445 26432
rect 12544 26404 13001 26432
rect 12400 26392 12406 26404
rect 12544 26373 12572 26404
rect 12989 26401 13001 26404
rect 13035 26432 13047 26435
rect 13446 26432 13452 26444
rect 13035 26404 13452 26432
rect 13035 26401 13047 26404
rect 12989 26395 13047 26401
rect 13446 26392 13452 26404
rect 13504 26392 13510 26444
rect 21818 26392 21824 26444
rect 21876 26432 21882 26444
rect 22278 26432 22284 26444
rect 21876 26404 22284 26432
rect 21876 26392 21882 26404
rect 22278 26392 22284 26404
rect 22336 26432 22342 26444
rect 22554 26432 22560 26444
rect 22336 26404 22560 26432
rect 22336 26392 22342 26404
rect 22554 26392 22560 26404
rect 22612 26392 22618 26444
rect 23106 26432 23112 26444
rect 22940 26404 23112 26432
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 13262 26324 13268 26376
rect 13320 26324 13326 26376
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13541 26367 13599 26373
rect 13412 26336 13457 26364
rect 13412 26324 13418 26336
rect 13541 26333 13553 26367
rect 13587 26364 13599 26367
rect 13814 26364 13820 26376
rect 13587 26336 13820 26364
rect 13587 26333 13599 26336
rect 13541 26327 13599 26333
rect 13814 26324 13820 26336
rect 13872 26364 13878 26376
rect 14458 26364 14464 26376
rect 13872 26336 14464 26364
rect 13872 26324 13878 26336
rect 14458 26324 14464 26336
rect 14516 26324 14522 26376
rect 14642 26364 14648 26376
rect 14603 26336 14648 26364
rect 14642 26324 14648 26336
rect 14700 26324 14706 26376
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 20254 26364 20260 26376
rect 19291 26336 20260 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 20254 26324 20260 26336
rect 20312 26364 20318 26376
rect 20530 26364 20536 26376
rect 20312 26336 20536 26364
rect 20312 26324 20318 26336
rect 20530 26324 20536 26336
rect 20588 26324 20594 26376
rect 21637 26367 21695 26373
rect 21637 26333 21649 26367
rect 21683 26364 21695 26367
rect 22002 26364 22008 26376
rect 21683 26336 22008 26364
rect 21683 26333 21695 26336
rect 21637 26327 21695 26333
rect 22002 26324 22008 26336
rect 22060 26324 22066 26376
rect 22646 26364 22652 26376
rect 22607 26336 22652 26364
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 22940 26373 22968 26404
rect 23106 26392 23112 26404
rect 23164 26432 23170 26444
rect 23477 26435 23535 26441
rect 23477 26432 23489 26435
rect 23164 26404 23489 26432
rect 23164 26392 23170 26404
rect 23477 26401 23489 26404
rect 23523 26401 23535 26435
rect 23477 26395 23535 26401
rect 23584 26373 23612 26472
rect 26510 26460 26516 26472
rect 26568 26460 26574 26512
rect 26620 26500 26648 26540
rect 31110 26528 31116 26540
rect 31168 26528 31174 26580
rect 26620 26472 31754 26500
rect 27706 26432 27712 26444
rect 26712 26404 27712 26432
rect 22925 26367 22983 26373
rect 22925 26333 22937 26367
rect 22971 26333 22983 26367
rect 22925 26327 22983 26333
rect 23385 26367 23443 26373
rect 23385 26333 23397 26367
rect 23431 26333 23443 26367
rect 23385 26327 23443 26333
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 10410 26256 10416 26308
rect 10468 26256 10474 26308
rect 13170 26296 13176 26308
rect 13131 26268 13176 26296
rect 13170 26256 13176 26268
rect 13228 26256 13234 26308
rect 7466 26228 7472 26240
rect 7427 26200 7472 26228
rect 7466 26188 7472 26200
rect 7524 26188 7530 26240
rect 13280 26237 13308 26324
rect 14366 26256 14372 26308
rect 14424 26296 14430 26308
rect 14829 26299 14887 26305
rect 14829 26296 14841 26299
rect 14424 26268 14841 26296
rect 14424 26256 14430 26268
rect 14829 26265 14841 26268
rect 14875 26265 14887 26299
rect 14829 26259 14887 26265
rect 21542 26256 21548 26308
rect 21600 26296 21606 26308
rect 21821 26299 21879 26305
rect 21821 26296 21833 26299
rect 21600 26268 21833 26296
rect 21600 26256 21606 26268
rect 21821 26265 21833 26268
rect 21867 26265 21879 26299
rect 21821 26259 21879 26265
rect 22465 26299 22523 26305
rect 22465 26265 22477 26299
rect 22511 26296 22523 26299
rect 22554 26296 22560 26308
rect 22511 26268 22560 26296
rect 22511 26265 22523 26268
rect 22465 26259 22523 26265
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 22738 26256 22744 26308
rect 22796 26296 22802 26308
rect 23400 26296 23428 26327
rect 23750 26324 23756 26376
rect 23808 26364 23814 26376
rect 26712 26373 26740 26404
rect 27706 26392 27712 26404
rect 27764 26392 27770 26444
rect 31726 26432 31754 26472
rect 46842 26432 46848 26444
rect 31726 26404 46848 26432
rect 46842 26392 46848 26404
rect 46900 26392 46906 26444
rect 26513 26367 26571 26373
rect 26513 26364 26525 26367
rect 23808 26336 26525 26364
rect 23808 26324 23814 26336
rect 26513 26333 26525 26336
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26333 26755 26367
rect 26697 26327 26755 26333
rect 26789 26367 26847 26373
rect 26789 26333 26801 26367
rect 26835 26333 26847 26367
rect 27246 26364 27252 26376
rect 27207 26336 27252 26364
rect 26789 26327 26847 26333
rect 22796 26268 23428 26296
rect 26804 26296 26832 26327
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 27433 26367 27491 26373
rect 27433 26333 27445 26367
rect 27479 26333 27491 26367
rect 27433 26327 27491 26333
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 26804 26268 27353 26296
rect 22796 26256 22802 26268
rect 27341 26265 27353 26268
rect 27387 26265 27399 26299
rect 27341 26259 27399 26265
rect 13265 26231 13323 26237
rect 13265 26197 13277 26231
rect 13311 26197 13323 26231
rect 13265 26191 13323 26197
rect 13446 26188 13452 26240
rect 13504 26228 13510 26240
rect 14461 26231 14519 26237
rect 14461 26228 14473 26231
rect 13504 26200 14473 26228
rect 13504 26188 13510 26200
rect 14461 26197 14473 26200
rect 14507 26197 14519 26231
rect 14461 26191 14519 26197
rect 14550 26188 14556 26240
rect 14608 26228 14614 26240
rect 14608 26200 14653 26228
rect 14608 26188 14614 26200
rect 22002 26188 22008 26240
rect 22060 26228 22066 26240
rect 22833 26231 22891 26237
rect 22833 26228 22845 26231
rect 22060 26200 22845 26228
rect 22060 26188 22066 26200
rect 22833 26197 22845 26200
rect 22879 26228 22891 26231
rect 23014 26228 23020 26240
rect 22879 26200 23020 26228
rect 22879 26197 22891 26200
rect 22833 26191 22891 26197
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 27448 26228 27476 26327
rect 30558 26324 30564 26376
rect 30616 26364 30622 26376
rect 31021 26367 31079 26373
rect 31021 26364 31033 26367
rect 30616 26336 31033 26364
rect 30616 26324 30622 26336
rect 31021 26333 31033 26336
rect 31067 26364 31079 26367
rect 31386 26364 31392 26376
rect 31067 26336 31392 26364
rect 31067 26333 31079 26336
rect 31021 26327 31079 26333
rect 31386 26324 31392 26336
rect 31444 26324 31450 26376
rect 26844 26200 27476 26228
rect 26844 26188 26850 26200
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10505 26027 10563 26033
rect 10505 26024 10517 26027
rect 10468 25996 10517 26024
rect 10468 25984 10474 25996
rect 10505 25993 10517 25996
rect 10551 25993 10563 26027
rect 10505 25987 10563 25993
rect 14274 25984 14280 26036
rect 14332 26024 14338 26036
rect 15657 26027 15715 26033
rect 15657 26024 15669 26027
rect 14332 25996 15669 26024
rect 14332 25984 14338 25996
rect 15657 25993 15669 25996
rect 15703 25993 15715 26027
rect 15657 25987 15715 25993
rect 23566 25984 23572 26036
rect 23624 26024 23630 26036
rect 24213 26027 24271 26033
rect 24213 26024 24225 26027
rect 23624 25996 24225 26024
rect 23624 25984 23630 25996
rect 24213 25993 24225 25996
rect 24259 25993 24271 26027
rect 27525 26027 27583 26033
rect 27525 26024 27537 26027
rect 24213 25987 24271 25993
rect 26068 25996 27537 26024
rect 7466 25916 7472 25968
rect 7524 25956 7530 25968
rect 8205 25959 8263 25965
rect 8205 25956 8217 25959
rect 7524 25928 8217 25956
rect 7524 25916 7530 25928
rect 8205 25925 8217 25928
rect 8251 25925 8263 25959
rect 8205 25919 8263 25925
rect 20254 25916 20260 25968
rect 20312 25916 20318 25968
rect 26068 25965 26096 25996
rect 27525 25993 27537 25996
rect 27571 25993 27583 26027
rect 27525 25987 27583 25993
rect 22741 25959 22799 25965
rect 22741 25925 22753 25959
rect 22787 25956 22799 25959
rect 26053 25959 26111 25965
rect 22787 25928 24072 25956
rect 22787 25925 22799 25928
rect 22741 25919 22799 25925
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 10413 25891 10471 25897
rect 10413 25888 10425 25891
rect 9916 25860 10425 25888
rect 9916 25848 9922 25860
rect 10413 25857 10425 25860
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 13078 25848 13084 25900
rect 13136 25848 13142 25900
rect 15286 25848 15292 25900
rect 15344 25848 15350 25900
rect 16114 25848 16120 25900
rect 16172 25888 16178 25900
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 16172 25860 17141 25888
rect 16172 25848 16178 25860
rect 17129 25857 17141 25860
rect 17175 25857 17187 25891
rect 17129 25851 17187 25857
rect 17313 25891 17371 25897
rect 17313 25857 17325 25891
rect 17359 25888 17371 25891
rect 17954 25888 17960 25900
rect 17359 25860 17960 25888
rect 17359 25857 17371 25860
rect 17313 25851 17371 25857
rect 17954 25848 17960 25860
rect 18012 25848 18018 25900
rect 23014 25888 23020 25900
rect 22975 25860 23020 25888
rect 23014 25848 23020 25860
rect 23072 25848 23078 25900
rect 23106 25891 23164 25897
rect 23106 25857 23118 25891
rect 23152 25857 23164 25891
rect 23106 25851 23164 25857
rect 23206 25891 23264 25897
rect 23206 25857 23218 25891
rect 23252 25857 23264 25891
rect 23382 25888 23388 25900
rect 23343 25860 23388 25888
rect 23206 25851 23264 25857
rect 8021 25823 8079 25829
rect 8021 25789 8033 25823
rect 8067 25820 8079 25823
rect 8294 25820 8300 25832
rect 8067 25792 8300 25820
rect 8067 25789 8079 25792
rect 8021 25783 8079 25789
rect 8294 25780 8300 25792
rect 8352 25780 8358 25832
rect 8481 25823 8539 25829
rect 8481 25789 8493 25823
rect 8527 25789 8539 25823
rect 8481 25783 8539 25789
rect 3510 25712 3516 25764
rect 3568 25752 3574 25764
rect 8496 25752 8524 25783
rect 11606 25780 11612 25832
rect 11664 25820 11670 25832
rect 11701 25823 11759 25829
rect 11701 25820 11713 25823
rect 11664 25792 11713 25820
rect 11664 25780 11670 25792
rect 11701 25789 11713 25792
rect 11747 25789 11759 25823
rect 11701 25783 11759 25789
rect 11977 25823 12035 25829
rect 11977 25789 11989 25823
rect 12023 25820 12035 25823
rect 12434 25820 12440 25832
rect 12023 25792 12440 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 12434 25780 12440 25792
rect 12492 25780 12498 25832
rect 13906 25820 13912 25832
rect 13867 25792 13912 25820
rect 13906 25780 13912 25792
rect 13964 25780 13970 25832
rect 14182 25820 14188 25832
rect 14143 25792 14188 25820
rect 14182 25780 14188 25792
rect 14240 25780 14246 25832
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19521 25823 19579 25829
rect 19521 25820 19533 25823
rect 19484 25792 19533 25820
rect 19484 25780 19490 25792
rect 19521 25789 19533 25792
rect 19567 25789 19579 25823
rect 19521 25783 19579 25789
rect 19797 25823 19855 25829
rect 19797 25789 19809 25823
rect 19843 25820 19855 25823
rect 19843 25792 22094 25820
rect 19843 25789 19855 25792
rect 19797 25783 19855 25789
rect 3568 25724 8524 25752
rect 3568 25712 3574 25724
rect 13446 25684 13452 25696
rect 13407 25656 13452 25684
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 17126 25684 17132 25696
rect 17087 25656 17132 25684
rect 17126 25644 17132 25656
rect 17184 25644 17190 25696
rect 21269 25687 21327 25693
rect 21269 25653 21281 25687
rect 21315 25684 21327 25687
rect 21542 25684 21548 25696
rect 21315 25656 21548 25684
rect 21315 25653 21327 25656
rect 21269 25647 21327 25653
rect 21542 25644 21548 25656
rect 21600 25644 21606 25696
rect 22066 25684 22094 25792
rect 23121 25764 23149 25851
rect 23106 25712 23112 25764
rect 23164 25712 23170 25764
rect 23216 25752 23244 25851
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 24044 25897 24072 25928
rect 26053 25925 26065 25959
rect 26099 25925 26111 25959
rect 26053 25919 26111 25925
rect 26237 25959 26295 25965
rect 26237 25925 26249 25959
rect 26283 25956 26295 25959
rect 26510 25956 26516 25968
rect 26283 25928 26516 25956
rect 26283 25925 26295 25928
rect 26237 25919 26295 25925
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 27154 25956 27160 25968
rect 27115 25928 27160 25956
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 24029 25891 24087 25897
rect 24029 25857 24041 25891
rect 24075 25857 24087 25891
rect 24029 25851 24087 25857
rect 24305 25891 24363 25897
rect 24305 25857 24317 25891
rect 24351 25888 24363 25891
rect 24394 25888 24400 25900
rect 24351 25860 24400 25888
rect 24351 25857 24363 25860
rect 24305 25851 24363 25857
rect 24394 25848 24400 25860
rect 24452 25848 24458 25900
rect 26786 25848 26792 25900
rect 26844 25888 26850 25900
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26844 25860 26985 25888
rect 26844 25848 26850 25860
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 27264 25820 27292 25851
rect 27338 25848 27344 25900
rect 27396 25888 27402 25900
rect 28902 25888 28908 25900
rect 27396 25860 27441 25888
rect 28863 25860 28908 25888
rect 27396 25848 27402 25860
rect 28902 25848 28908 25860
rect 28960 25848 28966 25900
rect 28442 25820 28448 25832
rect 26988 25792 27292 25820
rect 27586 25792 28448 25820
rect 26988 25764 27016 25792
rect 23216 25724 26556 25752
rect 23845 25687 23903 25693
rect 23845 25684 23857 25687
rect 22066 25656 23857 25684
rect 23845 25653 23857 25656
rect 23891 25653 23903 25687
rect 23845 25647 23903 25653
rect 25774 25644 25780 25696
rect 25832 25684 25838 25696
rect 26421 25687 26479 25693
rect 26421 25684 26433 25687
rect 25832 25656 26433 25684
rect 25832 25644 25838 25656
rect 26421 25653 26433 25656
rect 26467 25653 26479 25687
rect 26528 25684 26556 25724
rect 26970 25712 26976 25764
rect 27028 25712 27034 25764
rect 27586 25684 27614 25792
rect 28442 25780 28448 25792
rect 28500 25820 28506 25832
rect 28994 25820 29000 25832
rect 28500 25792 29000 25820
rect 28500 25780 28506 25792
rect 28994 25780 29000 25792
rect 29052 25780 29058 25832
rect 26528 25656 27614 25684
rect 26421 25647 26479 25653
rect 28626 25644 28632 25696
rect 28684 25684 28690 25696
rect 28997 25687 29055 25693
rect 28997 25684 29009 25687
rect 28684 25656 29009 25684
rect 28684 25644 28690 25656
rect 28997 25653 29009 25656
rect 29043 25653 29055 25687
rect 28997 25647 29055 25653
rect 46290 25644 46296 25696
rect 46348 25684 46354 25696
rect 47765 25687 47823 25693
rect 47765 25684 47777 25687
rect 46348 25656 47777 25684
rect 46348 25644 46354 25656
rect 47765 25653 47777 25656
rect 47811 25653 47823 25687
rect 47765 25647 47823 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 9398 25440 9404 25492
rect 9456 25480 9462 25492
rect 9493 25483 9551 25489
rect 9493 25480 9505 25483
rect 9456 25452 9505 25480
rect 9456 25440 9462 25452
rect 9493 25449 9505 25452
rect 9539 25449 9551 25483
rect 11606 25480 11612 25492
rect 11567 25452 11612 25480
rect 9493 25443 9551 25449
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 13078 25440 13084 25492
rect 13136 25480 13142 25492
rect 13173 25483 13231 25489
rect 13173 25480 13185 25483
rect 13136 25452 13185 25480
rect 13136 25440 13142 25452
rect 13173 25449 13185 25452
rect 13219 25449 13231 25483
rect 13173 25443 13231 25449
rect 14093 25483 14151 25489
rect 14093 25449 14105 25483
rect 14139 25480 14151 25483
rect 14182 25480 14188 25492
rect 14139 25452 14188 25480
rect 14139 25449 14151 25452
rect 14093 25443 14151 25449
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 14458 25480 14464 25492
rect 14419 25452 14464 25480
rect 14458 25440 14464 25452
rect 14516 25440 14522 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15286 25480 15292 25492
rect 15151 25452 15292 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15286 25440 15292 25452
rect 15344 25440 15350 25492
rect 16114 25480 16120 25492
rect 16075 25452 16120 25480
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25480 20223 25483
rect 20254 25480 20260 25492
rect 20211 25452 20260 25480
rect 20211 25449 20223 25452
rect 20165 25443 20223 25449
rect 20254 25440 20260 25452
rect 20312 25440 20318 25492
rect 22646 25480 22652 25492
rect 22607 25452 22652 25480
rect 22646 25440 22652 25452
rect 22704 25440 22710 25492
rect 27614 25480 27620 25492
rect 27575 25452 27620 25480
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 27798 25440 27804 25492
rect 27856 25480 27862 25492
rect 27893 25483 27951 25489
rect 27893 25480 27905 25483
rect 27856 25452 27905 25480
rect 27856 25440 27862 25452
rect 27893 25449 27905 25452
rect 27939 25480 27951 25483
rect 28902 25480 28908 25492
rect 27939 25452 28908 25480
rect 27939 25449 27951 25452
rect 27893 25443 27951 25449
rect 28902 25440 28908 25452
rect 28960 25440 28966 25492
rect 14274 25372 14280 25424
rect 14332 25412 14338 25424
rect 14332 25384 14596 25412
rect 14332 25372 14338 25384
rect 14568 25353 14596 25384
rect 19150 25372 19156 25424
rect 19208 25412 19214 25424
rect 23198 25412 23204 25424
rect 19208 25384 23204 25412
rect 19208 25372 19214 25384
rect 23198 25372 23204 25384
rect 23256 25372 23262 25424
rect 28721 25415 28779 25421
rect 28721 25381 28733 25415
rect 28767 25412 28779 25415
rect 30282 25412 30288 25424
rect 28767 25384 30288 25412
rect 28767 25381 28779 25384
rect 28721 25375 28779 25381
rect 30282 25372 30288 25384
rect 30340 25372 30346 25424
rect 14553 25347 14611 25353
rect 9508 25316 11468 25344
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 9508 25285 9536 25316
rect 11440 25288 11468 25316
rect 14553 25313 14565 25347
rect 14599 25313 14611 25347
rect 17126 25344 17132 25356
rect 17087 25316 17132 25344
rect 14553 25307 14611 25313
rect 17126 25304 17132 25316
rect 17184 25304 17190 25356
rect 18138 25304 18144 25356
rect 18196 25344 18202 25356
rect 22002 25344 22008 25356
rect 18196 25316 19288 25344
rect 21963 25316 22008 25344
rect 18196 25304 18202 25316
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 8536 25248 9505 25276
rect 8536 25236 8542 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 10042 25276 10048 25288
rect 10003 25248 10048 25276
rect 9493 25239 9551 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25276 10287 25279
rect 10318 25276 10324 25288
rect 10275 25248 10324 25276
rect 10275 25245 10287 25248
rect 10229 25239 10287 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 11422 25236 11428 25288
rect 11480 25276 11486 25288
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 11480 25248 11621 25276
rect 11480 25236 11486 25248
rect 11609 25245 11621 25248
rect 11655 25276 11667 25279
rect 11882 25276 11888 25288
rect 11655 25248 11888 25276
rect 11655 25245 11667 25248
rect 11609 25239 11667 25245
rect 11882 25236 11888 25248
rect 11940 25236 11946 25288
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 1670 25208 1676 25220
rect 1631 25180 1676 25208
rect 1670 25168 1676 25180
rect 1728 25168 1734 25220
rect 13096 25208 13124 25239
rect 13998 25236 14004 25288
rect 14056 25276 14062 25288
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 14056 25248 14289 25276
rect 14056 25236 14062 25248
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 15013 25279 15071 25285
rect 15013 25276 15025 25279
rect 14277 25239 14335 25245
rect 14844 25248 15025 25276
rect 14844 25220 14872 25248
rect 15013 25245 15025 25248
rect 15059 25245 15071 25279
rect 15013 25239 15071 25245
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 16117 25279 16175 25285
rect 16117 25276 16129 25279
rect 15436 25248 16129 25276
rect 15436 25236 15442 25248
rect 16117 25245 16129 25248
rect 16163 25245 16175 25279
rect 16390 25276 16396 25288
rect 16351 25248 16396 25276
rect 16117 25239 16175 25245
rect 14090 25208 14096 25220
rect 13096 25180 14096 25208
rect 14090 25168 14096 25180
rect 14148 25208 14154 25220
rect 14826 25208 14832 25220
rect 14148 25180 14832 25208
rect 14148 25168 14154 25180
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 16132 25208 16160 25239
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 16850 25276 16856 25288
rect 16811 25248 16856 25276
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 19260 25285 19288 25316
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 22490 25347 22548 25353
rect 22490 25344 22502 25347
rect 22220 25316 22502 25344
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 19978 25276 19984 25288
rect 19576 25248 19984 25276
rect 19576 25236 19582 25248
rect 19978 25236 19984 25248
rect 20036 25276 20042 25288
rect 20073 25279 20131 25285
rect 20073 25276 20085 25279
rect 20036 25248 20085 25276
rect 20036 25236 20042 25248
rect 20073 25245 20085 25248
rect 20119 25276 20131 25279
rect 20717 25279 20775 25285
rect 20717 25276 20729 25279
rect 20119 25248 20729 25276
rect 20119 25245 20131 25248
rect 20073 25239 20131 25245
rect 20717 25245 20729 25248
rect 20763 25245 20775 25279
rect 20717 25239 20775 25245
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25245 21603 25279
rect 21545 25239 21603 25245
rect 18414 25208 18420 25220
rect 16132 25180 16436 25208
rect 18354 25180 18420 25208
rect 10134 25140 10140 25152
rect 10095 25112 10140 25140
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 13538 25100 13544 25152
rect 13596 25140 13602 25152
rect 15838 25140 15844 25152
rect 13596 25112 15844 25140
rect 13596 25100 13602 25112
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 16298 25140 16304 25152
rect 16259 25112 16304 25140
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 16408 25140 16436 25180
rect 18414 25168 18420 25180
rect 18472 25168 18478 25220
rect 21560 25208 21588 25239
rect 22094 25208 22100 25220
rect 21560 25180 22100 25208
rect 22094 25168 22100 25180
rect 22152 25168 22158 25220
rect 18601 25143 18659 25149
rect 18601 25140 18613 25143
rect 16408 25112 18613 25140
rect 18601 25109 18613 25112
rect 18647 25109 18659 25143
rect 19334 25140 19340 25152
rect 19295 25112 19340 25140
rect 18601 25103 18659 25109
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 20809 25143 20867 25149
rect 20809 25109 20821 25143
rect 20855 25140 20867 25143
rect 21082 25140 21088 25152
rect 20855 25112 21088 25140
rect 20855 25109 20867 25112
rect 20809 25103 20867 25109
rect 21082 25100 21088 25112
rect 21140 25100 21146 25152
rect 21358 25140 21364 25152
rect 21319 25112 21364 25140
rect 21358 25100 21364 25112
rect 21416 25100 21422 25152
rect 21542 25100 21548 25152
rect 21600 25140 21606 25152
rect 22220 25140 22248 25316
rect 22490 25313 22502 25316
rect 22536 25344 22548 25347
rect 23382 25344 23388 25356
rect 22536 25316 23388 25344
rect 22536 25313 22548 25316
rect 22490 25307 22548 25313
rect 23382 25304 23388 25316
rect 23440 25304 23446 25356
rect 27246 25344 27252 25356
rect 26620 25316 27252 25344
rect 22278 25236 22284 25288
rect 22336 25276 22342 25288
rect 25774 25276 25780 25288
rect 22336 25248 22381 25276
rect 25735 25248 25780 25276
rect 22336 25236 22342 25248
rect 25774 25236 25780 25248
rect 25832 25236 25838 25288
rect 26234 25236 26240 25288
rect 26292 25276 26298 25288
rect 26620 25285 26648 25316
rect 27246 25304 27252 25316
rect 27304 25304 27310 25356
rect 29270 25304 29276 25356
rect 29328 25344 29334 25356
rect 30009 25347 30067 25353
rect 29328 25316 29776 25344
rect 29328 25304 29334 25316
rect 26605 25279 26663 25285
rect 26605 25276 26617 25279
rect 26292 25248 26617 25276
rect 26292 25236 26298 25248
rect 26605 25245 26617 25248
rect 26651 25245 26663 25279
rect 27617 25279 27675 25285
rect 27617 25276 27629 25279
rect 26605 25239 26663 25245
rect 26804 25248 27629 25276
rect 26804 25220 26832 25248
rect 27617 25245 27629 25248
rect 27663 25245 27675 25279
rect 27617 25239 27675 25245
rect 27709 25279 27767 25285
rect 27709 25245 27721 25279
rect 27755 25276 27767 25279
rect 28442 25276 28448 25288
rect 27755 25248 28448 25276
rect 27755 25245 27767 25248
rect 27709 25239 27767 25245
rect 28442 25236 28448 25248
rect 28500 25236 28506 25288
rect 28626 25276 28632 25288
rect 28587 25248 28632 25276
rect 28626 25236 28632 25248
rect 28684 25236 28690 25288
rect 28718 25236 28724 25288
rect 28776 25276 28782 25288
rect 29748 25285 29776 25316
rect 30009 25313 30021 25347
rect 30055 25344 30067 25347
rect 40402 25344 40408 25356
rect 30055 25316 40408 25344
rect 30055 25313 30067 25316
rect 30009 25307 30067 25313
rect 40402 25304 40408 25316
rect 40460 25304 40466 25356
rect 46290 25344 46296 25356
rect 46251 25316 46296 25344
rect 46290 25304 46296 25316
rect 46348 25304 46354 25356
rect 28813 25279 28871 25285
rect 28813 25276 28825 25279
rect 28776 25248 28825 25276
rect 28776 25236 28782 25248
rect 28813 25245 28825 25248
rect 28859 25245 28871 25279
rect 28813 25239 28871 25245
rect 28905 25279 28963 25285
rect 28905 25245 28917 25279
rect 28951 25276 28963 25279
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 28951 25248 29561 25276
rect 28951 25245 28963 25248
rect 28905 25239 28963 25245
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 29822 25236 29828 25288
rect 29880 25276 29886 25288
rect 30098 25276 30104 25288
rect 29880 25248 29960 25276
rect 30059 25248 30104 25276
rect 29880 25236 29886 25248
rect 22373 25211 22431 25217
rect 22373 25177 22385 25211
rect 22419 25208 22431 25211
rect 22738 25208 22744 25220
rect 22419 25180 22744 25208
rect 22419 25177 22431 25180
rect 22373 25171 22431 25177
rect 22738 25168 22744 25180
rect 22796 25168 22802 25220
rect 26786 25208 26792 25220
rect 26747 25180 26792 25208
rect 26786 25168 26792 25180
rect 26844 25168 26850 25220
rect 27246 25168 27252 25220
rect 27304 25208 27310 25220
rect 27433 25211 27491 25217
rect 27433 25208 27445 25211
rect 27304 25180 27445 25208
rect 27304 25168 27310 25180
rect 27433 25177 27445 25180
rect 27479 25177 27491 25211
rect 28460 25208 28488 25236
rect 29932 25208 29960 25248
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 30558 25276 30564 25288
rect 30519 25248 30564 25276
rect 30558 25236 30564 25248
rect 30616 25236 30622 25288
rect 48130 25276 48136 25288
rect 48091 25248 48136 25276
rect 48130 25236 48136 25248
rect 48188 25236 48194 25288
rect 28460 25180 29960 25208
rect 46477 25211 46535 25217
rect 27433 25171 27491 25177
rect 46477 25177 46489 25211
rect 46523 25208 46535 25211
rect 47670 25208 47676 25220
rect 46523 25180 47676 25208
rect 46523 25177 46535 25180
rect 46477 25171 46535 25177
rect 47670 25168 47676 25180
rect 47728 25168 47734 25220
rect 21600 25112 22248 25140
rect 21600 25100 21606 25112
rect 24946 25100 24952 25152
rect 25004 25140 25010 25152
rect 25593 25143 25651 25149
rect 25593 25140 25605 25143
rect 25004 25112 25605 25140
rect 25004 25100 25010 25112
rect 25593 25109 25605 25112
rect 25639 25109 25651 25143
rect 25593 25103 25651 25109
rect 26973 25143 27031 25149
rect 26973 25109 26985 25143
rect 27019 25140 27031 25143
rect 27706 25140 27712 25152
rect 27019 25112 27712 25140
rect 27019 25109 27031 25112
rect 26973 25103 27031 25109
rect 27706 25100 27712 25112
rect 27764 25100 27770 25152
rect 28445 25143 28503 25149
rect 28445 25109 28457 25143
rect 28491 25140 28503 25143
rect 29454 25140 29460 25152
rect 28491 25112 29460 25140
rect 28491 25109 28503 25112
rect 28445 25103 28503 25109
rect 29454 25100 29460 25112
rect 29512 25100 29518 25152
rect 30558 25100 30564 25152
rect 30616 25140 30622 25152
rect 30653 25143 30711 25149
rect 30653 25140 30665 25143
rect 30616 25112 30665 25140
rect 30616 25100 30622 25112
rect 30653 25109 30665 25112
rect 30699 25109 30711 25143
rect 30653 25103 30711 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 13906 24896 13912 24948
rect 13964 24936 13970 24948
rect 14553 24939 14611 24945
rect 14553 24936 14565 24939
rect 13964 24908 14565 24936
rect 13964 24896 13970 24908
rect 14553 24905 14565 24908
rect 14599 24905 14611 24939
rect 15838 24936 15844 24948
rect 15799 24908 15844 24936
rect 14553 24899 14611 24905
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 15933 24939 15991 24945
rect 15933 24905 15945 24939
rect 15979 24936 15991 24939
rect 16298 24936 16304 24948
rect 15979 24908 16304 24936
rect 15979 24905 15991 24908
rect 15933 24899 15991 24905
rect 16298 24896 16304 24908
rect 16356 24896 16362 24948
rect 16850 24936 16856 24948
rect 16811 24908 16856 24936
rect 16850 24896 16856 24908
rect 16908 24896 16914 24948
rect 22094 24896 22100 24948
rect 22152 24936 22158 24948
rect 22152 24908 22197 24936
rect 22152 24896 22158 24908
rect 29822 24896 29828 24948
rect 29880 24936 29886 24948
rect 30929 24939 30987 24945
rect 30929 24936 30941 24939
rect 29880 24908 30941 24936
rect 29880 24896 29886 24908
rect 30929 24905 30941 24908
rect 30975 24905 30987 24939
rect 30929 24899 30987 24905
rect 13262 24828 13268 24880
rect 13320 24868 13326 24880
rect 15749 24871 15807 24877
rect 15749 24868 15761 24871
rect 13320 24840 15761 24868
rect 13320 24828 13326 24840
rect 15749 24837 15761 24840
rect 15795 24837 15807 24871
rect 15749 24831 15807 24837
rect 46750 24828 46756 24880
rect 46808 24828 46814 24880
rect 8297 24803 8355 24809
rect 8297 24769 8309 24803
rect 8343 24800 8355 24803
rect 8478 24800 8484 24812
rect 8343 24772 8484 24800
rect 8343 24769 8355 24772
rect 8297 24763 8355 24769
rect 8478 24760 8484 24772
rect 8536 24760 8542 24812
rect 10226 24760 10232 24812
rect 10284 24760 10290 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 13173 24803 13231 24809
rect 13173 24800 13185 24803
rect 12860 24772 13185 24800
rect 12860 24760 12866 24772
rect 13173 24769 13185 24772
rect 13219 24800 13231 24803
rect 13354 24800 13360 24812
rect 13219 24772 13360 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 13354 24760 13360 24772
rect 13412 24800 13418 24812
rect 13817 24803 13875 24809
rect 13817 24800 13829 24803
rect 13412 24772 13829 24800
rect 13412 24760 13418 24772
rect 13817 24769 13829 24772
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 14001 24803 14059 24809
rect 14001 24769 14013 24803
rect 14047 24800 14059 24803
rect 14366 24800 14372 24812
rect 14047 24772 14372 24800
rect 14047 24769 14059 24772
rect 14001 24763 14059 24769
rect 14366 24760 14372 24772
rect 14424 24760 14430 24812
rect 14458 24760 14464 24812
rect 14516 24800 14522 24812
rect 14516 24772 14561 24800
rect 14516 24760 14522 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 15436 24772 15577 24800
rect 15436 24760 15442 24772
rect 15565 24769 15577 24772
rect 15611 24769 15623 24803
rect 16666 24800 16672 24812
rect 16627 24772 16672 24800
rect 15565 24763 15623 24769
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 18230 24800 18236 24812
rect 18191 24772 18236 24800
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24800 18383 24803
rect 18414 24800 18420 24812
rect 18371 24772 18420 24800
rect 18371 24769 18383 24772
rect 18325 24763 18383 24769
rect 18414 24760 18420 24772
rect 18472 24760 18478 24812
rect 22465 24803 22523 24809
rect 22465 24769 22477 24803
rect 22511 24769 22523 24803
rect 22465 24763 22523 24769
rect 8389 24735 8447 24741
rect 8389 24701 8401 24735
rect 8435 24732 8447 24735
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 8435 24704 8861 24732
rect 8435 24701 8447 24704
rect 8389 24695 8447 24701
rect 8849 24701 8861 24704
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 9125 24735 9183 24741
rect 9125 24701 9137 24735
rect 9171 24732 9183 24735
rect 10134 24732 10140 24744
rect 9171 24704 10140 24732
rect 9171 24701 9183 24704
rect 9125 24695 9183 24701
rect 10134 24692 10140 24704
rect 10192 24692 10198 24744
rect 16390 24732 16396 24744
rect 13372 24704 16396 24732
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 12158 24664 12164 24676
rect 10376 24636 12164 24664
rect 10376 24624 10382 24636
rect 12158 24624 12164 24636
rect 12216 24664 12222 24676
rect 13372 24673 13400 24704
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 18506 24692 18512 24744
rect 18564 24732 18570 24744
rect 18969 24735 19027 24741
rect 18969 24732 18981 24735
rect 18564 24704 18981 24732
rect 18564 24692 18570 24704
rect 18969 24701 18981 24704
rect 19015 24701 19027 24735
rect 18969 24695 19027 24701
rect 19153 24735 19211 24741
rect 19153 24701 19165 24735
rect 19199 24732 19211 24735
rect 19334 24732 19340 24744
rect 19199 24704 19340 24732
rect 19199 24701 19211 24704
rect 19153 24695 19211 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24732 20867 24735
rect 22278 24732 22284 24744
rect 20855 24704 22284 24732
rect 20855 24701 20867 24704
rect 20809 24695 20867 24701
rect 22278 24692 22284 24704
rect 22336 24692 22342 24744
rect 22480 24732 22508 24763
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 22612 24772 22657 24800
rect 22612 24760 22618 24772
rect 24670 24760 24676 24812
rect 24728 24760 24734 24812
rect 27614 24800 27620 24812
rect 27575 24772 27620 24800
rect 27614 24760 27620 24772
rect 27672 24760 27678 24812
rect 30558 24760 30564 24812
rect 30616 24760 30622 24812
rect 46566 24760 46572 24812
rect 46624 24800 46630 24812
rect 46768 24800 46796 24828
rect 46845 24803 46903 24809
rect 46845 24800 46857 24803
rect 46624 24772 46857 24800
rect 46624 24760 46630 24772
rect 46845 24769 46857 24772
rect 46891 24769 46903 24803
rect 46845 24763 46903 24769
rect 47486 24760 47492 24812
rect 47544 24800 47550 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47544 24772 47593 24800
rect 47544 24760 47550 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 47670 24760 47676 24812
rect 47728 24800 47734 24812
rect 47728 24772 47773 24800
rect 47728 24760 47734 24772
rect 22741 24735 22799 24741
rect 22480 24704 22600 24732
rect 13357 24667 13415 24673
rect 13357 24664 13369 24667
rect 12216 24636 13369 24664
rect 12216 24624 12222 24636
rect 13357 24633 13369 24636
rect 13403 24633 13415 24667
rect 13357 24627 13415 24633
rect 16117 24667 16175 24673
rect 16117 24633 16129 24667
rect 16163 24664 16175 24667
rect 20438 24664 20444 24676
rect 16163 24636 20444 24664
rect 16163 24633 16175 24636
rect 16117 24627 16175 24633
rect 20438 24624 20444 24636
rect 20496 24624 20502 24676
rect 22572 24664 22600 24704
rect 22741 24701 22753 24735
rect 22787 24732 22799 24735
rect 22922 24732 22928 24744
rect 22787 24704 22928 24732
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 22922 24692 22928 24704
rect 22980 24692 22986 24744
rect 23290 24732 23296 24744
rect 23251 24704 23296 24732
rect 23290 24692 23296 24704
rect 23348 24692 23354 24744
rect 23566 24732 23572 24744
rect 23527 24704 23572 24732
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 26234 24732 26240 24744
rect 25087 24704 26240 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 27706 24732 27712 24744
rect 27619 24704 27712 24732
rect 27706 24692 27712 24704
rect 27764 24732 27770 24744
rect 28902 24732 28908 24744
rect 27764 24704 28908 24732
rect 27764 24692 27770 24704
rect 28902 24692 28908 24704
rect 28960 24692 28966 24744
rect 29178 24732 29184 24744
rect 29139 24704 29184 24732
rect 29178 24692 29184 24704
rect 29236 24692 29242 24744
rect 29454 24732 29460 24744
rect 29415 24704 29460 24732
rect 29454 24692 29460 24704
rect 29512 24692 29518 24744
rect 46750 24732 46756 24744
rect 30484 24704 46756 24732
rect 22572 24636 22784 24664
rect 22756 24608 22784 24636
rect 25958 24624 25964 24676
rect 26016 24664 26022 24676
rect 26016 24636 29316 24664
rect 26016 24624 26022 24636
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 10597 24599 10655 24605
rect 10597 24596 10609 24599
rect 9364 24568 10609 24596
rect 9364 24556 9370 24568
rect 10597 24565 10609 24568
rect 10643 24565 10655 24599
rect 13906 24596 13912 24608
rect 13867 24568 13912 24596
rect 10597 24559 10655 24565
rect 13906 24556 13912 24568
rect 13964 24556 13970 24608
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 16666 24596 16672 24608
rect 14516 24568 16672 24596
rect 14516 24556 14522 24568
rect 16666 24556 16672 24568
rect 16724 24556 16730 24608
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 23109 24599 23167 24605
rect 23109 24596 23121 24599
rect 22796 24568 23121 24596
rect 22796 24556 22802 24568
rect 23109 24565 23121 24568
rect 23155 24565 23167 24599
rect 23109 24559 23167 24565
rect 27893 24599 27951 24605
rect 27893 24565 27905 24599
rect 27939 24596 27951 24599
rect 28994 24596 29000 24608
rect 27939 24568 29000 24596
rect 27939 24565 27951 24568
rect 27893 24559 27951 24565
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29288 24596 29316 24636
rect 30484 24596 30512 24704
rect 46750 24692 46756 24704
rect 46808 24692 46814 24744
rect 29288 24568 30512 24596
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 46937 24599 46995 24605
rect 46937 24596 46949 24599
rect 46532 24568 46949 24596
rect 46532 24556 46538 24568
rect 46937 24565 46949 24568
rect 46983 24565 46995 24599
rect 46937 24559 46995 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 9953 24395 10011 24401
rect 9953 24361 9965 24395
rect 9999 24392 10011 24395
rect 10226 24392 10232 24404
rect 9999 24364 10232 24392
rect 9999 24361 10011 24364
rect 9953 24355 10011 24361
rect 10226 24352 10232 24364
rect 10284 24352 10290 24404
rect 15286 24352 15292 24404
rect 15344 24392 15350 24404
rect 18506 24392 18512 24404
rect 15344 24364 18512 24392
rect 15344 24352 15350 24364
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 19797 24395 19855 24401
rect 19797 24361 19809 24395
rect 19843 24392 19855 24395
rect 20622 24392 20628 24404
rect 19843 24364 20628 24392
rect 19843 24361 19855 24364
rect 19797 24355 19855 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 22002 24352 22008 24404
rect 22060 24392 22066 24404
rect 22097 24395 22155 24401
rect 22097 24392 22109 24395
rect 22060 24364 22109 24392
rect 22060 24352 22066 24364
rect 22097 24361 22109 24364
rect 22143 24361 22155 24395
rect 22097 24355 22155 24361
rect 22278 24352 22284 24404
rect 22336 24392 22342 24404
rect 26421 24395 26479 24401
rect 22336 24364 26004 24392
rect 22336 24352 22342 24364
rect 25976 24324 26004 24364
rect 26421 24361 26433 24395
rect 26467 24392 26479 24395
rect 26786 24392 26792 24404
rect 26467 24364 26792 24392
rect 26467 24361 26479 24364
rect 26421 24355 26479 24361
rect 26786 24352 26792 24364
rect 26844 24352 26850 24404
rect 27525 24395 27583 24401
rect 27525 24361 27537 24395
rect 27571 24392 27583 24395
rect 27982 24392 27988 24404
rect 27571 24364 27988 24392
rect 27571 24361 27583 24364
rect 27525 24355 27583 24361
rect 27982 24352 27988 24364
rect 28040 24352 28046 24404
rect 28537 24395 28595 24401
rect 28537 24361 28549 24395
rect 28583 24392 28595 24395
rect 28718 24392 28724 24404
rect 28583 24364 28724 24392
rect 28583 24361 28595 24364
rect 28537 24355 28595 24361
rect 28718 24352 28724 24364
rect 28776 24352 28782 24404
rect 28902 24352 28908 24404
rect 28960 24392 28966 24404
rect 29914 24392 29920 24404
rect 28960 24364 29005 24392
rect 29875 24364 29920 24392
rect 28960 24352 28966 24364
rect 29914 24352 29920 24364
rect 29972 24352 29978 24404
rect 46382 24392 46388 24404
rect 31726 24364 46388 24392
rect 31726 24324 31754 24364
rect 46382 24352 46388 24364
rect 46440 24352 46446 24404
rect 25976 24296 31754 24324
rect 16025 24259 16083 24265
rect 16025 24225 16037 24259
rect 16071 24256 16083 24259
rect 17037 24259 17095 24265
rect 17037 24256 17049 24259
rect 16071 24228 17049 24256
rect 16071 24225 16083 24228
rect 16025 24219 16083 24225
rect 17037 24225 17049 24228
rect 17083 24225 17095 24259
rect 17037 24219 17095 24225
rect 19426 24216 19432 24268
rect 19484 24256 19490 24268
rect 20349 24259 20407 24265
rect 20349 24256 20361 24259
rect 19484 24228 20361 24256
rect 19484 24216 19490 24228
rect 20349 24225 20361 24228
rect 20395 24256 20407 24259
rect 23290 24256 23296 24268
rect 20395 24228 23296 24256
rect 20395 24225 20407 24228
rect 20349 24219 20407 24225
rect 23290 24216 23296 24228
rect 23348 24256 23354 24268
rect 24673 24259 24731 24265
rect 24673 24256 24685 24259
rect 23348 24228 24685 24256
rect 23348 24216 23354 24228
rect 24673 24225 24685 24228
rect 24719 24225 24731 24259
rect 24946 24256 24952 24268
rect 24907 24228 24952 24256
rect 24673 24219 24731 24225
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 27614 24216 27620 24268
rect 27672 24256 27678 24268
rect 27985 24259 28043 24265
rect 27985 24256 27997 24259
rect 27672 24228 27997 24256
rect 27672 24216 27678 24228
rect 27985 24225 27997 24228
rect 28031 24225 28043 24259
rect 27985 24219 28043 24225
rect 28276 24228 28856 24256
rect 9858 24188 9864 24200
rect 9819 24160 9864 24188
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12894 24188 12900 24200
rect 12492 24160 12900 24188
rect 12492 24148 12498 24160
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 15838 24188 15844 24200
rect 13219 24160 15700 24188
rect 15799 24160 15844 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 13354 24120 13360 24132
rect 13315 24092 13360 24120
rect 13354 24080 13360 24092
rect 13412 24080 13418 24132
rect 15672 24120 15700 24160
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 16390 24188 16396 24200
rect 16347 24160 16396 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 16390 24148 16396 24160
rect 16448 24148 16454 24200
rect 16758 24188 16764 24200
rect 16719 24160 16764 24188
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 18322 24120 18328 24132
rect 15672 24092 17448 24120
rect 18262 24092 18328 24120
rect 12526 24052 12532 24064
rect 12487 24024 12532 24052
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 16209 24055 16267 24061
rect 16209 24021 16221 24055
rect 16255 24052 16267 24055
rect 16298 24052 16304 24064
rect 16255 24024 16304 24052
rect 16255 24021 16267 24024
rect 16209 24015 16267 24021
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 17420 24052 17448 24092
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 19628 24120 19656 24151
rect 20530 24120 20536 24132
rect 19628 24092 20536 24120
rect 19628 24052 19656 24092
rect 20530 24080 20536 24092
rect 20588 24080 20594 24132
rect 20625 24123 20683 24129
rect 20625 24089 20637 24123
rect 20671 24089 20683 24123
rect 20625 24083 20683 24089
rect 17420 24024 19656 24052
rect 20640 24052 20668 24083
rect 21082 24080 21088 24132
rect 21140 24080 21146 24132
rect 25682 24080 25688 24132
rect 25740 24080 25746 24132
rect 21358 24052 21364 24064
rect 20640 24024 21364 24052
rect 21358 24012 21364 24024
rect 21416 24012 21422 24064
rect 27724 24052 27752 24151
rect 27798 24148 27804 24200
rect 27856 24188 27862 24200
rect 28077 24191 28135 24197
rect 27856 24160 27901 24188
rect 27856 24148 27862 24160
rect 28077 24157 28089 24191
rect 28123 24188 28135 24191
rect 28276 24188 28304 24228
rect 28123 24160 28304 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 28442 24148 28448 24200
rect 28500 24188 28506 24200
rect 28721 24191 28779 24197
rect 28721 24188 28733 24191
rect 28500 24160 28733 24188
rect 28500 24148 28506 24160
rect 28721 24157 28733 24160
rect 28767 24157 28779 24191
rect 28828 24188 28856 24228
rect 28902 24216 28908 24268
rect 28960 24256 28966 24268
rect 28997 24259 29055 24265
rect 28997 24256 29009 24259
rect 28960 24228 29009 24256
rect 28960 24216 28966 24228
rect 28997 24225 29009 24228
rect 29043 24225 29055 24259
rect 30009 24259 30067 24265
rect 28997 24219 29055 24225
rect 29104 24228 29868 24256
rect 29104 24188 29132 24228
rect 28828 24160 29132 24188
rect 29733 24191 29791 24197
rect 28721 24151 28779 24157
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 29840 24188 29868 24228
rect 30009 24225 30021 24259
rect 30055 24256 30067 24259
rect 30282 24256 30288 24268
rect 30055 24228 30288 24256
rect 30055 24225 30067 24228
rect 30009 24219 30067 24225
rect 30282 24216 30288 24228
rect 30340 24216 30346 24268
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 30098 24188 30104 24200
rect 29840 24160 30104 24188
rect 29733 24151 29791 24157
rect 27982 24080 27988 24132
rect 28040 24120 28046 24132
rect 29748 24120 29776 24151
rect 30098 24148 30104 24160
rect 30156 24148 30162 24200
rect 46293 24191 46351 24197
rect 46293 24157 46305 24191
rect 46339 24157 46351 24191
rect 46293 24151 46351 24157
rect 28040 24092 29776 24120
rect 46308 24120 46336 24151
rect 47762 24120 47768 24132
rect 46308 24092 47768 24120
rect 28040 24080 28046 24092
rect 47762 24080 47768 24092
rect 47820 24080 47826 24132
rect 29270 24052 29276 24064
rect 27724 24024 29276 24052
rect 29270 24012 29276 24024
rect 29328 24012 29334 24064
rect 29546 24052 29552 24064
rect 29507 24024 29552 24052
rect 29546 24012 29552 24024
rect 29604 24012 29610 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 1762 23848 1768 23860
rect 1627 23820 1768 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 1762 23808 1768 23820
rect 1820 23808 1826 23860
rect 12802 23848 12808 23860
rect 12763 23820 12808 23848
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 14366 23808 14372 23860
rect 14424 23848 14430 23860
rect 14553 23851 14611 23857
rect 14553 23848 14565 23851
rect 14424 23820 14565 23848
rect 14424 23808 14430 23820
rect 14553 23817 14565 23820
rect 14599 23848 14611 23851
rect 15657 23851 15715 23857
rect 15657 23848 15669 23851
rect 14599 23820 15669 23848
rect 14599 23817 14611 23820
rect 14553 23811 14611 23817
rect 15657 23817 15669 23820
rect 15703 23817 15715 23851
rect 15657 23811 15715 23817
rect 15841 23851 15899 23857
rect 15841 23817 15853 23851
rect 15887 23848 15899 23851
rect 16298 23848 16304 23860
rect 15887 23820 16304 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 16853 23851 16911 23857
rect 16853 23848 16865 23851
rect 16816 23820 16865 23848
rect 16816 23808 16822 23820
rect 16853 23817 16865 23820
rect 16899 23817 16911 23851
rect 18322 23848 18328 23860
rect 18283 23820 18328 23848
rect 16853 23811 16911 23817
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 24397 23851 24455 23857
rect 24397 23817 24409 23851
rect 24443 23848 24455 23851
rect 24670 23848 24676 23860
rect 24443 23820 24676 23848
rect 24443 23817 24455 23820
rect 24397 23811 24455 23817
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 27890 23808 27896 23860
rect 27948 23848 27954 23860
rect 28721 23851 28779 23857
rect 28721 23848 28733 23851
rect 27948 23820 28733 23848
rect 27948 23808 27954 23820
rect 28721 23817 28733 23820
rect 28767 23848 28779 23851
rect 28902 23848 28908 23860
rect 28767 23820 28908 23848
rect 28767 23817 28779 23820
rect 28721 23811 28779 23817
rect 28902 23808 28908 23820
rect 28960 23808 28966 23860
rect 9306 23740 9312 23792
rect 9364 23780 9370 23792
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 9364 23752 9413 23780
rect 9364 23740 9370 23752
rect 9401 23749 9413 23752
rect 9447 23780 9459 23783
rect 11517 23783 11575 23789
rect 11517 23780 11529 23783
rect 9447 23752 11529 23780
rect 9447 23749 9459 23752
rect 9401 23743 9459 23749
rect 11517 23749 11529 23752
rect 11563 23749 11575 23783
rect 11517 23743 11575 23749
rect 11733 23783 11791 23789
rect 11733 23749 11745 23783
rect 11779 23780 11791 23783
rect 12066 23780 12072 23792
rect 11779 23752 12072 23780
rect 11779 23749 11791 23752
rect 11733 23743 11791 23749
rect 12066 23740 12072 23752
rect 12124 23740 12130 23792
rect 13633 23783 13691 23789
rect 13633 23780 13645 23783
rect 12636 23752 13645 23780
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 8478 23712 8484 23724
rect 8439 23684 8484 23712
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23681 9643 23715
rect 9585 23675 9643 23681
rect 9122 23604 9128 23656
rect 9180 23644 9186 23656
rect 9600 23644 9628 23675
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 9732 23684 9777 23712
rect 9732 23672 9738 23684
rect 9858 23672 9864 23724
rect 9916 23712 9922 23724
rect 12636 23721 12664 23752
rect 13633 23749 13645 23752
rect 13679 23780 13691 23783
rect 14645 23783 14703 23789
rect 14645 23780 14657 23783
rect 13679 23752 14657 23780
rect 13679 23749 13691 23752
rect 13633 23743 13691 23749
rect 14645 23749 14657 23752
rect 14691 23749 14703 23783
rect 15286 23780 15292 23792
rect 15247 23752 15292 23780
rect 14645 23743 14703 23749
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 26329 23783 26387 23789
rect 26329 23749 26341 23783
rect 26375 23780 26387 23783
rect 45370 23780 45376 23792
rect 26375 23752 27738 23780
rect 45331 23752 45376 23780
rect 26375 23749 26387 23752
rect 26329 23743 26387 23749
rect 45370 23740 45376 23752
rect 45428 23740 45434 23792
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 9916 23684 10149 23712
rect 9916 23672 9922 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 13262 23712 13268 23724
rect 13223 23684 13268 23712
rect 12621 23675 12679 23681
rect 13262 23672 13268 23684
rect 13320 23672 13326 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13538 23712 13544 23724
rect 13495 23684 13544 23712
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 13740 23684 14473 23712
rect 12437 23647 12495 23653
rect 9180 23616 10456 23644
rect 9180 23604 9186 23616
rect 9401 23579 9459 23585
rect 9401 23545 9413 23579
rect 9447 23576 9459 23579
rect 10042 23576 10048 23588
rect 9447 23548 10048 23576
rect 9447 23545 9459 23548
rect 9401 23539 9459 23545
rect 10042 23536 10048 23548
rect 10100 23536 10106 23588
rect 10428 23520 10456 23616
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12526 23644 12532 23656
rect 12483 23616 12532 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12526 23604 12532 23616
rect 12584 23644 12590 23656
rect 13740 23644 13768 23684
rect 14461 23681 14473 23684
rect 14507 23712 14519 23715
rect 15194 23712 15200 23724
rect 14507 23684 15200 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 15470 23712 15476 23724
rect 15431 23684 15476 23712
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 15565 23675 15623 23681
rect 12584 23616 13768 23644
rect 12584 23604 12590 23616
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14277 23647 14335 23653
rect 14277 23644 14289 23647
rect 13872 23616 14289 23644
rect 13872 23604 13878 23616
rect 14277 23613 14289 23616
rect 14323 23644 14335 23647
rect 15102 23644 15108 23656
rect 14323 23616 15108 23644
rect 14323 23613 14335 23616
rect 14277 23607 14335 23613
rect 15102 23604 15108 23616
rect 15160 23644 15166 23656
rect 15580 23644 15608 23675
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 18230 23712 18236 23724
rect 18191 23684 18236 23712
rect 18230 23672 18236 23684
rect 18288 23672 18294 23724
rect 18877 23715 18935 23721
rect 18877 23681 18889 23715
rect 18923 23712 18935 23715
rect 19978 23712 19984 23724
rect 18923 23684 19984 23712
rect 18923 23681 18935 23684
rect 18877 23675 18935 23681
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 24305 23715 24363 23721
rect 24305 23681 24317 23715
rect 24351 23712 24363 23715
rect 24670 23712 24676 23724
rect 24351 23684 24676 23712
rect 24351 23681 24363 23684
rect 24305 23675 24363 23681
rect 24670 23672 24676 23684
rect 24728 23712 24734 23724
rect 25593 23715 25651 23721
rect 25593 23712 25605 23715
rect 24728 23684 25605 23712
rect 24728 23672 24734 23684
rect 25593 23681 25605 23684
rect 25639 23712 25651 23715
rect 26237 23715 26295 23721
rect 26237 23712 26249 23715
rect 25639 23684 26249 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 26237 23681 26249 23684
rect 26283 23681 26295 23715
rect 26237 23675 26295 23681
rect 26973 23715 27031 23721
rect 26973 23681 26985 23715
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 15160 23616 15608 23644
rect 18248 23644 18276 23672
rect 19426 23644 19432 23656
rect 18248 23616 19432 23644
rect 15160 23604 15166 23616
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 13262 23576 13268 23588
rect 11931 23548 13268 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 13262 23536 13268 23548
rect 13320 23536 13326 23588
rect 15194 23536 15200 23588
rect 15252 23576 15258 23588
rect 15746 23576 15752 23588
rect 15252 23548 15752 23576
rect 15252 23536 15258 23548
rect 15746 23536 15752 23548
rect 15804 23536 15810 23588
rect 8297 23511 8355 23517
rect 8297 23477 8309 23511
rect 8343 23508 8355 23511
rect 8386 23508 8392 23520
rect 8343 23480 8392 23508
rect 8343 23477 8355 23480
rect 8297 23471 8355 23477
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 10134 23468 10140 23520
rect 10192 23508 10198 23520
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 10192 23480 10241 23508
rect 10192 23468 10198 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10229 23471 10287 23477
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 11701 23511 11759 23517
rect 11701 23508 11713 23511
rect 10468 23480 11713 23508
rect 10468 23468 10474 23480
rect 11701 23477 11713 23480
rect 11747 23477 11759 23511
rect 11701 23471 11759 23477
rect 14829 23511 14887 23517
rect 14829 23477 14841 23511
rect 14875 23508 14887 23511
rect 15930 23508 15936 23520
rect 14875 23480 15936 23508
rect 14875 23477 14887 23480
rect 14829 23471 14887 23477
rect 15930 23468 15936 23480
rect 15988 23468 15994 23520
rect 18966 23508 18972 23520
rect 18927 23480 18972 23508
rect 18966 23468 18972 23480
rect 19024 23468 19030 23520
rect 26988 23508 27016 23675
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 30006 23712 30012 23724
rect 28776 23684 30012 23712
rect 28776 23672 28782 23684
rect 30006 23672 30012 23684
rect 30064 23672 30070 23724
rect 47762 23712 47768 23724
rect 47723 23684 47768 23712
rect 47762 23672 47768 23684
rect 47820 23672 47826 23724
rect 27249 23647 27307 23653
rect 27249 23613 27261 23647
rect 27295 23644 27307 23647
rect 29546 23644 29552 23656
rect 27295 23616 29552 23644
rect 27295 23613 27307 23616
rect 27249 23607 27307 23613
rect 29546 23604 29552 23616
rect 29604 23604 29610 23656
rect 45189 23647 45247 23653
rect 45189 23613 45201 23647
rect 45235 23644 45247 23647
rect 45738 23644 45744 23656
rect 45235 23616 45744 23644
rect 45235 23613 45247 23616
rect 45189 23607 45247 23613
rect 45738 23604 45744 23616
rect 45796 23604 45802 23656
rect 46750 23644 46756 23656
rect 46711 23616 46756 23644
rect 46750 23604 46756 23616
rect 46808 23604 46814 23656
rect 29178 23508 29184 23520
rect 26988 23480 29184 23508
rect 29178 23468 29184 23480
rect 29236 23468 29242 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 9493 23307 9551 23313
rect 9493 23304 9505 23307
rect 8352 23276 9505 23304
rect 8352 23264 8358 23276
rect 9493 23273 9505 23276
rect 9539 23304 9551 23307
rect 9582 23304 9588 23316
rect 9539 23276 9588 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 10226 23304 10232 23316
rect 10187 23276 10232 23304
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 10410 23304 10416 23316
rect 10371 23276 10416 23304
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 11882 23304 11888 23316
rect 11843 23276 11888 23304
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 15838 23304 15844 23316
rect 15519 23276 15844 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 19426 23304 19432 23316
rect 19387 23276 19432 23304
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 22094 23304 22100 23316
rect 20916 23276 22100 23304
rect 2314 23196 2320 23248
rect 2372 23236 2378 23248
rect 2372 23208 15148 23236
rect 2372 23196 2378 23208
rect 9674 23168 9680 23180
rect 9508 23140 9680 23168
rect 9122 23100 9128 23112
rect 9083 23072 9128 23100
rect 9122 23060 9128 23072
rect 9180 23060 9186 23112
rect 8294 22924 8300 22976
rect 8352 22964 8358 22976
rect 8941 22967 8999 22973
rect 8941 22964 8953 22967
rect 8352 22936 8953 22964
rect 8352 22924 8358 22936
rect 8941 22933 8953 22936
rect 8987 22933 8999 22967
rect 8941 22927 8999 22933
rect 9125 22967 9183 22973
rect 9125 22933 9137 22967
rect 9171 22964 9183 22967
rect 9508 22964 9536 23140
rect 9674 23128 9680 23140
rect 9732 23168 9738 23180
rect 13265 23171 13323 23177
rect 9732 23140 11192 23168
rect 9732 23128 9738 23140
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 9766 23100 9772 23112
rect 9631 23072 9772 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 9766 23060 9772 23072
rect 9824 23100 9830 23112
rect 10594 23100 10600 23112
rect 9824 23072 10600 23100
rect 9824 23060 9830 23072
rect 10594 23060 10600 23072
rect 10652 23060 10658 23112
rect 10045 23035 10103 23041
rect 10045 23001 10057 23035
rect 10091 23001 10103 23035
rect 10962 23032 10968 23044
rect 10923 23004 10968 23032
rect 10045 22995 10103 23001
rect 9171 22936 9536 22964
rect 9171 22933 9183 22936
rect 9125 22927 9183 22933
rect 9582 22924 9588 22976
rect 9640 22964 9646 22976
rect 10060 22964 10088 22995
rect 10962 22992 10968 23004
rect 11020 22992 11026 23044
rect 11164 23041 11192 23140
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13906 23168 13912 23180
rect 13311 23140 13912 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15120 23168 15148 23208
rect 17954 23196 17960 23248
rect 18012 23236 18018 23248
rect 20916 23236 20944 23276
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 18012 23208 20944 23236
rect 18012 23196 18018 23208
rect 21082 23196 21088 23248
rect 21140 23236 21146 23248
rect 22005 23239 22063 23245
rect 22005 23236 22017 23239
rect 21140 23208 22017 23236
rect 21140 23196 21146 23208
rect 22005 23205 22017 23208
rect 22051 23205 22063 23239
rect 22005 23199 22063 23205
rect 27341 23171 27399 23177
rect 27341 23168 27353 23171
rect 15120 23140 27353 23168
rect 27341 23137 27353 23140
rect 27387 23137 27399 23171
rect 27341 23131 27399 23137
rect 45738 23128 45744 23180
rect 45796 23168 45802 23180
rect 46293 23171 46351 23177
rect 46293 23168 46305 23171
rect 45796 23140 46305 23168
rect 45796 23128 45802 23140
rect 46293 23137 46305 23140
rect 46339 23137 46351 23171
rect 46842 23168 46848 23180
rect 46803 23140 46848 23168
rect 46293 23131 46351 23137
rect 46842 23128 46848 23140
rect 46900 23128 46906 23180
rect 13173 23103 13231 23109
rect 13173 23069 13185 23103
rect 13219 23100 13231 23103
rect 13814 23100 13820 23112
rect 13219 23072 13820 23100
rect 13219 23069 13231 23072
rect 13173 23063 13231 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14458 23100 14464 23112
rect 14323 23072 14464 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14458 23060 14464 23072
rect 14516 23060 14522 23112
rect 14826 23100 14832 23112
rect 14787 23072 14832 23100
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15344 23072 15669 23100
rect 15344 23060 15350 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 15930 23100 15936 23112
rect 15891 23072 15936 23100
rect 15657 23063 15715 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 19242 23100 19248 23112
rect 19203 23072 19248 23100
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 20956 23072 22248 23100
rect 20956 23060 20962 23072
rect 11149 23035 11207 23041
rect 11149 23001 11161 23035
rect 11195 23032 11207 23035
rect 11238 23032 11244 23044
rect 11195 23004 11244 23032
rect 11195 23001 11207 23004
rect 11149 22995 11207 23001
rect 11238 22992 11244 23004
rect 11296 22992 11302 23044
rect 11790 23032 11796 23044
rect 11751 23004 11796 23032
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 12618 22992 12624 23044
rect 12676 23032 12682 23044
rect 13354 23032 13360 23044
rect 12676 23004 13360 23032
rect 12676 22992 12682 23004
rect 13354 22992 13360 23004
rect 13412 23032 13418 23044
rect 13412 23004 15056 23032
rect 13412 22992 13418 23004
rect 9640 22936 10088 22964
rect 9640 22924 9646 22936
rect 10226 22924 10232 22976
rect 10284 22973 10290 22976
rect 10284 22967 10303 22973
rect 10291 22933 10303 22967
rect 10284 22927 10303 22933
rect 13541 22967 13599 22973
rect 13541 22933 13553 22967
rect 13587 22964 13599 22967
rect 13630 22964 13636 22976
rect 13587 22936 13636 22964
rect 13587 22933 13599 22936
rect 13541 22927 13599 22933
rect 10284 22924 10290 22927
rect 13630 22924 13636 22936
rect 13688 22924 13694 22976
rect 14274 22964 14280 22976
rect 14235 22936 14280 22964
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14918 22964 14924 22976
rect 14879 22936 14924 22964
rect 14918 22924 14924 22936
rect 14976 22924 14982 22976
rect 15028 22964 15056 23004
rect 15470 22992 15476 23044
rect 15528 23032 15534 23044
rect 15841 23035 15899 23041
rect 15841 23032 15853 23035
rect 15528 23004 15853 23032
rect 15528 22992 15534 23004
rect 15841 23001 15853 23004
rect 15887 23001 15899 23035
rect 15841 22995 15899 23001
rect 16114 22992 16120 23044
rect 16172 23032 16178 23044
rect 20806 23032 20812 23044
rect 16172 23004 20812 23032
rect 16172 22992 16178 23004
rect 20806 22992 20812 23004
rect 20864 22992 20870 23044
rect 22002 23032 22008 23044
rect 21963 23004 22008 23032
rect 22002 22992 22008 23004
rect 22060 22992 22066 23044
rect 22220 23032 22248 23072
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 22741 23103 22799 23109
rect 22336 23072 22381 23100
rect 22336 23060 22342 23072
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 27154 23100 27160 23112
rect 27115 23072 27160 23100
rect 22741 23063 22799 23069
rect 22756 23032 22784 23063
rect 27154 23060 27160 23072
rect 27212 23060 27218 23112
rect 44453 23103 44511 23109
rect 44453 23069 44465 23103
rect 44499 23069 44511 23103
rect 44453 23063 44511 23069
rect 45373 23103 45431 23109
rect 45373 23069 45385 23103
rect 45419 23100 45431 23103
rect 45462 23100 45468 23112
rect 45419 23072 45468 23100
rect 45419 23069 45431 23072
rect 45373 23063 45431 23069
rect 22220 23004 22784 23032
rect 28997 23035 29055 23041
rect 28997 23001 29009 23035
rect 29043 23032 29055 23035
rect 30374 23032 30380 23044
rect 29043 23004 30380 23032
rect 29043 23001 29055 23004
rect 28997 22995 29055 23001
rect 30374 22992 30380 23004
rect 30432 22992 30438 23044
rect 44468 23032 44496 23063
rect 45462 23060 45468 23072
rect 45520 23060 45526 23112
rect 45557 23103 45615 23109
rect 45557 23069 45569 23103
rect 45603 23100 45615 23103
rect 45830 23100 45836 23112
rect 45603 23072 45836 23100
rect 45603 23069 45615 23072
rect 45557 23063 45615 23069
rect 45830 23060 45836 23072
rect 45888 23060 45894 23112
rect 46106 23032 46112 23044
rect 44468 23004 46112 23032
rect 46106 22992 46112 23004
rect 46164 22992 46170 23044
rect 46477 23035 46535 23041
rect 46477 23001 46489 23035
rect 46523 23032 46535 23035
rect 47670 23032 47676 23044
rect 46523 23004 47676 23032
rect 46523 23001 46535 23004
rect 46477 22995 46535 23001
rect 47670 22992 47676 23004
rect 47728 22992 47734 23044
rect 19242 22964 19248 22976
rect 15028 22936 19248 22964
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 22186 22964 22192 22976
rect 22147 22936 22192 22964
rect 22186 22924 22192 22936
rect 22244 22924 22250 22976
rect 22833 22967 22891 22973
rect 22833 22933 22845 22967
rect 22879 22964 22891 22967
rect 22922 22964 22928 22976
rect 22879 22936 22928 22964
rect 22879 22933 22891 22936
rect 22833 22927 22891 22933
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 42794 22924 42800 22976
rect 42852 22964 42858 22976
rect 44269 22967 44327 22973
rect 44269 22964 44281 22967
rect 42852 22936 44281 22964
rect 42852 22924 42858 22936
rect 44269 22933 44281 22936
rect 44315 22933 44327 22967
rect 44269 22927 44327 22933
rect 45186 22924 45192 22976
rect 45244 22964 45250 22976
rect 45465 22967 45523 22973
rect 45465 22964 45477 22967
rect 45244 22936 45477 22964
rect 45244 22924 45250 22936
rect 45465 22933 45477 22936
rect 45511 22933 45523 22967
rect 45465 22927 45523 22933
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 9582 22720 9588 22772
rect 9640 22760 9646 22772
rect 9769 22763 9827 22769
rect 9769 22760 9781 22763
rect 9640 22732 9781 22760
rect 9640 22720 9646 22732
rect 9769 22729 9781 22732
rect 9815 22729 9827 22763
rect 9769 22723 9827 22729
rect 10439 22763 10497 22769
rect 10439 22729 10451 22763
rect 10485 22760 10497 22763
rect 10962 22760 10968 22772
rect 10485 22732 10968 22760
rect 10485 22729 10497 22732
rect 10439 22723 10497 22729
rect 10962 22720 10968 22732
rect 11020 22760 11026 22772
rect 11977 22763 12035 22769
rect 11977 22760 11989 22763
rect 11020 22732 11989 22760
rect 11020 22720 11026 22732
rect 11977 22729 11989 22732
rect 12023 22729 12035 22763
rect 12894 22760 12900 22772
rect 11977 22723 12035 22729
rect 12406 22732 12900 22760
rect 8294 22692 8300 22704
rect 8255 22664 8300 22692
rect 8294 22652 8300 22664
rect 8352 22652 8358 22704
rect 10134 22692 10140 22704
rect 9522 22664 10140 22692
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 10229 22695 10287 22701
rect 10229 22661 10241 22695
rect 10275 22692 10287 22695
rect 10318 22692 10324 22704
rect 10275 22664 10324 22692
rect 10275 22661 10287 22664
rect 10229 22655 10287 22661
rect 10318 22652 10324 22664
rect 10376 22652 10382 22704
rect 11609 22695 11667 22701
rect 11609 22661 11621 22695
rect 11655 22661 11667 22695
rect 11609 22655 11667 22661
rect 11825 22695 11883 22701
rect 11825 22661 11837 22695
rect 11871 22692 11883 22695
rect 12406 22692 12434 22732
rect 12894 22720 12900 22732
rect 12952 22760 12958 22772
rect 13538 22760 13544 22772
rect 12952 22732 13544 22760
rect 12952 22720 12958 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 15102 22760 15108 22772
rect 15063 22732 15108 22760
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 23937 22763 23995 22769
rect 23937 22760 23949 22763
rect 22060 22732 23949 22760
rect 22060 22720 22066 22732
rect 23937 22729 23949 22732
rect 23983 22729 23995 22763
rect 23937 22723 23995 22729
rect 13630 22692 13636 22704
rect 11871 22664 12434 22692
rect 13591 22664 13636 22692
rect 11871 22661 11883 22664
rect 11825 22655 11883 22661
rect 11624 22624 11652 22655
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 14918 22692 14924 22704
rect 14858 22664 14924 22692
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 21177 22695 21235 22701
rect 21177 22661 21189 22695
rect 21223 22692 21235 22695
rect 22465 22695 22523 22701
rect 22465 22692 22477 22695
rect 21223 22664 22477 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 22465 22661 22477 22664
rect 22511 22661 22523 22695
rect 22465 22655 22523 22661
rect 22922 22652 22928 22704
rect 22980 22652 22986 22704
rect 12434 22624 12440 22636
rect 11624 22596 12440 22624
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12618 22624 12624 22636
rect 12579 22596 12624 22624
rect 12618 22584 12624 22596
rect 12676 22584 12682 22636
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22624 15899 22627
rect 16666 22624 16672 22636
rect 15887 22596 16672 22624
rect 15887 22593 15899 22596
rect 15841 22587 15899 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 18506 22624 18512 22636
rect 18467 22596 18512 22624
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22624 19395 22627
rect 19426 22624 19432 22636
rect 19383 22596 19432 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 19426 22584 19432 22596
rect 19484 22624 19490 22636
rect 20898 22624 20904 22636
rect 19484 22596 20904 22624
rect 19484 22584 19490 22596
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 21082 22624 21088 22636
rect 21043 22596 21088 22624
rect 21082 22584 21088 22596
rect 21140 22584 21146 22636
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 23952 22624 23980 22723
rect 27062 22720 27068 22772
rect 27120 22760 27126 22772
rect 47670 22760 47676 22772
rect 27120 22732 29500 22760
rect 47631 22732 47676 22760
rect 27120 22720 27126 22732
rect 26421 22695 26479 22701
rect 26421 22661 26433 22695
rect 26467 22692 26479 22695
rect 26467 22664 29408 22692
rect 26467 22661 26479 22664
rect 26421 22655 26479 22661
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 23952 22596 24593 22624
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 8021 22559 8079 22565
rect 8021 22525 8033 22559
rect 8067 22556 8079 22559
rect 8386 22556 8392 22568
rect 8067 22528 8392 22556
rect 8067 22525 8079 22528
rect 8021 22519 8079 22525
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 13357 22559 13415 22565
rect 13357 22525 13369 22559
rect 13403 22556 13415 22559
rect 14274 22556 14280 22568
rect 13403 22528 14280 22556
rect 13403 22525 13415 22528
rect 13357 22519 13415 22525
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 22189 22559 22247 22565
rect 22189 22525 22201 22559
rect 22235 22556 22247 22559
rect 22830 22556 22836 22568
rect 22235 22528 22836 22556
rect 22235 22525 22247 22528
rect 22189 22519 22247 22525
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 24765 22559 24823 22565
rect 24765 22525 24777 22559
rect 24811 22556 24823 22559
rect 24946 22556 24952 22568
rect 24811 22528 24952 22556
rect 24811 22525 24823 22528
rect 24765 22519 24823 22525
rect 24946 22516 24952 22528
rect 25004 22516 25010 22568
rect 27154 22516 27160 22568
rect 27212 22556 27218 22568
rect 27617 22559 27675 22565
rect 27617 22556 27629 22559
rect 27212 22528 27629 22556
rect 27212 22516 27218 22528
rect 27617 22525 27629 22528
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 27801 22559 27859 22565
rect 27801 22525 27813 22559
rect 27847 22556 27859 22559
rect 29270 22556 29276 22568
rect 27847 22528 29276 22556
rect 27847 22525 27859 22528
rect 27801 22519 27859 22525
rect 10594 22488 10600 22500
rect 10555 22460 10600 22488
rect 10594 22448 10600 22460
rect 10652 22448 10658 22500
rect 27632 22488 27660 22519
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 29380 22556 29408 22664
rect 29472 22633 29500 22732
rect 47670 22720 47676 22732
rect 47728 22720 47734 22772
rect 29457 22627 29515 22633
rect 29457 22593 29469 22627
rect 29503 22593 29515 22627
rect 44634 22624 44640 22636
rect 44595 22596 44640 22624
rect 29457 22587 29515 22593
rect 44634 22584 44640 22596
rect 44692 22584 44698 22636
rect 44910 22624 44916 22636
rect 44871 22596 44916 22624
rect 44910 22584 44916 22596
rect 44968 22584 44974 22636
rect 46477 22627 46535 22633
rect 46477 22624 46489 22627
rect 45526 22596 46489 22624
rect 40034 22556 40040 22568
rect 29380 22528 40040 22556
rect 40034 22516 40040 22528
rect 40092 22516 40098 22568
rect 45370 22516 45376 22568
rect 45428 22556 45434 22568
rect 45526 22556 45554 22596
rect 46477 22593 46489 22596
rect 46523 22593 46535 22627
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 46477 22587 46535 22593
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 46198 22556 46204 22568
rect 45428 22528 45554 22556
rect 46159 22528 46204 22556
rect 45428 22516 45434 22528
rect 46198 22516 46204 22528
rect 46256 22516 46262 22568
rect 45097 22491 45155 22497
rect 45097 22488 45109 22491
rect 27632 22460 45109 22488
rect 45097 22457 45109 22460
rect 45143 22457 45155 22491
rect 45097 22451 45155 22457
rect 10042 22380 10048 22432
rect 10100 22420 10106 22432
rect 10226 22420 10232 22432
rect 10100 22392 10232 22420
rect 10100 22380 10106 22392
rect 10226 22380 10232 22392
rect 10284 22420 10290 22432
rect 10413 22423 10471 22429
rect 10413 22420 10425 22423
rect 10284 22392 10425 22420
rect 10284 22380 10290 22392
rect 10413 22389 10425 22392
rect 10459 22389 10471 22423
rect 10413 22383 10471 22389
rect 11793 22423 11851 22429
rect 11793 22389 11805 22423
rect 11839 22420 11851 22423
rect 12066 22420 12072 22432
rect 11839 22392 12072 22420
rect 11839 22389 11851 22392
rect 11793 22383 11851 22389
rect 12066 22380 12072 22392
rect 12124 22380 12130 22432
rect 12805 22423 12863 22429
rect 12805 22389 12817 22423
rect 12851 22420 12863 22423
rect 14826 22420 14832 22432
rect 12851 22392 14832 22420
rect 12851 22389 12863 22392
rect 12805 22383 12863 22389
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 15657 22423 15715 22429
rect 15657 22420 15669 22423
rect 15252 22392 15669 22420
rect 15252 22380 15258 22392
rect 15657 22389 15669 22392
rect 15703 22389 15715 22423
rect 18690 22420 18696 22432
rect 18651 22392 18696 22420
rect 15657 22383 15715 22389
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 19429 22423 19487 22429
rect 19429 22389 19441 22423
rect 19475 22420 19487 22423
rect 19978 22420 19984 22432
rect 19475 22392 19984 22420
rect 19475 22389 19487 22392
rect 19429 22383 19487 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 14277 22219 14335 22225
rect 14277 22185 14289 22219
rect 14323 22216 14335 22219
rect 14458 22216 14464 22228
rect 14323 22188 14464 22216
rect 14323 22185 14335 22188
rect 14277 22179 14335 22185
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 22186 22216 22192 22228
rect 22147 22188 22192 22216
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 22830 22216 22836 22228
rect 22791 22188 22836 22216
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 8110 22040 8116 22092
rect 8168 22080 8174 22092
rect 11238 22080 11244 22092
rect 8168 22052 11244 22080
rect 8168 22040 8174 22052
rect 10152 22021 10180 22052
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 15194 22080 15200 22092
rect 11940 22052 12434 22080
rect 15155 22052 15200 22080
rect 11940 22040 11946 22052
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10594 22012 10600 22024
rect 10555 21984 10600 22012
rect 10137 21975 10195 21981
rect 9876 21944 9904 21975
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 12406 22012 12434 22052
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15562 22040 15568 22092
rect 15620 22080 15626 22092
rect 16482 22080 16488 22092
rect 15620 22052 16488 22080
rect 15620 22040 15626 22052
rect 16482 22040 16488 22052
rect 16540 22080 16546 22092
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16540 22052 16957 22080
rect 16540 22040 16546 22052
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 17954 22080 17960 22092
rect 17915 22052 17960 22080
rect 16945 22043 17003 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 18417 22083 18475 22089
rect 18417 22049 18429 22083
rect 18463 22080 18475 22083
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 18463 22052 19533 22080
rect 18463 22049 18475 22052
rect 18417 22043 18475 22049
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 19521 22043 19579 22049
rect 20993 22083 21051 22089
rect 20993 22049 21005 22083
rect 21039 22080 21051 22083
rect 22204 22080 22232 22176
rect 44910 22148 44916 22160
rect 44468 22120 44916 22148
rect 22554 22080 22560 22092
rect 21039 22052 22560 22080
rect 21039 22049 21051 22052
rect 20993 22043 21051 22049
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 12406 21984 14105 22012
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 21981 18107 22015
rect 18049 21975 18107 21981
rect 10870 21944 10876 21956
rect 9876 21916 10180 21944
rect 10831 21916 10876 21944
rect 9674 21876 9680 21888
rect 9635 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10152 21876 10180 21916
rect 10870 21904 10876 21916
rect 10928 21904 10934 21956
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 10318 21876 10324 21888
rect 10152 21848 10324 21876
rect 10318 21836 10324 21848
rect 10376 21876 10382 21888
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 10376 21848 12357 21876
rect 10376 21836 10382 21848
rect 12345 21845 12357 21848
rect 12391 21876 12403 21879
rect 12618 21876 12624 21888
rect 12391 21848 12624 21876
rect 12391 21845 12403 21848
rect 12345 21839 12403 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 14108 21876 14136 21975
rect 15470 21944 15476 21956
rect 15431 21916 15476 21944
rect 15470 21904 15476 21916
rect 15528 21904 15534 21956
rect 16758 21944 16764 21956
rect 16698 21916 16764 21944
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 17954 21876 17960 21888
rect 14108 21848 17960 21876
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18064 21876 18092 21975
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18748 21984 19257 22012
rect 18748 21972 18754 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 19978 21904 19984 21956
rect 20036 21904 20042 21956
rect 18230 21876 18236 21888
rect 18064 21848 18236 21876
rect 18230 21836 18236 21848
rect 18288 21876 18294 21888
rect 21008 21876 21036 22043
rect 22554 22040 22560 22052
rect 22612 22040 22618 22092
rect 24946 22080 24952 22092
rect 24907 22052 24952 22080
rect 24946 22040 24952 22052
rect 25004 22040 25010 22092
rect 27982 22040 27988 22092
rect 28040 22080 28046 22092
rect 28040 22052 28764 22080
rect 28040 22040 28046 22052
rect 21266 21972 21272 22024
rect 21324 22012 21330 22024
rect 22646 22012 22652 22024
rect 21324 21984 22652 22012
rect 21324 21972 21330 21984
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25130 22012 25136 22024
rect 24903 21984 25136 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 22002 21944 22008 21956
rect 21963 21916 22008 21944
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 22848 21944 22876 21975
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 25498 22012 25504 22024
rect 25459 21984 25504 22012
rect 25498 21972 25504 21984
rect 25556 21972 25562 22024
rect 28736 22021 28764 22052
rect 29362 22040 29368 22092
rect 29420 22080 29426 22092
rect 29733 22083 29791 22089
rect 29733 22080 29745 22083
rect 29420 22052 29745 22080
rect 29420 22040 29426 22052
rect 29733 22049 29745 22052
rect 29779 22049 29791 22083
rect 44361 22083 44419 22089
rect 29733 22043 29791 22049
rect 30944 22052 35894 22080
rect 27341 22015 27399 22021
rect 27341 21981 27353 22015
rect 27387 22012 27399 22015
rect 28721 22015 28779 22021
rect 27387 21984 28672 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 22112 21916 22876 21944
rect 25685 21947 25743 21953
rect 18288 21848 21036 21876
rect 18288 21836 18294 21848
rect 21910 21836 21916 21888
rect 21968 21876 21974 21888
rect 22112 21876 22140 21916
rect 25685 21913 25697 21947
rect 25731 21944 25743 21947
rect 26234 21944 26240 21956
rect 25731 21916 26240 21944
rect 25731 21913 25743 21916
rect 25685 21907 25743 21913
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 27522 21904 27528 21956
rect 27580 21944 27586 21956
rect 27893 21947 27951 21953
rect 27893 21944 27905 21947
rect 27580 21916 27905 21944
rect 27580 21904 27586 21916
rect 27893 21913 27905 21916
rect 27939 21913 27951 21947
rect 28644 21944 28672 21984
rect 28721 21981 28733 22015
rect 28767 21981 28779 22015
rect 29546 22012 29552 22024
rect 29507 21984 29552 22012
rect 28721 21975 28779 21981
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 30944 21944 30972 22052
rect 35866 22012 35894 22052
rect 44361 22049 44373 22083
rect 44407 22080 44419 22083
rect 44468 22080 44496 22120
rect 44910 22108 44916 22120
rect 44968 22108 44974 22160
rect 44407 22052 44496 22080
rect 46293 22083 46351 22089
rect 44407 22049 44419 22052
rect 44361 22043 44419 22049
rect 46293 22049 46305 22083
rect 46339 22080 46351 22083
rect 46566 22080 46572 22092
rect 46339 22052 46572 22080
rect 46339 22049 46351 22052
rect 46293 22043 46351 22049
rect 46566 22040 46572 22052
rect 46624 22040 46630 22092
rect 46658 22040 46664 22092
rect 46716 22080 46722 22092
rect 46937 22083 46995 22089
rect 46937 22080 46949 22083
rect 46716 22052 46949 22080
rect 46716 22040 46722 22052
rect 46937 22049 46949 22052
rect 46983 22049 46995 22083
rect 46937 22043 46995 22049
rect 37274 22012 37280 22024
rect 35866 21984 37280 22012
rect 37274 21972 37280 21984
rect 37332 21972 37338 22024
rect 43438 22012 43444 22024
rect 43399 21984 43444 22012
rect 43438 21972 43444 21984
rect 43496 21972 43502 22024
rect 43622 22012 43628 22024
rect 43583 21984 43628 22012
rect 43622 21972 43628 21984
rect 43680 21972 43686 22024
rect 45278 22012 45284 22024
rect 45239 21984 45284 22012
rect 45278 21972 45284 21984
rect 45336 21972 45342 22024
rect 45557 22015 45615 22021
rect 45557 22012 45569 22015
rect 45388 21984 45569 22012
rect 28644 21916 30972 21944
rect 31389 21947 31447 21953
rect 27893 21907 27951 21913
rect 31389 21913 31401 21947
rect 31435 21944 31447 21947
rect 39574 21944 39580 21956
rect 31435 21916 39580 21944
rect 31435 21913 31447 21916
rect 31389 21907 31447 21913
rect 21968 21848 22140 21876
rect 21968 21836 21974 21848
rect 22186 21836 22192 21888
rect 22244 21885 22250 21888
rect 22244 21879 22263 21885
rect 22251 21845 22263 21879
rect 22244 21839 22263 21845
rect 22373 21879 22431 21885
rect 22373 21845 22385 21879
rect 22419 21876 22431 21879
rect 22646 21876 22652 21888
rect 22419 21848 22652 21876
rect 22419 21845 22431 21848
rect 22373 21839 22431 21845
rect 22244 21836 22250 21839
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 27982 21876 27988 21888
rect 27943 21848 27988 21876
rect 27982 21836 27988 21848
rect 28040 21836 28046 21888
rect 28810 21876 28816 21888
rect 28771 21848 28816 21876
rect 28810 21836 28816 21848
rect 28868 21836 28874 21888
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 31404 21876 31432 21907
rect 39574 21904 39580 21916
rect 39632 21904 39638 21956
rect 44450 21904 44456 21956
rect 44508 21944 44514 21956
rect 45186 21944 45192 21956
rect 44508 21916 45192 21944
rect 44508 21904 44514 21916
rect 45186 21904 45192 21916
rect 45244 21944 45250 21956
rect 45388 21944 45416 21984
rect 45557 21981 45569 21984
rect 45603 21981 45615 22015
rect 45557 21975 45615 21981
rect 45646 21944 45652 21956
rect 45244 21916 45416 21944
rect 45607 21916 45652 21944
rect 45244 21904 45250 21916
rect 45646 21904 45652 21916
rect 45704 21904 45710 21956
rect 46477 21947 46535 21953
rect 46477 21913 46489 21947
rect 46523 21944 46535 21947
rect 47670 21944 47676 21956
rect 46523 21916 47676 21944
rect 46523 21913 46535 21916
rect 46477 21907 46535 21913
rect 47670 21904 47676 21916
rect 47728 21904 47734 21956
rect 28960 21848 31432 21876
rect 28960 21836 28966 21848
rect 38562 21836 38568 21888
rect 38620 21876 38626 21888
rect 45922 21876 45928 21888
rect 38620 21848 45928 21876
rect 38620 21836 38626 21848
rect 45922 21836 45928 21848
rect 45980 21836 45986 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 10873 21675 10931 21681
rect 10873 21641 10885 21675
rect 10919 21672 10931 21675
rect 11330 21672 11336 21684
rect 10919 21644 11336 21672
rect 10919 21641 10931 21644
rect 10873 21635 10931 21641
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 16758 21672 16764 21684
rect 14884 21644 15516 21672
rect 16719 21644 16764 21672
rect 14884 21632 14890 21644
rect 9766 21604 9772 21616
rect 9727 21576 9772 21604
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 15378 21564 15384 21616
rect 15436 21564 15442 21616
rect 15488 21604 15516 21644
rect 16758 21632 16764 21644
rect 16816 21632 16822 21684
rect 21910 21672 21916 21684
rect 20088 21644 21916 21672
rect 15488 21576 16712 21604
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10781 21539 10839 21545
rect 10781 21536 10793 21539
rect 9916 21508 10793 21536
rect 9916 21496 9922 21508
rect 10781 21505 10793 21508
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 12434 21536 12440 21548
rect 11931 21508 12440 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 10045 21403 10103 21409
rect 10045 21400 10057 21403
rect 9732 21372 10057 21400
rect 9732 21360 9738 21372
rect 10045 21369 10057 21372
rect 10091 21369 10103 21403
rect 10796 21400 10824 21499
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21536 14427 21539
rect 15289 21539 15347 21545
rect 14415 21508 15240 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 12069 21403 12127 21409
rect 12069 21400 12081 21403
rect 10796 21372 12081 21400
rect 10045 21363 10103 21369
rect 12069 21369 12081 21372
rect 12115 21369 12127 21403
rect 12069 21363 12127 21369
rect 1578 21292 1584 21344
rect 1636 21332 1642 21344
rect 9950 21332 9956 21344
rect 1636 21304 9956 21332
rect 1636 21292 1642 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10229 21335 10287 21341
rect 10229 21301 10241 21335
rect 10275 21332 10287 21335
rect 10686 21332 10692 21344
rect 10275 21304 10692 21332
rect 10275 21301 10287 21304
rect 10229 21295 10287 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 14461 21335 14519 21341
rect 14461 21332 14473 21335
rect 14332 21304 14473 21332
rect 14332 21292 14338 21304
rect 14461 21301 14473 21304
rect 14507 21301 14519 21335
rect 15212 21332 15240 21508
rect 15289 21505 15301 21539
rect 15335 21536 15347 21539
rect 15396 21536 15424 21564
rect 16684 21545 16712 21576
rect 15335 21508 15424 21536
rect 16669 21539 16727 21545
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 16669 21505 16681 21539
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21505 17371 21539
rect 17313 21499 17371 21505
rect 15381 21471 15439 21477
rect 15381 21437 15393 21471
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 15396 21400 15424 21431
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 15528 21440 15669 21468
rect 15528 21428 15534 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 17328 21468 17356 21499
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18322 21536 18328 21548
rect 18012 21508 18328 21536
rect 18012 21496 18018 21508
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 20088 21536 20116 21644
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22060 21644 22477 21672
rect 22060 21632 22066 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 22554 21632 22560 21684
rect 22612 21672 22618 21684
rect 26234 21672 26240 21684
rect 22612 21644 22657 21672
rect 26195 21644 26240 21672
rect 22612 21632 22618 21644
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 27430 21632 27436 21684
rect 27488 21672 27494 21684
rect 28902 21672 28908 21684
rect 27488 21644 28908 21672
rect 27488 21632 27494 21644
rect 28902 21632 28908 21644
rect 28960 21632 28966 21684
rect 29270 21632 29276 21684
rect 29328 21672 29334 21684
rect 29917 21675 29975 21681
rect 29917 21672 29929 21675
rect 29328 21644 29929 21672
rect 29328 21632 29334 21644
rect 29917 21641 29929 21644
rect 29963 21641 29975 21675
rect 29917 21635 29975 21641
rect 43993 21675 44051 21681
rect 43993 21641 44005 21675
rect 44039 21672 44051 21675
rect 44450 21672 44456 21684
rect 44039 21644 44456 21672
rect 44039 21641 44051 21644
rect 43993 21635 44051 21641
rect 44450 21632 44456 21644
rect 44508 21632 44514 21684
rect 44634 21672 44640 21684
rect 44595 21644 44640 21672
rect 44634 21632 44640 21644
rect 44692 21632 44698 21684
rect 22373 21607 22431 21613
rect 22373 21604 22385 21607
rect 20272 21576 22385 21604
rect 20272 21548 20300 21576
rect 22373 21573 22385 21576
rect 22419 21573 22431 21607
rect 22373 21567 22431 21573
rect 27338 21564 27344 21616
rect 27396 21604 27402 21616
rect 42794 21604 42800 21616
rect 27396 21576 38700 21604
rect 27396 21564 27402 21576
rect 20254 21536 20260 21548
rect 19567 21508 20116 21536
rect 20215 21508 20260 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 18138 21468 18144 21480
rect 15657 21431 15715 21437
rect 16040 21440 18144 21468
rect 15930 21400 15936 21412
rect 15396 21372 15936 21400
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 16040 21332 16068 21440
rect 18138 21428 18144 21440
rect 18196 21428 18202 21480
rect 18506 21400 18512 21412
rect 18419 21372 18512 21400
rect 18506 21360 18512 21372
rect 18564 21400 18570 21412
rect 19536 21400 19564 21499
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20956 21508 21097 21536
rect 20956 21496 20962 21508
rect 21085 21505 21097 21508
rect 21131 21505 21143 21539
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 21085 21499 21143 21505
rect 22664 21508 23397 21536
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 20162 21468 20168 21480
rect 19668 21440 20168 21468
rect 19668 21428 19674 21440
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21468 20407 21471
rect 21266 21468 21272 21480
rect 20395 21440 21272 21468
rect 20395 21437 20407 21440
rect 20349 21431 20407 21437
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 22094 21428 22100 21480
rect 22152 21468 22158 21480
rect 22664 21468 22692 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25501 21539 25559 21545
rect 25501 21536 25513 21539
rect 25188 21508 25513 21536
rect 25188 21496 25194 21508
rect 25501 21505 25513 21508
rect 25547 21536 25559 21539
rect 26145 21539 26203 21545
rect 26145 21536 26157 21539
rect 25547 21508 26157 21536
rect 25547 21505 25559 21508
rect 25501 21499 25559 21505
rect 26145 21505 26157 21508
rect 26191 21505 26203 21539
rect 27522 21536 27528 21548
rect 27483 21508 27528 21536
rect 26145 21499 26203 21505
rect 27522 21496 27528 21508
rect 27580 21536 27586 21548
rect 28997 21539 29055 21545
rect 28997 21536 29009 21539
rect 27580 21508 29009 21536
rect 27580 21496 27586 21508
rect 28997 21505 29009 21508
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29365 21539 29423 21545
rect 29365 21505 29377 21539
rect 29411 21536 29423 21539
rect 29825 21539 29883 21545
rect 29825 21536 29837 21539
rect 29411 21508 29837 21536
rect 29411 21505 29423 21508
rect 29365 21499 29423 21505
rect 29825 21505 29837 21508
rect 29871 21536 29883 21539
rect 31386 21536 31392 21548
rect 29871 21508 31392 21536
rect 29871 21505 29883 21508
rect 29825 21499 29883 21505
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 22152 21440 22692 21468
rect 22741 21471 22799 21477
rect 22152 21428 22158 21440
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 23201 21471 23259 21477
rect 23201 21468 23213 21471
rect 22787 21440 23213 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 23201 21437 23213 21440
rect 23247 21437 23259 21471
rect 23201 21431 23259 21437
rect 24578 21428 24584 21480
rect 24636 21468 24642 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 24636 21440 28273 21468
rect 24636 21428 24642 21440
rect 28261 21437 28273 21440
rect 28307 21468 28319 21471
rect 28442 21468 28448 21480
rect 28307 21440 28448 21468
rect 28307 21437 28319 21440
rect 28261 21431 28319 21437
rect 28442 21428 28448 21440
rect 28500 21468 28506 21480
rect 28500 21440 31754 21468
rect 28500 21428 28506 21440
rect 22186 21400 22192 21412
rect 18564 21372 19564 21400
rect 22147 21372 22192 21400
rect 18564 21360 18570 21372
rect 22186 21360 22192 21372
rect 22244 21360 22250 21412
rect 31726 21400 31754 21440
rect 38562 21400 38568 21412
rect 31726 21372 38568 21400
rect 38562 21360 38568 21372
rect 38620 21360 38626 21412
rect 38672 21400 38700 21576
rect 39132 21576 42800 21604
rect 39132 21545 39160 21576
rect 42794 21564 42800 21576
rect 42852 21564 42858 21616
rect 45278 21604 45284 21616
rect 44284 21576 45284 21604
rect 39117 21539 39175 21545
rect 39117 21505 39129 21539
rect 39163 21505 39175 21539
rect 39117 21499 39175 21505
rect 39298 21468 39304 21480
rect 39259 21440 39304 21468
rect 39298 21428 39304 21440
rect 39356 21428 39362 21480
rect 39574 21468 39580 21480
rect 39535 21440 39580 21468
rect 39574 21428 39580 21440
rect 39632 21428 39638 21480
rect 44284 21468 44312 21576
rect 45278 21564 45284 21576
rect 45336 21564 45342 21616
rect 47946 21604 47952 21616
rect 47907 21576 47952 21604
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 44450 21536 44456 21548
rect 44363 21508 44456 21536
rect 44450 21496 44456 21508
rect 44508 21536 44514 21548
rect 45189 21539 45247 21545
rect 45189 21536 45201 21539
rect 44508 21508 45201 21536
rect 44508 21496 44514 21508
rect 45189 21505 45201 21508
rect 45235 21505 45247 21539
rect 45646 21536 45652 21548
rect 45607 21508 45652 21536
rect 45189 21499 45247 21505
rect 45646 21496 45652 21508
rect 45704 21496 45710 21548
rect 44361 21471 44419 21477
rect 44361 21468 44373 21471
rect 44284 21440 44373 21468
rect 44361 21437 44373 21440
rect 44407 21437 44419 21471
rect 44361 21431 44419 21437
rect 48133 21403 48191 21409
rect 48133 21400 48145 21403
rect 38672 21372 48145 21400
rect 48133 21369 48145 21372
rect 48179 21369 48191 21403
rect 48133 21363 48191 21369
rect 15212 21304 16068 21332
rect 14461 21295 14519 21301
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17092 21304 17417 21332
rect 17092 21292 17098 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 19521 21335 19579 21341
rect 19521 21301 19533 21335
rect 19567 21332 19579 21335
rect 20162 21332 20168 21344
rect 19567 21304 20168 21332
rect 19567 21301 19579 21304
rect 19521 21295 19579 21301
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 20625 21335 20683 21341
rect 20625 21332 20637 21335
rect 20496 21304 20637 21332
rect 20496 21292 20502 21304
rect 20625 21301 20637 21304
rect 20671 21301 20683 21335
rect 21174 21332 21180 21344
rect 21135 21304 21180 21332
rect 20625 21295 20683 21301
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 23569 21335 23627 21341
rect 23569 21332 23581 21335
rect 22888 21304 23581 21332
rect 22888 21292 22894 21304
rect 23569 21301 23581 21304
rect 23615 21301 23627 21335
rect 23569 21295 23627 21301
rect 25593 21335 25651 21341
rect 25593 21301 25605 21335
rect 25639 21332 25651 21335
rect 25774 21332 25780 21344
rect 25639 21304 25780 21332
rect 25639 21301 25651 21304
rect 25593 21295 25651 21301
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 46566 21292 46572 21344
rect 46624 21332 46630 21344
rect 46661 21335 46719 21341
rect 46661 21332 46673 21335
rect 46624 21304 46673 21332
rect 46624 21292 46630 21304
rect 46661 21301 46673 21304
rect 46707 21301 46719 21335
rect 46661 21295 46719 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9950 21088 9956 21140
rect 10008 21128 10014 21140
rect 10008 21100 28856 21128
rect 10008 21088 10014 21100
rect 10594 21020 10600 21072
rect 10652 21060 10658 21072
rect 11241 21063 11299 21069
rect 11241 21060 11253 21063
rect 10652 21032 11253 21060
rect 10652 21020 10658 21032
rect 11241 21029 11253 21032
rect 11287 21029 11299 21063
rect 11241 21023 11299 21029
rect 22373 21063 22431 21069
rect 22373 21029 22385 21063
rect 22419 21060 22431 21063
rect 22554 21060 22560 21072
rect 22419 21032 22560 21060
rect 22419 21029 22431 21032
rect 22373 21023 22431 21029
rect 22554 21020 22560 21032
rect 22612 21020 22618 21072
rect 8110 20992 8116 21004
rect 8071 20964 8116 20992
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20992 8447 20995
rect 9217 20995 9275 21001
rect 9217 20992 9229 20995
rect 8435 20964 9229 20992
rect 8435 20961 8447 20964
rect 8389 20955 8447 20961
rect 9217 20961 9229 20964
rect 9263 20961 9275 20995
rect 9217 20955 9275 20961
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14093 20995 14151 21001
rect 14093 20992 14105 20995
rect 13872 20964 14105 20992
rect 13872 20952 13878 20964
rect 14093 20961 14105 20964
rect 14139 20961 14151 20995
rect 14274 20992 14280 21004
rect 14235 20964 14280 20992
rect 14093 20955 14151 20961
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 15470 20992 15476 21004
rect 15431 20964 15476 20992
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 16482 20952 16488 21004
rect 16540 20992 16546 21004
rect 16853 20995 16911 21001
rect 16853 20992 16865 20995
rect 16540 20964 16865 20992
rect 16540 20952 16546 20964
rect 16853 20961 16865 20964
rect 16899 20961 16911 20995
rect 17034 20992 17040 21004
rect 16995 20964 17040 20992
rect 16853 20955 16911 20961
rect 17034 20952 17040 20964
rect 17092 20952 17098 21004
rect 20162 20992 20168 21004
rect 20123 20964 20168 20992
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 20438 20992 20444 21004
rect 20399 20964 20444 20992
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 25774 20992 25780 21004
rect 22060 20964 23152 20992
rect 25735 20964 25780 20992
rect 22060 20952 22066 20964
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7616 20896 8033 20924
rect 7616 20884 7622 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8938 20924 8944 20936
rect 8899 20896 8944 20924
rect 8021 20887 8079 20893
rect 8036 20788 8064 20887
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11974 20924 11980 20936
rect 11471 20896 11980 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19978 20924 19984 20936
rect 19291 20896 19984 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19978 20884 19984 20896
rect 20036 20884 20042 20936
rect 22646 20924 22652 20936
rect 22607 20896 22652 20924
rect 22646 20884 22652 20896
rect 22704 20884 22710 20936
rect 23124 20933 23152 20964
rect 25774 20952 25780 20964
rect 25832 20952 25838 21004
rect 27433 20995 27491 21001
rect 27433 20961 27445 20995
rect 27479 20992 27491 20995
rect 28718 20992 28724 21004
rect 27479 20964 28724 20992
rect 27479 20961 27491 20964
rect 27433 20955 27491 20961
rect 28718 20952 28724 20964
rect 28776 20952 28782 21004
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 23658 20884 23664 20936
rect 23716 20924 23722 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23716 20896 24409 20924
rect 23716 20884 23722 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25593 20927 25651 20933
rect 25593 20924 25605 20927
rect 24912 20896 25605 20924
rect 24912 20884 24918 20896
rect 25593 20893 25605 20896
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 27893 20927 27951 20933
rect 27893 20893 27905 20927
rect 27939 20893 27951 20927
rect 27893 20887 27951 20893
rect 9950 20816 9956 20868
rect 10008 20816 10014 20868
rect 18690 20856 18696 20868
rect 18651 20828 18696 20856
rect 18690 20816 18696 20828
rect 18748 20816 18754 20868
rect 21174 20816 21180 20868
rect 21232 20816 21238 20868
rect 22186 20816 22192 20868
rect 22244 20856 22250 20868
rect 22373 20859 22431 20865
rect 22373 20856 22385 20859
rect 22244 20828 22385 20856
rect 22244 20816 22250 20828
rect 22373 20825 22385 20828
rect 22419 20856 22431 20859
rect 25498 20856 25504 20868
rect 22419 20828 25504 20856
rect 22419 20825 22431 20828
rect 22373 20819 22431 20825
rect 25498 20816 25504 20828
rect 25556 20816 25562 20868
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 27522 20856 27528 20868
rect 26844 20828 27528 20856
rect 26844 20816 26850 20828
rect 27522 20816 27528 20828
rect 27580 20856 27586 20868
rect 27908 20856 27936 20887
rect 27580 20828 27936 20856
rect 27580 20816 27586 20828
rect 28626 20816 28632 20868
rect 28684 20856 28690 20868
rect 28721 20859 28779 20865
rect 28721 20856 28733 20859
rect 28684 20828 28733 20856
rect 28684 20816 28690 20828
rect 28721 20825 28733 20828
rect 28767 20825 28779 20859
rect 28828 20856 28856 21100
rect 45278 21088 45284 21140
rect 45336 21128 45342 21140
rect 45741 21131 45799 21137
rect 45741 21128 45753 21131
rect 45336 21100 45753 21128
rect 45336 21088 45342 21100
rect 45741 21097 45753 21100
rect 45787 21097 45799 21131
rect 45741 21091 45799 21097
rect 29549 20995 29607 21001
rect 29549 20961 29561 20995
rect 29595 20992 29607 20995
rect 30190 20992 30196 21004
rect 29595 20964 30196 20992
rect 29595 20961 29607 20964
rect 29549 20955 29607 20961
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 30466 20992 30472 21004
rect 30427 20964 30472 20992
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 45373 20927 45431 20933
rect 45373 20893 45385 20927
rect 45419 20924 45431 20927
rect 45462 20924 45468 20936
rect 45419 20896 45468 20924
rect 45419 20893 45431 20896
rect 45373 20887 45431 20893
rect 45462 20884 45468 20896
rect 45520 20884 45526 20936
rect 46290 20924 46296 20936
rect 46251 20896 46296 20924
rect 46290 20884 46296 20896
rect 46348 20884 46354 20936
rect 29733 20859 29791 20865
rect 29733 20856 29745 20859
rect 28828 20828 29745 20856
rect 28721 20819 28779 20825
rect 29733 20825 29745 20828
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 45557 20859 45615 20865
rect 45557 20825 45569 20859
rect 45603 20856 45615 20859
rect 45830 20856 45836 20868
rect 45603 20828 45836 20856
rect 45603 20825 45615 20828
rect 45557 20819 45615 20825
rect 10042 20788 10048 20800
rect 8036 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20788 10106 20800
rect 10689 20791 10747 20797
rect 10689 20788 10701 20791
rect 10100 20760 10701 20788
rect 10100 20748 10106 20760
rect 10689 20757 10701 20760
rect 10735 20757 10747 20791
rect 19334 20788 19340 20800
rect 19295 20760 19340 20788
rect 10689 20751 10747 20757
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 21913 20791 21971 20797
rect 21913 20788 21925 20791
rect 20312 20760 21925 20788
rect 20312 20748 20318 20760
rect 21913 20757 21925 20760
rect 21959 20788 21971 20791
rect 22557 20791 22615 20797
rect 22557 20788 22569 20791
rect 21959 20760 22569 20788
rect 21959 20757 21971 20760
rect 21913 20751 21971 20757
rect 22557 20757 22569 20760
rect 22603 20757 22615 20791
rect 22557 20751 22615 20757
rect 23198 20748 23204 20800
rect 23256 20788 23262 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 23256 20760 23305 20788
rect 23256 20748 23262 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 24486 20788 24492 20800
rect 24447 20760 24492 20788
rect 23293 20751 23351 20757
rect 24486 20748 24492 20760
rect 24544 20748 24550 20800
rect 28736 20788 28764 20819
rect 45830 20816 45836 20828
rect 45888 20816 45894 20868
rect 46477 20859 46535 20865
rect 46477 20825 46489 20859
rect 46523 20856 46535 20859
rect 47302 20856 47308 20868
rect 46523 20828 47308 20856
rect 46523 20825 46535 20828
rect 46477 20819 46535 20825
rect 47302 20816 47308 20828
rect 47360 20816 47366 20868
rect 32582 20788 32588 20800
rect 28736 20760 32588 20788
rect 32582 20748 32588 20760
rect 32640 20748 32646 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 25222 20584 25228 20596
rect 3568 20556 25228 20584
rect 3568 20544 3574 20556
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 25406 20544 25412 20596
rect 25464 20584 25470 20596
rect 33778 20584 33784 20596
rect 25464 20556 33784 20584
rect 25464 20544 25470 20556
rect 33778 20544 33784 20556
rect 33836 20544 33842 20596
rect 43717 20587 43775 20593
rect 43717 20553 43729 20587
rect 43763 20584 43775 20587
rect 44450 20584 44456 20596
rect 43763 20556 44456 20584
rect 43763 20553 43775 20556
rect 43717 20547 43775 20553
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 47670 20584 47676 20596
rect 44652 20556 45508 20584
rect 47631 20556 47676 20584
rect 3418 20476 3424 20528
rect 3476 20516 3482 20528
rect 9950 20516 9956 20528
rect 3476 20488 9674 20516
rect 9911 20488 9956 20516
rect 3476 20476 3482 20488
rect 7558 20448 7564 20460
rect 7519 20420 7564 20448
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20380 7803 20383
rect 7926 20380 7932 20392
rect 7791 20352 7932 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20349 8079 20383
rect 9646 20380 9674 20488
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 15010 20476 15016 20528
rect 15068 20516 15074 20528
rect 15657 20519 15715 20525
rect 15657 20516 15669 20519
rect 15068 20488 15669 20516
rect 15068 20476 15074 20488
rect 15657 20485 15669 20488
rect 15703 20485 15715 20519
rect 15657 20479 15715 20485
rect 18417 20519 18475 20525
rect 18417 20485 18429 20519
rect 18463 20516 18475 20519
rect 19334 20516 19340 20528
rect 18463 20488 19340 20516
rect 18463 20485 18475 20488
rect 18417 20479 18475 20485
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 24486 20476 24492 20528
rect 24544 20476 24550 20528
rect 27893 20519 27951 20525
rect 27893 20485 27905 20519
rect 27939 20516 27951 20519
rect 28810 20516 28816 20528
rect 27939 20488 28816 20516
rect 27939 20485 27951 20488
rect 27893 20479 27951 20485
rect 28810 20476 28816 20488
rect 28868 20476 28874 20528
rect 44652 20516 44680 20556
rect 45370 20516 45376 20528
rect 31864 20488 44680 20516
rect 45331 20488 45376 20516
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 10686 20448 10692 20460
rect 9916 20420 9961 20448
rect 10647 20420 10692 20448
rect 9916 20408 9922 20420
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 11790 20448 11796 20460
rect 11751 20420 11796 20448
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 12618 20448 12624 20460
rect 12579 20420 12624 20448
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 15335 20420 16865 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 16853 20417 16865 20420
rect 16899 20448 16911 20451
rect 17402 20448 17408 20460
rect 16899 20420 17408 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 18230 20448 18236 20460
rect 18191 20420 18236 20448
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 20036 20420 20545 20448
rect 20036 20408 20042 20420
rect 20533 20417 20545 20420
rect 20579 20448 20591 20451
rect 22554 20448 22560 20460
rect 20579 20420 22094 20448
rect 22515 20420 22560 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 12802 20380 12808 20392
rect 9646 20352 11008 20380
rect 12763 20352 12808 20380
rect 8021 20343 8079 20349
rect 4798 20204 4804 20256
rect 4856 20244 4862 20256
rect 8036 20244 8064 20343
rect 10505 20315 10563 20321
rect 10505 20281 10517 20315
rect 10551 20312 10563 20315
rect 10870 20312 10876 20324
rect 10551 20284 10876 20312
rect 10551 20281 10563 20284
rect 10505 20275 10563 20281
rect 10870 20272 10876 20284
rect 10928 20272 10934 20324
rect 10980 20312 11008 20352
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 14366 20380 14372 20392
rect 14327 20352 14372 20380
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 17034 20380 17040 20392
rect 16632 20352 17040 20380
rect 16632 20340 16638 20352
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20349 18751 20383
rect 22066 20380 22094 20420
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 22741 20451 22799 20457
rect 22741 20417 22753 20451
rect 22787 20448 22799 20451
rect 22830 20448 22836 20460
rect 22787 20420 22836 20448
rect 22787 20417 22799 20420
rect 22741 20411 22799 20417
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 23198 20448 23204 20460
rect 23159 20420 23204 20448
rect 23198 20408 23204 20420
rect 23256 20408 23262 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26786 20448 26792 20460
rect 26099 20420 26792 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26786 20408 26792 20420
rect 26844 20408 26850 20460
rect 27065 20451 27123 20457
rect 27065 20417 27077 20451
rect 27111 20448 27123 20451
rect 27246 20448 27252 20460
rect 27111 20420 27252 20448
rect 27111 20417 27123 20420
rect 27065 20411 27123 20417
rect 27246 20408 27252 20420
rect 27304 20408 27310 20460
rect 22649 20383 22707 20389
rect 22066 20352 22600 20380
rect 18693 20343 18751 20349
rect 18708 20312 18736 20343
rect 10980 20284 18736 20312
rect 18892 20284 20760 20312
rect 11974 20244 11980 20256
rect 4856 20216 8064 20244
rect 11935 20216 11980 20244
rect 4856 20204 4862 20216
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 16666 20204 16672 20256
rect 16724 20244 16730 20256
rect 16942 20244 16948 20256
rect 16724 20216 16948 20244
rect 16724 20204 16730 20216
rect 16942 20204 16948 20216
rect 17000 20244 17006 20256
rect 18892 20244 18920 20284
rect 17000 20216 18920 20244
rect 17000 20204 17006 20216
rect 19702 20204 19708 20256
rect 19760 20244 19766 20256
rect 20625 20247 20683 20253
rect 20625 20244 20637 20247
rect 19760 20216 20637 20244
rect 19760 20204 19766 20216
rect 20625 20213 20637 20216
rect 20671 20213 20683 20247
rect 20732 20244 20760 20284
rect 22462 20244 22468 20256
rect 20732 20216 22468 20244
rect 20625 20207 20683 20213
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 22572 20244 22600 20352
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 23477 20383 23535 20389
rect 23477 20380 23489 20383
rect 22695 20352 23489 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 23477 20349 23489 20352
rect 23523 20349 23535 20383
rect 23477 20343 23535 20349
rect 24949 20383 25007 20389
rect 24949 20349 24961 20383
rect 24995 20380 25007 20383
rect 25498 20380 25504 20392
rect 24995 20352 25504 20380
rect 24995 20349 25007 20352
rect 24949 20343 25007 20349
rect 25498 20340 25504 20352
rect 25556 20340 25562 20392
rect 27706 20380 27712 20392
rect 27667 20352 27712 20380
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 28169 20383 28227 20389
rect 28169 20349 28181 20383
rect 28215 20349 28227 20383
rect 28169 20343 28227 20349
rect 25222 20272 25228 20324
rect 25280 20312 25286 20324
rect 28184 20312 28212 20343
rect 25280 20284 28212 20312
rect 25280 20272 25286 20284
rect 25130 20244 25136 20256
rect 22572 20216 25136 20244
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 26142 20244 26148 20256
rect 26103 20216 26148 20244
rect 26142 20204 26148 20216
rect 26200 20204 26206 20256
rect 26786 20204 26792 20256
rect 26844 20244 26850 20256
rect 27157 20247 27215 20253
rect 27157 20244 27169 20247
rect 26844 20216 27169 20244
rect 26844 20204 26850 20216
rect 27157 20213 27169 20216
rect 27203 20213 27215 20247
rect 27157 20207 27215 20213
rect 27246 20204 27252 20256
rect 27304 20244 27310 20256
rect 31864 20244 31892 20488
rect 45370 20476 45376 20488
rect 45428 20476 45434 20528
rect 45480 20516 45508 20556
rect 47670 20544 47676 20556
rect 47728 20544 47734 20596
rect 47854 20516 47860 20528
rect 45480 20488 47860 20516
rect 47854 20476 47860 20488
rect 47912 20476 47918 20528
rect 43806 20448 43812 20460
rect 43767 20420 43812 20448
rect 43806 20408 43812 20420
rect 43864 20408 43870 20460
rect 44174 20448 44180 20460
rect 44135 20420 44180 20448
rect 44174 20408 44180 20420
rect 44232 20408 44238 20460
rect 45094 20408 45100 20460
rect 45152 20438 45158 20460
rect 47578 20448 47584 20460
rect 45152 20423 45232 20438
rect 45152 20417 45247 20423
rect 47539 20420 47584 20448
rect 45152 20410 45201 20417
rect 45152 20408 45158 20410
rect 33778 20340 33784 20392
rect 33836 20380 33842 20392
rect 44450 20380 44456 20392
rect 33836 20352 44456 20380
rect 33836 20340 33842 20352
rect 44450 20340 44456 20352
rect 44508 20340 44514 20392
rect 44634 20380 44640 20392
rect 44595 20352 44640 20380
rect 44634 20340 44640 20352
rect 44692 20340 44698 20392
rect 45189 20383 45201 20410
rect 45235 20383 45247 20417
rect 47578 20408 47584 20420
rect 47636 20408 47642 20460
rect 45189 20377 45247 20383
rect 46658 20380 46664 20392
rect 46619 20352 46664 20380
rect 46658 20340 46664 20352
rect 46716 20340 46722 20392
rect 40770 20272 40776 20324
rect 40828 20312 40834 20324
rect 44266 20312 44272 20324
rect 40828 20284 44272 20312
rect 40828 20272 40834 20284
rect 44266 20272 44272 20284
rect 44324 20272 44330 20324
rect 44358 20272 44364 20324
rect 44416 20312 44422 20324
rect 45370 20312 45376 20324
rect 44416 20284 45376 20312
rect 44416 20272 44422 20284
rect 45370 20272 45376 20284
rect 45428 20272 45434 20324
rect 27304 20216 31892 20244
rect 27304 20204 27310 20216
rect 40678 20204 40684 20256
rect 40736 20244 40742 20256
rect 46014 20244 46020 20256
rect 40736 20216 46020 20244
rect 40736 20204 40742 20216
rect 46014 20204 46020 20216
rect 46072 20204 46078 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 7926 20040 7932 20052
rect 7887 20012 7932 20040
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 8938 20040 8944 20052
rect 8899 20012 8944 20040
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 28534 20040 28540 20052
rect 16500 20012 28540 20040
rect 3786 19932 3792 19984
rect 3844 19972 3850 19984
rect 16500 19972 16528 20012
rect 28534 20000 28540 20012
rect 28592 20000 28598 20052
rect 44266 20000 44272 20052
rect 44324 20040 44330 20052
rect 47578 20040 47584 20052
rect 44324 20012 47584 20040
rect 44324 20000 44330 20012
rect 47578 20000 47584 20012
rect 47636 20000 47642 20052
rect 3844 19944 16528 19972
rect 3844 19932 3850 19944
rect 18230 19932 18236 19984
rect 18288 19972 18294 19984
rect 19426 19972 19432 19984
rect 18288 19944 19432 19972
rect 18288 19932 18294 19944
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 20254 19972 20260 19984
rect 19536 19944 20260 19972
rect 7852 19876 12756 19904
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 7852 19845 7880 19876
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 7837 19839 7895 19845
rect 7837 19805 7849 19839
rect 7883 19805 7895 19839
rect 9122 19836 9128 19848
rect 9083 19808 9128 19836
rect 7837 19799 7895 19805
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 12728 19845 12756 19876
rect 13722 19864 13728 19916
rect 13780 19904 13786 19916
rect 16390 19904 16396 19916
rect 13780 19876 16252 19904
rect 16351 19876 16396 19904
rect 13780 19864 13786 19876
rect 12713 19839 12771 19845
rect 12713 19805 12725 19839
rect 12759 19836 12771 19839
rect 15010 19836 15016 19848
rect 12759 19808 15016 19836
rect 12759 19805 12771 19808
rect 12713 19799 12771 19805
rect 15010 19796 15016 19808
rect 15068 19796 15074 19848
rect 15194 19836 15200 19848
rect 15155 19808 15200 19836
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 15381 19703 15439 19709
rect 15381 19669 15393 19703
rect 15427 19700 15439 19703
rect 16132 19700 16160 19799
rect 16224 19768 16252 19876
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 19536 19913 19564 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 22462 19932 22468 19984
rect 22520 19972 22526 19984
rect 25130 19972 25136 19984
rect 22520 19944 24992 19972
rect 25091 19944 25136 19972
rect 22520 19932 22526 19944
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19873 19579 19907
rect 19702 19904 19708 19916
rect 19663 19876 19708 19904
rect 19521 19867 19579 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 22646 19904 22652 19916
rect 20916 19876 22652 19904
rect 17402 19836 17408 19848
rect 17363 19808 17408 19836
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17512 19808 18368 19836
rect 17512 19768 17540 19808
rect 18230 19768 18236 19780
rect 16224 19740 17540 19768
rect 18191 19740 18236 19768
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 18340 19768 18368 19808
rect 20916 19768 20944 19876
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 22925 19907 22983 19913
rect 22925 19873 22937 19907
rect 22971 19904 22983 19907
rect 23014 19904 23020 19916
rect 22971 19876 23020 19904
rect 22971 19873 22983 19876
rect 22925 19867 22983 19873
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 23201 19907 23259 19913
rect 23201 19873 23213 19907
rect 23247 19904 23259 19907
rect 23382 19904 23388 19916
rect 23247 19876 23388 19904
rect 23247 19873 23259 19876
rect 23201 19867 23259 19873
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 24964 19904 24992 19944
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 26510 19932 26516 19984
rect 26568 19972 26574 19984
rect 44634 19972 44640 19984
rect 26568 19944 31754 19972
rect 26568 19932 26574 19944
rect 27982 19904 27988 19916
rect 24964 19876 27988 19904
rect 27982 19864 27988 19876
rect 28040 19864 28046 19916
rect 31726 19904 31754 19944
rect 43732 19944 44640 19972
rect 40773 19907 40831 19913
rect 31726 19876 35894 19904
rect 22002 19836 22008 19848
rect 21963 19808 22008 19836
rect 22002 19796 22008 19808
rect 22060 19796 22066 19848
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19838 22891 19839
rect 22879 19810 22968 19838
rect 23658 19836 23664 19848
rect 22879 19805 22891 19810
rect 22833 19799 22891 19805
rect 21358 19768 21364 19780
rect 18340 19740 20944 19768
rect 21319 19740 21364 19768
rect 21358 19728 21364 19740
rect 21416 19728 21422 19780
rect 22940 19768 22968 19810
rect 23619 19808 23664 19836
rect 23658 19796 23664 19808
rect 23716 19836 23722 19848
rect 24302 19836 24308 19848
rect 23716 19808 24308 19836
rect 23716 19796 23722 19808
rect 24302 19796 24308 19808
rect 24360 19796 24366 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25774 19836 25780 19848
rect 24995 19808 25780 19836
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25774 19796 25780 19808
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19836 25927 19839
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 25915 19808 27169 19836
rect 25915 19805 25927 19808
rect 25869 19799 25927 19805
rect 27157 19805 27169 19808
rect 27203 19805 27215 19839
rect 27157 19799 27215 19805
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 28629 19839 28687 19845
rect 28629 19836 28641 19839
rect 27304 19808 28641 19836
rect 27304 19796 27310 19808
rect 28629 19805 28641 19808
rect 28675 19805 28687 19839
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 28629 19799 28687 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 28920 19808 31754 19836
rect 23290 19768 23296 19780
rect 22940 19740 23296 19768
rect 23290 19728 23296 19740
rect 23348 19768 23354 19780
rect 24854 19768 24860 19780
rect 23348 19740 24860 19768
rect 23348 19728 23354 19740
rect 24854 19728 24860 19740
rect 24912 19728 24918 19780
rect 26510 19768 26516 19780
rect 26471 19740 26516 19768
rect 26510 19728 26516 19740
rect 26568 19728 26574 19780
rect 27798 19728 27804 19780
rect 27856 19768 27862 19780
rect 27985 19771 28043 19777
rect 27985 19768 27997 19771
rect 27856 19740 27997 19768
rect 27856 19728 27862 19740
rect 27985 19737 27997 19740
rect 28031 19768 28043 19771
rect 28920 19768 28948 19808
rect 28031 19740 28948 19768
rect 28997 19771 29055 19777
rect 28031 19737 28043 19740
rect 27985 19731 28043 19737
rect 28997 19737 29009 19771
rect 29043 19768 29055 19771
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 29043 19740 30021 19768
rect 29043 19737 29055 19740
rect 28997 19731 29055 19737
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 30009 19731 30067 19737
rect 17402 19700 17408 19712
rect 15427 19672 17408 19700
rect 15427 19669 15439 19672
rect 15381 19663 15439 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 19426 19700 19432 19712
rect 18196 19672 19432 19700
rect 18196 19660 18202 19672
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 22097 19703 22155 19709
rect 22097 19669 22109 19703
rect 22143 19700 22155 19703
rect 23106 19700 23112 19712
rect 22143 19672 23112 19700
rect 22143 19669 22155 19672
rect 22097 19663 22155 19669
rect 23106 19660 23112 19672
rect 23164 19660 23170 19712
rect 23753 19703 23811 19709
rect 23753 19669 23765 19703
rect 23799 19700 23811 19703
rect 23842 19700 23848 19712
rect 23799 19672 23848 19700
rect 23799 19669 23811 19672
rect 23753 19663 23811 19669
rect 23842 19660 23848 19672
rect 23900 19660 23906 19712
rect 23934 19660 23940 19712
rect 23992 19700 23998 19712
rect 26528 19700 26556 19728
rect 23992 19672 26556 19700
rect 23992 19660 23998 19672
rect 27706 19660 27712 19712
rect 27764 19700 27770 19712
rect 28902 19700 28908 19712
rect 27764 19672 28908 19700
rect 27764 19660 27770 19672
rect 28902 19660 28908 19672
rect 28960 19700 28966 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 28960 19672 30113 19700
rect 28960 19660 28966 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 31726 19700 31754 19808
rect 35866 19768 35894 19876
rect 40773 19873 40785 19907
rect 40819 19904 40831 19907
rect 43625 19907 43683 19913
rect 40819 19876 43484 19904
rect 40819 19873 40831 19876
rect 40773 19867 40831 19873
rect 40678 19768 40684 19780
rect 35866 19740 40684 19768
rect 40678 19728 40684 19740
rect 40736 19728 40742 19780
rect 40954 19768 40960 19780
rect 40915 19740 40960 19768
rect 40954 19728 40960 19740
rect 41012 19728 41018 19780
rect 42610 19768 42616 19780
rect 42571 19740 42616 19768
rect 42610 19728 42616 19740
rect 42668 19728 42674 19780
rect 43456 19768 43484 19876
rect 43625 19873 43637 19907
rect 43671 19904 43683 19907
rect 43732 19904 43760 19944
rect 44634 19932 44640 19944
rect 44692 19932 44698 19984
rect 45370 19972 45376 19984
rect 45331 19944 45376 19972
rect 45370 19932 45376 19944
rect 45428 19932 45434 19984
rect 45465 19907 45523 19913
rect 45465 19904 45477 19907
rect 43671 19876 43760 19904
rect 43824 19876 45477 19904
rect 43671 19873 43683 19876
rect 43625 19867 43683 19873
rect 43824 19845 43852 19876
rect 45465 19873 45477 19876
rect 45511 19873 45523 19907
rect 45465 19867 45523 19873
rect 46477 19907 46535 19913
rect 46477 19873 46489 19907
rect 46523 19904 46535 19907
rect 48038 19904 48044 19916
rect 46523 19876 48044 19904
rect 46523 19873 46535 19876
rect 46477 19867 46535 19873
rect 48038 19864 48044 19876
rect 48096 19864 48102 19916
rect 43809 19839 43867 19845
rect 43809 19805 43821 19839
rect 43855 19805 43867 19839
rect 43809 19799 43867 19805
rect 43990 19796 43996 19848
rect 44048 19836 44054 19848
rect 46293 19839 46351 19845
rect 46293 19836 46305 19839
rect 44048 19808 46305 19836
rect 44048 19796 44054 19808
rect 46293 19805 46305 19808
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 43456 19740 43576 19768
rect 43438 19700 43444 19712
rect 31726 19672 43444 19700
rect 30101 19663 30159 19669
rect 43438 19660 43444 19672
rect 43496 19660 43502 19712
rect 43548 19700 43576 19740
rect 43898 19728 43904 19780
rect 43956 19768 43962 19780
rect 45005 19771 45063 19777
rect 45005 19768 45017 19771
rect 43956 19740 45017 19768
rect 43956 19728 43962 19740
rect 45005 19737 45017 19740
rect 45051 19737 45063 19771
rect 45005 19731 45063 19737
rect 46658 19728 46664 19780
rect 46716 19768 46722 19780
rect 48133 19771 48191 19777
rect 48133 19768 48145 19771
rect 46716 19740 48145 19768
rect 46716 19728 46722 19740
rect 48133 19737 48145 19740
rect 48179 19737 48191 19771
rect 48133 19731 48191 19737
rect 44453 19703 44511 19709
rect 44453 19700 44465 19703
rect 43548 19672 44465 19700
rect 44453 19669 44465 19672
rect 44499 19700 44511 19703
rect 45094 19700 45100 19712
rect 44499 19672 45100 19700
rect 44499 19669 44511 19672
rect 44453 19663 44511 19669
rect 45094 19660 45100 19672
rect 45152 19660 45158 19712
rect 45554 19660 45560 19712
rect 45612 19700 45618 19712
rect 47026 19700 47032 19712
rect 45612 19672 47032 19700
rect 45612 19660 45618 19672
rect 47026 19660 47032 19672
rect 47084 19660 47090 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 23014 19496 23020 19508
rect 15252 19468 23020 19496
rect 15252 19456 15258 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 26142 19496 26148 19508
rect 23216 19468 26148 19496
rect 8205 19431 8263 19437
rect 8205 19397 8217 19431
rect 8251 19428 8263 19431
rect 8294 19428 8300 19440
rect 8251 19400 8300 19428
rect 8251 19397 8263 19400
rect 8205 19391 8263 19397
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 14369 19431 14427 19437
rect 14369 19397 14381 19431
rect 14415 19428 14427 19431
rect 16761 19431 16819 19437
rect 16761 19428 16773 19431
rect 14415 19400 16773 19428
rect 14415 19397 14427 19400
rect 14369 19391 14427 19397
rect 16761 19397 16773 19400
rect 16807 19397 16819 19431
rect 18506 19428 18512 19440
rect 16761 19391 16819 19397
rect 17420 19400 18512 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 8036 19292 8064 19323
rect 8386 19292 8392 19304
rect 8036 19264 8392 19292
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 8478 19224 8484 19236
rect 3108 19196 8484 19224
rect 3108 19184 3114 19196
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 14 19116 20 19168
rect 72 19156 78 19168
rect 8588 19156 8616 19255
rect 9122 19252 9128 19304
rect 9180 19292 9186 19304
rect 11900 19292 11928 19323
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 12860 19332 13185 19360
rect 12860 19320 12866 19332
rect 13173 19329 13185 19332
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 14185 19363 14243 19369
rect 14185 19360 14197 19363
rect 13504 19332 14197 19360
rect 13504 19320 13510 19332
rect 14185 19329 14197 19332
rect 14231 19329 14243 19363
rect 16666 19360 16672 19372
rect 16627 19332 16672 19360
rect 14185 19323 14243 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17420 19369 17448 19400
rect 18506 19388 18512 19400
rect 18564 19388 18570 19440
rect 19150 19388 19156 19440
rect 19208 19428 19214 19440
rect 19245 19431 19303 19437
rect 19245 19428 19257 19431
rect 19208 19400 19257 19428
rect 19208 19388 19214 19400
rect 19245 19397 19257 19400
rect 19291 19397 19303 19431
rect 19245 19391 19303 19397
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 23216 19428 23244 19468
rect 26142 19456 26148 19468
rect 26200 19456 26206 19508
rect 40865 19499 40923 19505
rect 40865 19465 40877 19499
rect 40911 19496 40923 19499
rect 40954 19496 40960 19508
rect 40911 19468 40960 19496
rect 40911 19465 40923 19468
rect 40865 19459 40923 19465
rect 40954 19456 40960 19468
rect 41012 19456 41018 19508
rect 43806 19456 43812 19508
rect 43864 19496 43870 19508
rect 43993 19499 44051 19505
rect 43993 19496 44005 19499
rect 43864 19468 44005 19496
rect 43864 19456 43870 19468
rect 43993 19465 44005 19468
rect 44039 19465 44051 19499
rect 43993 19459 44051 19465
rect 44836 19468 45324 19496
rect 23382 19428 23388 19440
rect 19484 19400 23244 19428
rect 23343 19400 23388 19428
rect 19484 19388 19490 19400
rect 23382 19388 23388 19400
rect 23440 19388 23446 19440
rect 23842 19388 23848 19440
rect 23900 19388 23906 19440
rect 27154 19428 27160 19440
rect 27115 19400 27160 19428
rect 27154 19388 27160 19400
rect 27212 19388 27218 19440
rect 27341 19431 27399 19437
rect 27341 19397 27353 19431
rect 27387 19428 27399 19431
rect 27430 19428 27436 19440
rect 27387 19400 27436 19428
rect 27387 19397 27399 19400
rect 27341 19391 27399 19397
rect 27430 19388 27436 19400
rect 27488 19388 27494 19440
rect 30282 19388 30288 19440
rect 30340 19428 30346 19440
rect 44836 19428 44864 19468
rect 30340 19400 30972 19428
rect 30340 19388 30346 19400
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19392 19332 19717 19360
rect 19392 19320 19398 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 21818 19320 21824 19372
rect 21876 19360 21882 19372
rect 21913 19363 21971 19369
rect 21913 19360 21925 19363
rect 21876 19332 21925 19360
rect 21876 19320 21882 19332
rect 21913 19329 21925 19332
rect 21959 19329 21971 19363
rect 23106 19360 23112 19372
rect 23067 19332 23112 19360
rect 21913 19323 21971 19329
rect 23106 19320 23112 19332
rect 23164 19320 23170 19372
rect 25774 19360 25780 19372
rect 25735 19332 25780 19360
rect 25774 19320 25780 19332
rect 25832 19320 25838 19372
rect 25866 19320 25872 19372
rect 25924 19360 25930 19372
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 25924 19332 26157 19360
rect 25924 19320 25930 19332
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 28350 19360 28356 19372
rect 28311 19332 28356 19360
rect 26145 19323 26203 19329
rect 28350 19320 28356 19332
rect 28408 19320 28414 19372
rect 28534 19360 28540 19372
rect 28495 19332 28540 19360
rect 28534 19320 28540 19332
rect 28592 19320 28598 19372
rect 29641 19363 29699 19369
rect 29641 19329 29653 19363
rect 29687 19360 29699 19363
rect 29822 19360 29828 19372
rect 29687 19332 29828 19360
rect 29687 19329 29699 19332
rect 29641 19323 29699 19329
rect 29822 19320 29828 19332
rect 29880 19360 29886 19372
rect 30944 19369 30972 19400
rect 43916 19400 44864 19428
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 29880 19332 30757 19360
rect 29880 19320 29886 19332
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19329 30987 19363
rect 30929 19323 30987 19329
rect 31297 19363 31355 19369
rect 31297 19329 31309 19363
rect 31343 19329 31355 19363
rect 31297 19323 31355 19329
rect 11974 19292 11980 19304
rect 9180 19264 11980 19292
rect 9180 19252 9186 19264
rect 11974 19252 11980 19264
rect 12032 19292 12038 19304
rect 13538 19292 13544 19304
rect 12032 19264 13544 19292
rect 12032 19252 12038 19264
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 13780 19264 14657 19292
rect 13780 19252 13786 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 17586 19292 17592 19304
rect 17547 19264 17592 19292
rect 14645 19255 14703 19261
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 27525 19295 27583 19301
rect 22066 19264 26280 19292
rect 8662 19184 8668 19236
rect 8720 19224 8726 19236
rect 22066 19224 22094 19264
rect 24854 19224 24860 19236
rect 8720 19196 22094 19224
rect 24815 19196 24860 19224
rect 8720 19184 8726 19196
rect 24854 19184 24860 19196
rect 24912 19184 24918 19236
rect 26252 19224 26280 19264
rect 27525 19261 27537 19295
rect 27571 19292 27583 19295
rect 28810 19292 28816 19304
rect 27571 19264 28816 19292
rect 27571 19261 27583 19264
rect 27525 19255 27583 19261
rect 28810 19252 28816 19264
rect 28868 19252 28874 19304
rect 29730 19292 29736 19304
rect 29691 19264 29736 19292
rect 29730 19252 29736 19264
rect 29788 19252 29794 19304
rect 30190 19292 30196 19304
rect 30151 19264 30196 19292
rect 30190 19252 30196 19264
rect 30248 19252 30254 19304
rect 31312 19292 31340 19323
rect 31386 19320 31392 19372
rect 31444 19360 31450 19372
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31444 19332 32137 19360
rect 31444 19320 31450 19332
rect 32125 19329 32137 19332
rect 32171 19360 32183 19363
rect 40770 19360 40776 19372
rect 32171 19332 40776 19360
rect 32171 19329 32183 19332
rect 32125 19323 32183 19329
rect 40770 19320 40776 19332
rect 40828 19320 40834 19372
rect 42978 19320 42984 19372
rect 43036 19360 43042 19372
rect 43916 19369 43944 19400
rect 44910 19388 44916 19440
rect 44968 19388 44974 19440
rect 45296 19428 45324 19468
rect 45370 19456 45376 19508
rect 45428 19496 45434 19508
rect 46201 19499 46259 19505
rect 46201 19496 46213 19499
rect 45428 19468 46213 19496
rect 45428 19456 45434 19468
rect 46201 19465 46213 19468
rect 46247 19465 46259 19499
rect 46201 19459 46259 19465
rect 47302 19456 47308 19508
rect 47360 19496 47366 19508
rect 47673 19499 47731 19505
rect 47673 19496 47685 19499
rect 47360 19468 47685 19496
rect 47360 19456 47366 19468
rect 47673 19465 47685 19468
rect 47719 19465 47731 19499
rect 47673 19459 47731 19465
rect 45296 19400 46152 19428
rect 43901 19363 43959 19369
rect 43901 19360 43913 19363
rect 43036 19332 43913 19360
rect 43036 19320 43042 19332
rect 43901 19329 43913 19332
rect 43947 19329 43959 19363
rect 43901 19323 43959 19329
rect 44085 19363 44143 19369
rect 44085 19329 44097 19363
rect 44131 19360 44143 19363
rect 44821 19363 44879 19369
rect 44131 19332 44772 19360
rect 44131 19329 44143 19332
rect 44085 19323 44143 19329
rect 30392 19264 31340 19292
rect 44744 19292 44772 19332
rect 44821 19329 44833 19363
rect 44867 19358 44879 19363
rect 44928 19358 44956 19388
rect 46124 19369 46152 19400
rect 47026 19388 47032 19440
rect 47084 19428 47090 19440
rect 47084 19400 47624 19428
rect 47084 19388 47090 19400
rect 46109 19363 46167 19369
rect 44867 19330 44956 19358
rect 45020 19332 46060 19360
rect 44867 19329 44879 19330
rect 44821 19323 44879 19329
rect 45020 19292 45048 19332
rect 44744 19264 45048 19292
rect 30392 19236 30420 19264
rect 45094 19252 45100 19304
rect 45152 19292 45158 19304
rect 45649 19295 45707 19301
rect 45152 19264 45197 19292
rect 45152 19252 45158 19264
rect 45649 19261 45661 19295
rect 45695 19292 45707 19295
rect 45738 19292 45744 19304
rect 45695 19264 45744 19292
rect 45695 19261 45707 19264
rect 45649 19255 45707 19261
rect 45738 19252 45744 19264
rect 45796 19252 45802 19304
rect 46032 19292 46060 19332
rect 46109 19329 46121 19363
rect 46155 19329 46167 19363
rect 46293 19363 46351 19369
rect 46293 19360 46305 19363
rect 46109 19323 46167 19329
rect 46216 19332 46305 19360
rect 46216 19292 46244 19332
rect 46293 19329 46305 19332
rect 46339 19360 46351 19363
rect 46382 19360 46388 19372
rect 46339 19332 46388 19360
rect 46339 19329 46351 19332
rect 46293 19323 46351 19329
rect 46382 19320 46388 19332
rect 46440 19360 46446 19372
rect 46750 19360 46756 19372
rect 46440 19332 46756 19360
rect 46440 19320 46446 19332
rect 46750 19320 46756 19332
rect 46808 19320 46814 19372
rect 47596 19369 47624 19400
rect 47581 19363 47639 19369
rect 47581 19329 47593 19363
rect 47627 19329 47639 19363
rect 47581 19323 47639 19329
rect 46032 19264 46244 19292
rect 27890 19224 27896 19236
rect 26252 19196 27896 19224
rect 27890 19184 27896 19196
rect 27948 19184 27954 19236
rect 28445 19227 28503 19233
rect 28445 19193 28457 19227
rect 28491 19224 28503 19227
rect 30374 19224 30380 19236
rect 28491 19196 30380 19224
rect 28491 19193 28503 19196
rect 28445 19187 28503 19193
rect 30374 19184 30380 19196
rect 30432 19184 30438 19236
rect 43438 19184 43444 19236
rect 43496 19224 43502 19236
rect 46106 19224 46112 19236
rect 43496 19196 46112 19224
rect 43496 19184 43502 19196
rect 46106 19184 46112 19196
rect 46164 19184 46170 19236
rect 46290 19184 46296 19236
rect 46348 19224 46354 19236
rect 47029 19227 47087 19233
rect 47029 19224 47041 19227
rect 46348 19196 47041 19224
rect 46348 19184 46354 19196
rect 47029 19193 47041 19196
rect 47075 19193 47087 19227
rect 47029 19187 47087 19193
rect 72 19128 8616 19156
rect 72 19116 78 19128
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 11238 19156 11244 19168
rect 9824 19128 11244 19156
rect 9824 19116 9830 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 11790 19156 11796 19168
rect 11747 19128 11796 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 12802 19156 12808 19168
rect 12667 19128 12808 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13170 19116 13176 19168
rect 13228 19156 13234 19168
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 13228 19128 13277 19156
rect 13228 19116 13234 19128
rect 13265 19125 13277 19128
rect 13311 19125 13323 19159
rect 13265 19119 13323 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 18230 19156 18236 19168
rect 13412 19128 18236 19156
rect 13412 19116 13418 19128
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20254 19156 20260 19168
rect 19935 19128 20260 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21968 19128 22017 19156
rect 21968 19116 21974 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 29546 19156 29552 19168
rect 22704 19128 29552 19156
rect 22704 19116 22710 19128
rect 29546 19116 29552 19128
rect 29604 19116 29610 19168
rect 31202 19156 31208 19168
rect 31163 19128 31208 19156
rect 31202 19116 31208 19128
rect 31260 19116 31266 19168
rect 32217 19159 32275 19165
rect 32217 19125 32229 19159
rect 32263 19156 32275 19159
rect 32306 19156 32312 19168
rect 32263 19128 32312 19156
rect 32263 19125 32275 19128
rect 32217 19119 32275 19125
rect 32306 19116 32312 19128
rect 32364 19116 32370 19168
rect 33502 19116 33508 19168
rect 33560 19156 33566 19168
rect 43806 19156 43812 19168
rect 33560 19128 43812 19156
rect 33560 19116 33566 19128
rect 43806 19116 43812 19128
rect 43864 19116 43870 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 2225 18915 2283 18921
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 16298 18952 16304 18964
rect 9232 18924 16304 18952
rect 2038 18844 2044 18896
rect 2096 18884 2102 18896
rect 9232 18884 9260 18924
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 30466 18952 30472 18964
rect 16632 18924 30472 18952
rect 16632 18912 16638 18924
rect 30466 18912 30472 18924
rect 30524 18912 30530 18964
rect 32122 18912 32128 18964
rect 32180 18952 32186 18964
rect 33321 18955 33379 18961
rect 33321 18952 33333 18955
rect 32180 18924 33333 18952
rect 32180 18912 32186 18924
rect 33321 18921 33333 18924
rect 33367 18952 33379 18955
rect 43990 18952 43996 18964
rect 33367 18924 43996 18952
rect 33367 18921 33379 18924
rect 33321 18915 33379 18921
rect 43990 18912 43996 18924
rect 44048 18912 44054 18964
rect 44269 18955 44327 18961
rect 44269 18921 44281 18955
rect 44315 18952 44327 18955
rect 45094 18952 45100 18964
rect 44315 18924 45100 18952
rect 44315 18921 44327 18924
rect 44269 18915 44327 18921
rect 45094 18912 45100 18924
rect 45152 18912 45158 18964
rect 18322 18884 18328 18896
rect 2096 18856 9260 18884
rect 10428 18856 11928 18884
rect 2096 18844 2102 18856
rect 10428 18816 10456 18856
rect 11790 18816 11796 18828
rect 6886 18788 10456 18816
rect 11751 18788 11796 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 6886 18748 6914 18788
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 11900 18816 11928 18856
rect 14384 18856 15332 18884
rect 18283 18856 18328 18884
rect 14384 18816 14412 18856
rect 15194 18816 15200 18828
rect 11900 18788 14412 18816
rect 14476 18788 15200 18816
rect 2188 18720 6914 18748
rect 2188 18708 2194 18720
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 8168 18720 8217 18748
rect 8168 18708 8174 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 9030 18708 9036 18760
rect 9088 18748 9094 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 9088 18720 9137 18748
rect 9088 18708 9094 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 13170 18708 13176 18760
rect 13228 18708 13234 18760
rect 14476 18757 14504 18788
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 15304 18816 15332 18856
rect 18322 18844 18328 18856
rect 18380 18844 18386 18896
rect 18414 18844 18420 18896
rect 18472 18884 18478 18896
rect 19150 18884 19156 18896
rect 18472 18856 19156 18884
rect 18472 18844 18478 18856
rect 19150 18844 19156 18856
rect 19208 18884 19214 18896
rect 22646 18884 22652 18896
rect 19208 18856 22652 18884
rect 19208 18844 19214 18856
rect 16482 18816 16488 18828
rect 15304 18788 16488 18816
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 19260 18825 19288 18856
rect 22646 18844 22652 18856
rect 22704 18844 22710 18896
rect 23014 18844 23020 18896
rect 23072 18884 23078 18896
rect 31113 18887 31171 18893
rect 23072 18856 25084 18884
rect 23072 18844 23078 18856
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18816 19303 18819
rect 19429 18819 19487 18825
rect 19291 18788 19325 18816
rect 19291 18785 19303 18788
rect 19245 18779 19303 18785
rect 19429 18785 19441 18819
rect 19475 18816 19487 18819
rect 20070 18816 20076 18828
rect 19475 18788 20076 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 21910 18816 21916 18828
rect 21871 18788 21916 18816
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 22278 18816 22284 18828
rect 22239 18788 22284 18816
rect 22278 18776 22284 18788
rect 22336 18776 22342 18828
rect 25056 18816 25084 18856
rect 31113 18853 31125 18887
rect 31159 18884 31171 18887
rect 33502 18884 33508 18896
rect 31159 18856 33508 18884
rect 31159 18853 31171 18856
rect 31113 18847 31171 18853
rect 33502 18844 33508 18856
rect 33560 18844 33566 18896
rect 43257 18887 43315 18893
rect 43257 18853 43269 18887
rect 43303 18853 43315 18887
rect 43257 18847 43315 18853
rect 27062 18816 27068 18828
rect 25056 18788 27068 18816
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14461 18711 14519 18717
rect 14660 18720 15301 18748
rect 9398 18680 9404 18692
rect 9359 18652 9404 18680
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 10778 18680 10784 18692
rect 10626 18652 10784 18680
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 12069 18683 12127 18689
rect 12069 18649 12081 18683
rect 12115 18649 12127 18683
rect 12069 18643 12127 18649
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 10226 18612 10232 18624
rect 8444 18584 10232 18612
rect 8444 18572 8450 18584
rect 10226 18572 10232 18584
rect 10284 18612 10290 18624
rect 10870 18612 10876 18624
rect 10284 18584 10876 18612
rect 10284 18572 10290 18584
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 12084 18612 12112 18643
rect 14660 18624 14688 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 16574 18748 16580 18760
rect 16535 18720 16580 18748
rect 15289 18711 15347 18717
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 25056 18757 25084 18788
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 28077 18819 28135 18825
rect 28077 18785 28089 18819
rect 28123 18816 28135 18819
rect 29822 18816 29828 18828
rect 28123 18788 29828 18816
rect 28123 18785 28135 18788
rect 28077 18779 28135 18785
rect 29822 18776 29828 18788
rect 29880 18776 29886 18828
rect 43272 18816 43300 18847
rect 45094 18816 45100 18828
rect 33980 18788 43300 18816
rect 43456 18788 45100 18816
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18717 21787 18751
rect 21729 18711 21787 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18748 25283 18751
rect 25685 18751 25743 18757
rect 25685 18748 25697 18751
rect 25271 18720 25697 18748
rect 25271 18717 25283 18720
rect 25225 18711 25283 18717
rect 25685 18717 25697 18720
rect 25731 18748 25743 18751
rect 25774 18748 25780 18760
rect 25731 18720 25780 18748
rect 25731 18717 25743 18720
rect 25685 18711 25743 18717
rect 15654 18680 15660 18692
rect 15615 18652 15660 18680
rect 15654 18640 15660 18652
rect 15712 18640 15718 18692
rect 16853 18683 16911 18689
rect 16853 18649 16865 18683
rect 16899 18649 16911 18683
rect 18966 18680 18972 18692
rect 18078 18652 18972 18680
rect 16853 18643 16911 18649
rect 13078 18612 13084 18624
rect 12084 18584 13084 18612
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 13541 18615 13599 18621
rect 13541 18581 13553 18615
rect 13587 18612 13599 18615
rect 14274 18612 14280 18624
rect 13587 18584 14280 18612
rect 13587 18581 13599 18584
rect 13541 18575 13599 18581
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 14642 18612 14648 18624
rect 14603 18584 14648 18612
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 16868 18612 16896 18643
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 21085 18683 21143 18689
rect 21085 18649 21097 18683
rect 21131 18649 21143 18683
rect 21744 18680 21772 18711
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 26697 18751 26755 18757
rect 26697 18748 26709 18751
rect 26292 18720 26709 18748
rect 26292 18708 26298 18720
rect 26697 18717 26709 18720
rect 26743 18717 26755 18751
rect 26697 18711 26755 18717
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 27154 18748 27160 18760
rect 27028 18720 27160 18748
rect 27028 18708 27034 18720
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27430 18748 27436 18760
rect 27391 18720 27436 18748
rect 27430 18708 27436 18720
rect 27488 18708 27494 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 27801 18751 27859 18757
rect 27801 18748 27813 18751
rect 27672 18720 27813 18748
rect 27672 18708 27678 18720
rect 27801 18717 27813 18720
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 28629 18751 28687 18757
rect 28629 18748 28641 18751
rect 28592 18720 28641 18748
rect 28592 18708 28598 18720
rect 28629 18717 28641 18720
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29546 18748 29552 18760
rect 29043 18720 29552 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 22186 18680 22192 18692
rect 21744 18652 22192 18680
rect 21085 18643 21143 18649
rect 18138 18612 18144 18624
rect 16868 18584 18144 18612
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 21100 18612 21128 18643
rect 22186 18640 22192 18652
rect 22244 18640 22250 18692
rect 25958 18680 25964 18692
rect 25919 18652 25964 18680
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 28350 18640 28356 18692
rect 28408 18680 28414 18692
rect 28828 18680 28856 18711
rect 29546 18708 29552 18720
rect 29604 18748 29610 18760
rect 30193 18751 30251 18757
rect 30193 18748 30205 18751
rect 29604 18720 30205 18748
rect 29604 18708 29610 18720
rect 30193 18717 30205 18720
rect 30239 18748 30251 18751
rect 30282 18748 30288 18760
rect 30239 18720 30288 18748
rect 30239 18717 30251 18720
rect 30193 18711 30251 18717
rect 30282 18708 30288 18720
rect 30340 18708 30346 18760
rect 30374 18708 30380 18760
rect 30432 18748 30438 18760
rect 30837 18751 30895 18757
rect 30432 18720 30477 18748
rect 30432 18708 30438 18720
rect 30837 18717 30849 18751
rect 30883 18717 30895 18751
rect 30837 18711 30895 18717
rect 28408 18652 28856 18680
rect 30852 18680 30880 18711
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 31665 18751 31723 18757
rect 31665 18748 31677 18751
rect 31260 18720 31677 18748
rect 31260 18708 31266 18720
rect 31665 18717 31677 18720
rect 31711 18717 31723 18751
rect 31665 18711 31723 18717
rect 32585 18751 32643 18757
rect 32585 18717 32597 18751
rect 32631 18748 32643 18751
rect 33980 18748 34008 18788
rect 43456 18757 43484 18788
rect 43257 18751 43315 18757
rect 43257 18748 43269 18751
rect 32631 18720 34008 18748
rect 35866 18720 43269 18748
rect 32631 18717 32643 18720
rect 32585 18711 32643 18717
rect 30852 18652 33456 18680
rect 28408 18640 28414 18652
rect 25590 18612 25596 18624
rect 21100 18584 25596 18612
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 33428 18612 33456 18652
rect 35866 18612 35894 18720
rect 43257 18717 43269 18720
rect 43303 18717 43315 18751
rect 43257 18711 43315 18717
rect 43441 18751 43499 18757
rect 43441 18717 43453 18751
rect 43487 18717 43499 18751
rect 43441 18711 43499 18717
rect 43272 18680 43300 18711
rect 43806 18708 43812 18760
rect 43864 18748 43870 18760
rect 44376 18757 44404 18788
rect 45094 18776 45100 18788
rect 45152 18776 45158 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 44177 18751 44235 18757
rect 44177 18748 44189 18751
rect 43864 18720 44189 18748
rect 43864 18708 43870 18720
rect 44177 18717 44189 18720
rect 44223 18717 44235 18751
rect 44177 18711 44235 18717
rect 44361 18751 44419 18757
rect 44361 18717 44373 18751
rect 44407 18717 44419 18751
rect 45002 18748 45008 18760
rect 44963 18720 45008 18748
rect 44361 18711 44419 18717
rect 45002 18708 45008 18720
rect 45060 18708 45066 18760
rect 45186 18748 45192 18760
rect 45147 18720 45192 18748
rect 45186 18708 45192 18720
rect 45244 18708 45250 18760
rect 46290 18748 46296 18760
rect 46251 18720 46296 18748
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 45373 18683 45431 18689
rect 45373 18680 45385 18683
rect 43272 18652 45385 18680
rect 45373 18649 45385 18652
rect 45419 18649 45431 18683
rect 45373 18643 45431 18649
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 33428 18584 35894 18612
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 9585 18411 9643 18417
rect 9585 18408 9597 18411
rect 9456 18380 9597 18408
rect 9456 18368 9462 18380
rect 9585 18377 9597 18380
rect 9631 18377 9643 18411
rect 10686 18408 10692 18420
rect 9585 18371 9643 18377
rect 9968 18380 10692 18408
rect 8110 18300 8116 18352
rect 8168 18340 8174 18352
rect 9968 18340 9996 18380
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 10836 18380 10885 18408
rect 10836 18368 10842 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 11885 18411 11943 18417
rect 11885 18408 11897 18411
rect 11572 18380 11897 18408
rect 11572 18368 11578 18380
rect 11885 18377 11897 18380
rect 11931 18377 11943 18411
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 11885 18371 11943 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 16390 18408 16396 18420
rect 12492 18380 16396 18408
rect 12492 18368 12498 18380
rect 16390 18368 16396 18380
rect 16448 18368 16454 18420
rect 17497 18411 17555 18417
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 17586 18408 17592 18420
rect 17543 18380 17592 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 18138 18408 18144 18420
rect 18099 18380 18144 18408
rect 18138 18368 18144 18380
rect 18196 18368 18202 18420
rect 25866 18368 25872 18420
rect 25924 18408 25930 18420
rect 46017 18411 46075 18417
rect 25924 18380 35894 18408
rect 25924 18368 25930 18380
rect 11330 18340 11336 18352
rect 8168 18312 9996 18340
rect 10060 18312 11336 18340
rect 8168 18300 8174 18312
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2406 18272 2412 18284
rect 2179 18244 2412 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2406 18232 2412 18244
rect 2464 18272 2470 18284
rect 8570 18272 8576 18284
rect 2464 18244 8576 18272
rect 2464 18232 2470 18244
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 9033 18275 9091 18281
rect 8680 18244 8892 18272
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 8680 18136 8708 18244
rect 8864 18204 8892 18244
rect 9033 18241 9045 18275
rect 9079 18272 9091 18275
rect 9122 18272 9128 18284
rect 9079 18244 9128 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9766 18272 9772 18284
rect 9727 18244 9772 18272
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10060 18281 10088 18312
rect 11330 18300 11336 18312
rect 11388 18300 11394 18352
rect 16114 18340 16120 18352
rect 11716 18312 14320 18340
rect 16075 18312 16120 18340
rect 11716 18284 11744 18312
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18241 10103 18275
rect 10226 18272 10232 18284
rect 10187 18244 10232 18272
rect 10045 18235 10103 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10778 18272 10784 18284
rect 10739 18244 10784 18272
rect 10778 18232 10784 18244
rect 10836 18232 10842 18284
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 10928 18244 11529 18272
rect 10928 18232 10934 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 11517 18235 11575 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 11974 18272 11980 18284
rect 11839 18244 11980 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 12728 18281 12756 18312
rect 14292 18284 14320 18312
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 18322 18340 18328 18352
rect 16684 18312 18328 18340
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 13538 18272 13544 18284
rect 13499 18244 13544 18272
rect 12713 18235 12771 18241
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 14274 18272 14280 18284
rect 14235 18244 14280 18272
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 16684 18281 16712 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 25222 18340 25228 18352
rect 18432 18312 25228 18340
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 17402 18272 17408 18284
rect 17363 18244 17408 18272
rect 16669 18235 16727 18241
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 17770 18232 17776 18284
rect 17828 18272 17834 18284
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 17828 18244 18061 18272
rect 17828 18232 17834 18244
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 12618 18204 12624 18216
rect 8864 18176 11928 18204
rect 12579 18176 12624 18204
rect 1627 18108 8708 18136
rect 11900 18136 11928 18176
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 13078 18204 13084 18216
rect 13039 18176 13084 18204
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 14458 18204 14464 18216
rect 14419 18176 14464 18204
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 18432 18204 18460 18312
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 28994 18300 29000 18352
rect 29052 18340 29058 18352
rect 29825 18343 29883 18349
rect 29825 18340 29837 18343
rect 29052 18312 29837 18340
rect 29052 18300 29058 18312
rect 29825 18309 29837 18312
rect 29871 18309 29883 18343
rect 32306 18340 32312 18352
rect 32267 18312 32312 18340
rect 29825 18303 29883 18309
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 20714 18272 20720 18284
rect 20487 18244 20720 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21818 18272 21824 18284
rect 21779 18244 21824 18272
rect 21818 18232 21824 18244
rect 21876 18272 21882 18284
rect 25958 18272 25964 18284
rect 21876 18244 25964 18272
rect 21876 18232 21882 18244
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26053 18275 26111 18281
rect 26053 18241 26065 18275
rect 26099 18272 26111 18275
rect 27062 18272 27068 18284
rect 26099 18244 27068 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 27062 18232 27068 18244
rect 27120 18232 27126 18284
rect 32122 18272 32128 18284
rect 32083 18244 32128 18272
rect 32122 18232 32128 18244
rect 32180 18232 32186 18284
rect 15712 18176 18460 18204
rect 20533 18207 20591 18213
rect 15712 18164 15718 18176
rect 20533 18173 20545 18207
rect 20579 18204 20591 18207
rect 21266 18204 21272 18216
rect 20579 18176 21272 18204
rect 20579 18173 20591 18176
rect 20533 18167 20591 18173
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 26145 18207 26203 18213
rect 26145 18173 26157 18207
rect 26191 18204 26203 18207
rect 26234 18204 26240 18216
rect 26191 18176 26240 18204
rect 26191 18173 26203 18176
rect 26145 18167 26203 18173
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 27157 18207 27215 18213
rect 27157 18173 27169 18207
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 27341 18207 27399 18213
rect 27341 18173 27353 18207
rect 27387 18204 27399 18207
rect 27798 18204 27804 18216
rect 27387 18176 27804 18204
rect 27387 18173 27399 18176
rect 27341 18167 27399 18173
rect 26421 18139 26479 18145
rect 11900 18108 22094 18136
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 1946 18028 1952 18080
rect 2004 18068 2010 18080
rect 2225 18071 2283 18077
rect 2225 18068 2237 18071
rect 2004 18040 2237 18068
rect 2004 18028 2010 18040
rect 2225 18037 2237 18040
rect 2271 18037 2283 18071
rect 2225 18031 2283 18037
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 13262 18068 13268 18080
rect 8628 18040 13268 18068
rect 8628 18028 8634 18040
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13412 18040 13645 18068
rect 13412 18028 13418 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 13633 18031 13691 18037
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16816 18040 16865 18068
rect 16816 18028 16822 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 20806 18068 20812 18080
rect 20767 18040 20812 18068
rect 16853 18031 16911 18037
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21913 18071 21971 18077
rect 21913 18068 21925 18071
rect 20956 18040 21925 18068
rect 20956 18028 20962 18040
rect 21913 18037 21925 18040
rect 21959 18037 21971 18071
rect 22066 18068 22094 18108
rect 26421 18105 26433 18139
rect 26467 18136 26479 18139
rect 27172 18136 27200 18167
rect 27798 18164 27804 18176
rect 27856 18164 27862 18216
rect 27890 18164 27896 18216
rect 27948 18204 27954 18216
rect 29641 18207 29699 18213
rect 27948 18176 27993 18204
rect 27948 18164 27954 18176
rect 29641 18173 29653 18207
rect 29687 18204 29699 18207
rect 30190 18204 30196 18216
rect 29687 18176 30196 18204
rect 29687 18173 29699 18176
rect 29641 18167 29699 18173
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 31478 18204 31484 18216
rect 31439 18176 31484 18204
rect 31478 18164 31484 18176
rect 31536 18164 31542 18216
rect 33962 18204 33968 18216
rect 33923 18176 33968 18204
rect 33962 18164 33968 18176
rect 34020 18164 34026 18216
rect 28166 18136 28172 18148
rect 26467 18108 28172 18136
rect 26467 18105 26479 18108
rect 26421 18099 26479 18105
rect 28166 18096 28172 18108
rect 28224 18096 28230 18148
rect 28258 18068 28264 18080
rect 22066 18040 28264 18068
rect 21913 18031 21971 18037
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 35866 18068 35894 18380
rect 46017 18377 46029 18411
rect 46063 18377 46075 18411
rect 47670 18408 47676 18420
rect 47631 18380 47676 18408
rect 46017 18371 46075 18377
rect 44910 18340 44916 18352
rect 44652 18312 44916 18340
rect 43806 18232 43812 18284
rect 43864 18272 43870 18284
rect 44652 18281 44680 18312
rect 44910 18300 44916 18312
rect 44968 18340 44974 18352
rect 46032 18340 46060 18371
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 44968 18312 46060 18340
rect 44968 18300 44974 18312
rect 44177 18275 44235 18281
rect 44177 18272 44189 18275
rect 43864 18244 44189 18272
rect 43864 18232 43870 18244
rect 44177 18241 44189 18244
rect 44223 18241 44235 18275
rect 44177 18235 44235 18241
rect 44637 18275 44695 18281
rect 44637 18241 44649 18275
rect 44683 18241 44695 18275
rect 44637 18235 44695 18241
rect 45005 18275 45063 18281
rect 45005 18241 45017 18275
rect 45051 18272 45063 18275
rect 45094 18272 45100 18284
rect 45051 18244 45100 18272
rect 45051 18241 45063 18244
rect 45005 18235 45063 18241
rect 45094 18232 45100 18244
rect 45152 18232 45158 18284
rect 45922 18272 45928 18284
rect 45883 18244 45928 18272
rect 45922 18232 45928 18244
rect 45980 18232 45986 18284
rect 46109 18275 46167 18281
rect 46109 18241 46121 18275
rect 46155 18241 46167 18275
rect 46109 18235 46167 18241
rect 44450 18164 44456 18216
rect 44508 18204 44514 18216
rect 45281 18207 45339 18213
rect 45281 18204 45293 18207
rect 44508 18176 45293 18204
rect 44508 18164 44514 18176
rect 45281 18173 45293 18176
rect 45327 18204 45339 18207
rect 46124 18204 46152 18235
rect 46290 18232 46296 18284
rect 46348 18272 46354 18284
rect 47029 18275 47087 18281
rect 47029 18272 47041 18275
rect 46348 18244 47041 18272
rect 46348 18232 46354 18244
rect 47029 18241 47041 18244
rect 47075 18241 47087 18275
rect 47029 18235 47087 18241
rect 47394 18232 47400 18284
rect 47452 18272 47458 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47452 18244 47593 18272
rect 47452 18232 47458 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 45327 18176 46152 18204
rect 45327 18173 45339 18176
rect 45281 18167 45339 18173
rect 44634 18096 44640 18148
rect 44692 18136 44698 18148
rect 45373 18139 45431 18145
rect 45373 18136 45385 18139
rect 44692 18108 45385 18136
rect 44692 18096 44698 18108
rect 45373 18105 45385 18108
rect 45419 18105 45431 18139
rect 45373 18099 45431 18105
rect 47596 18068 47624 18235
rect 35866 18040 47624 18068
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 13722 17864 13728 17876
rect 3108 17836 13728 17864
rect 3108 17824 3114 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14516 17836 14657 17864
rect 14516 17824 14522 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 23569 17867 23627 17873
rect 23569 17864 23581 17867
rect 21324 17836 23581 17864
rect 21324 17824 21330 17836
rect 23569 17833 23581 17836
rect 23615 17833 23627 17867
rect 23569 17827 23627 17833
rect 27249 17867 27307 17873
rect 27249 17833 27261 17867
rect 27295 17864 27307 17867
rect 27614 17864 27620 17876
rect 27295 17836 27620 17864
rect 27295 17833 27307 17836
rect 27249 17827 27307 17833
rect 27614 17824 27620 17836
rect 27672 17824 27678 17876
rect 27798 17864 27804 17876
rect 27759 17836 27804 17864
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 28258 17824 28264 17876
rect 28316 17864 28322 17876
rect 28442 17864 28448 17876
rect 28316 17836 28448 17864
rect 28316 17824 28322 17836
rect 28442 17824 28448 17836
rect 28500 17824 28506 17876
rect 28905 17867 28963 17873
rect 28905 17833 28917 17867
rect 28951 17864 28963 17867
rect 28994 17864 29000 17876
rect 28951 17836 29000 17864
rect 28951 17833 28963 17836
rect 28905 17827 28963 17833
rect 28994 17824 29000 17836
rect 29052 17824 29058 17876
rect 29730 17824 29736 17876
rect 29788 17864 29794 17876
rect 30009 17867 30067 17873
rect 30009 17864 30021 17867
rect 29788 17836 30021 17864
rect 29788 17824 29794 17836
rect 30009 17833 30021 17836
rect 30055 17833 30067 17867
rect 44450 17864 44456 17876
rect 44411 17836 44456 17864
rect 30009 17827 30067 17833
rect 44450 17824 44456 17836
rect 44508 17824 44514 17876
rect 45094 17824 45100 17876
rect 45152 17864 45158 17876
rect 45281 17867 45339 17873
rect 45281 17864 45293 17867
rect 45152 17836 45293 17864
rect 45152 17824 45158 17836
rect 45281 17833 45293 17836
rect 45327 17833 45339 17867
rect 45281 17827 45339 17833
rect 10781 17799 10839 17805
rect 10781 17765 10793 17799
rect 10827 17796 10839 17799
rect 11698 17796 11704 17808
rect 10827 17768 11704 17796
rect 10827 17765 10839 17768
rect 10781 17759 10839 17765
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 16390 17756 16396 17808
rect 16448 17796 16454 17808
rect 29917 17799 29975 17805
rect 16448 17768 26556 17796
rect 16448 17756 16454 17768
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 3752 17700 21189 17728
rect 3752 17688 3758 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 24670 17728 24676 17740
rect 21177 17691 21235 17697
rect 22112 17700 24676 17728
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1820 17632 2053 17660
rect 1820 17620 1826 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11146 17660 11152 17672
rect 11011 17632 11152 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 11330 17660 11336 17672
rect 11291 17632 11336 17660
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11057 17595 11115 17601
rect 11057 17561 11069 17595
rect 11103 17592 11115 17595
rect 11514 17592 11520 17604
rect 11103 17564 11520 17592
rect 11103 17561 11115 17564
rect 11057 17555 11115 17561
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 11808 17592 11836 17623
rect 13170 17620 13176 17672
rect 13228 17620 13234 17672
rect 14550 17660 14556 17672
rect 14511 17632 14556 17660
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17660 17647 17663
rect 17770 17660 17776 17672
rect 17635 17632 17776 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 20714 17660 20720 17672
rect 20627 17632 20720 17660
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 12066 17592 12072 17604
rect 11808 17564 11928 17592
rect 12027 17564 12072 17592
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11606 17524 11612 17536
rect 11195 17496 11612 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 11900 17524 11928 17564
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 15197 17595 15255 17601
rect 15197 17592 15209 17595
rect 15160 17564 15209 17592
rect 15160 17552 15166 17564
rect 15197 17561 15209 17564
rect 15243 17561 15255 17595
rect 15197 17555 15255 17561
rect 13354 17524 13360 17536
rect 11900 17496 13360 17524
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 13538 17524 13544 17536
rect 13499 17496 13544 17524
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 16448 17496 16497 17524
rect 16448 17484 16454 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 16908 17496 17601 17524
rect 16908 17484 16914 17496
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 20732 17524 20760 17620
rect 20898 17592 20904 17604
rect 20859 17564 20904 17592
rect 20898 17552 20904 17564
rect 20956 17552 20962 17604
rect 21174 17524 21180 17536
rect 20732 17496 21180 17524
rect 17589 17487 17647 17493
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 22112 17524 22140 17700
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 25590 17688 25596 17740
rect 25648 17728 25654 17740
rect 26142 17728 26148 17740
rect 25648 17700 26148 17728
rect 25648 17688 25654 17700
rect 26142 17688 26148 17700
rect 26200 17688 26206 17740
rect 26234 17688 26240 17740
rect 26292 17728 26298 17740
rect 26329 17731 26387 17737
rect 26329 17728 26341 17731
rect 26292 17700 26341 17728
rect 26292 17688 26298 17700
rect 26329 17697 26341 17700
rect 26375 17697 26387 17731
rect 26528 17728 26556 17768
rect 29917 17765 29929 17799
rect 29963 17796 29975 17799
rect 30282 17796 30288 17808
rect 29963 17768 30288 17796
rect 29963 17765 29975 17768
rect 29917 17759 29975 17765
rect 30282 17756 30288 17768
rect 30340 17756 30346 17808
rect 26528 17700 35894 17728
rect 26329 17691 26387 17697
rect 25504 17672 25556 17678
rect 22922 17620 22928 17672
rect 22980 17660 22986 17672
rect 23106 17660 23112 17672
rect 22980 17632 23112 17660
rect 22980 17620 22986 17632
rect 23106 17620 23112 17632
rect 23164 17660 23170 17672
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 23164 17632 23397 17660
rect 23164 17620 23170 17632
rect 23385 17629 23397 17632
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 26160 17660 26188 17688
rect 26881 17663 26939 17669
rect 26881 17660 26893 17663
rect 25556 17626 25636 17654
rect 26160 17632 26893 17660
rect 25504 17614 25556 17620
rect 22186 17552 22192 17604
rect 22244 17592 22250 17604
rect 23017 17595 23075 17601
rect 23017 17592 23029 17595
rect 22244 17564 23029 17592
rect 22244 17552 22250 17564
rect 23017 17561 23029 17564
rect 23063 17561 23075 17595
rect 23017 17555 23075 17561
rect 23201 17595 23259 17601
rect 23201 17561 23213 17595
rect 23247 17592 23259 17595
rect 23474 17592 23480 17604
rect 23247 17564 23480 17592
rect 23247 17561 23259 17564
rect 23201 17555 23259 17561
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 25608 17592 25636 17626
rect 26881 17629 26893 17632
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17660 27767 17663
rect 27982 17660 27988 17672
rect 27755 17632 27988 17660
rect 27755 17629 27767 17632
rect 27709 17623 27767 17629
rect 27080 17592 27108 17623
rect 27982 17620 27988 17632
rect 28040 17660 28046 17672
rect 28813 17663 28871 17669
rect 28813 17660 28825 17663
rect 28040 17632 28825 17660
rect 28040 17620 28046 17632
rect 28813 17629 28825 17632
rect 28859 17629 28871 17663
rect 29546 17660 29552 17672
rect 29507 17632 29552 17660
rect 28813 17623 28871 17629
rect 29546 17620 29552 17632
rect 29604 17620 29610 17672
rect 25608 17564 27108 17592
rect 23290 17524 23296 17536
rect 21324 17496 22140 17524
rect 23251 17496 23296 17524
rect 21324 17484 21330 17496
rect 23290 17484 23296 17496
rect 23348 17524 23354 17536
rect 23934 17524 23940 17536
rect 23348 17496 23940 17524
rect 23348 17484 23354 17496
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 35866 17524 35894 17700
rect 43530 17620 43536 17672
rect 43588 17660 43594 17672
rect 44085 17663 44143 17669
rect 44085 17660 44097 17663
rect 43588 17632 44097 17660
rect 43588 17620 43594 17632
rect 44085 17629 44097 17632
rect 44131 17629 44143 17663
rect 44266 17660 44272 17672
rect 44227 17632 44272 17660
rect 44085 17623 44143 17629
rect 44100 17592 44128 17623
rect 44266 17620 44272 17632
rect 44324 17620 44330 17672
rect 46290 17660 46296 17672
rect 46251 17632 46296 17660
rect 46290 17620 46296 17632
rect 46348 17620 46354 17672
rect 44450 17592 44456 17604
rect 44100 17564 44456 17592
rect 44450 17552 44456 17564
rect 44508 17552 44514 17604
rect 45002 17592 45008 17604
rect 44963 17564 45008 17592
rect 45002 17552 45008 17564
rect 45060 17552 45066 17604
rect 45186 17592 45192 17604
rect 45147 17564 45192 17592
rect 45186 17552 45192 17564
rect 45244 17552 45250 17604
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 44818 17524 44824 17536
rect 35866 17496 44824 17524
rect 44818 17484 44824 17496
rect 44876 17524 44882 17536
rect 47394 17524 47400 17536
rect 44876 17496 47400 17524
rect 44876 17484 44882 17496
rect 47394 17484 47400 17496
rect 47452 17484 47458 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 11885 17323 11943 17329
rect 11885 17289 11897 17323
rect 11931 17320 11943 17323
rect 12618 17320 12624 17332
rect 11931 17292 12624 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 13170 17320 13176 17332
rect 13131 17292 13176 17320
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 21174 17320 21180 17332
rect 21135 17292 21180 17320
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 23106 17280 23112 17332
rect 23164 17329 23170 17332
rect 23164 17323 23183 17329
rect 23171 17320 23183 17323
rect 23171 17292 24072 17320
rect 23171 17289 23183 17292
rect 23164 17283 23183 17289
rect 23164 17280 23170 17283
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 11517 17255 11575 17261
rect 11517 17252 11529 17255
rect 11204 17224 11529 17252
rect 11204 17212 11210 17224
rect 11517 17221 11529 17224
rect 11563 17221 11575 17255
rect 11517 17215 11575 17221
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 11532 17184 11560 17215
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 11733 17255 11791 17261
rect 11733 17252 11745 17255
rect 11664 17224 11745 17252
rect 11664 17212 11670 17224
rect 11733 17221 11745 17224
rect 11779 17252 11791 17255
rect 18598 17252 18604 17264
rect 11779 17224 12664 17252
rect 18354 17224 18604 17252
rect 11779 17221 11791 17224
rect 11733 17215 11791 17221
rect 11974 17184 11980 17196
rect 11532 17156 11980 17184
rect 11974 17144 11980 17156
rect 12032 17184 12038 17196
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 12032 17156 12357 17184
rect 12032 17144 12038 17156
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12636 17193 12664 17224
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 20714 17212 20720 17264
rect 20772 17212 20778 17264
rect 22925 17255 22983 17261
rect 22925 17221 22937 17255
rect 22971 17252 22983 17255
rect 23474 17252 23480 17264
rect 22971 17224 23480 17252
rect 22971 17221 22983 17224
rect 22925 17215 22983 17221
rect 23474 17212 23480 17224
rect 23532 17252 23538 17264
rect 23934 17252 23940 17264
rect 23532 17224 23796 17252
rect 23895 17224 23940 17252
rect 23532 17212 23538 17224
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12492 17156 12541 17184
rect 12492 17144 12498 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17184 12679 17187
rect 12710 17184 12716 17196
rect 12667 17156 12716 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12860 17156 13093 17184
rect 12860 17144 12866 17156
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 13170 17184 13176 17196
rect 13127 17156 13176 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 14056 17156 14381 17184
rect 14056 17144 14062 17156
rect 14369 17153 14381 17156
rect 14415 17184 14427 17187
rect 14550 17184 14556 17196
rect 14415 17156 14556 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 14642 17144 14648 17196
rect 14700 17184 14706 17196
rect 15102 17184 15108 17196
rect 14700 17156 15108 17184
rect 14700 17144 14706 17156
rect 15102 17144 15108 17156
rect 15160 17184 15166 17196
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 15160 17156 15209 17184
rect 15160 17144 15166 17156
rect 15197 17153 15209 17156
rect 15243 17153 15255 17187
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 15197 17147 15255 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 23768 17193 23796 17224
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 23842 17184 23848 17196
rect 23799 17156 23848 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 24044 17193 24072 17292
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 25501 17323 25559 17329
rect 25501 17320 25513 17323
rect 24728 17292 25513 17320
rect 24728 17280 24734 17292
rect 25501 17289 25513 17292
rect 25547 17289 25559 17323
rect 25501 17283 25559 17289
rect 27157 17323 27215 17329
rect 27157 17289 27169 17323
rect 27203 17320 27215 17323
rect 27246 17320 27252 17332
rect 27203 17292 27252 17320
rect 27203 17289 27215 17292
rect 27157 17283 27215 17289
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 45002 17280 45008 17332
rect 45060 17320 45066 17332
rect 46201 17323 46259 17329
rect 46201 17320 46213 17323
rect 45060 17292 46213 17320
rect 45060 17280 45066 17292
rect 46201 17289 46213 17292
rect 46247 17289 46259 17323
rect 47670 17320 47676 17332
rect 47631 17292 47676 17320
rect 46201 17283 46259 17289
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 44361 17255 44419 17261
rect 44361 17221 44373 17255
rect 44407 17252 44419 17255
rect 45922 17252 45928 17264
rect 44407 17224 45928 17252
rect 44407 17221 44419 17224
rect 44361 17215 44419 17221
rect 45922 17212 45928 17224
rect 45980 17212 45986 17264
rect 46290 17212 46296 17264
rect 46348 17252 46354 17264
rect 46348 17224 47072 17252
rect 46348 17212 46354 17224
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 25409 17187 25467 17193
rect 25409 17153 25421 17187
rect 25455 17153 25467 17187
rect 26970 17184 26976 17196
rect 26931 17156 26976 17184
rect 25409 17147 25467 17153
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 15930 17116 15936 17128
rect 3016 17088 12388 17116
rect 15891 17088 15936 17116
rect 3016 17076 3022 17088
rect 12360 17048 12388 17088
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 18322 17116 18328 17128
rect 17175 17088 18328 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18564 17088 18613 17116
rect 18564 17076 18570 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 19426 17116 19432 17128
rect 19387 17088 19432 17116
rect 18601 17079 18659 17085
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 19751 17088 20852 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 15948 17048 15976 17076
rect 20824 17060 20852 17088
rect 21082 17076 21088 17128
rect 21140 17116 21146 17128
rect 25424 17116 25452 17147
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27430 17184 27436 17196
rect 27203 17156 27436 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 44266 17184 44272 17196
rect 44179 17156 44272 17184
rect 44266 17144 44272 17156
rect 44324 17144 44330 17196
rect 44450 17184 44456 17196
rect 44411 17156 44456 17184
rect 44450 17144 44456 17156
rect 44508 17144 44514 17196
rect 46382 17184 46388 17196
rect 46343 17156 46388 17184
rect 46382 17144 46388 17156
rect 46440 17144 46446 17196
rect 47044 17193 47072 17224
rect 47029 17187 47087 17193
rect 47029 17153 47041 17187
rect 47075 17153 47087 17187
rect 47029 17147 47087 17153
rect 47394 17144 47400 17196
rect 47452 17184 47458 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47452 17156 47593 17184
rect 47452 17144 47458 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 21140 17088 25452 17116
rect 44284 17116 44312 17144
rect 46198 17116 46204 17128
rect 44284 17088 46204 17116
rect 21140 17076 21146 17088
rect 46198 17076 46204 17088
rect 46256 17076 46262 17128
rect 12360 17020 15976 17048
rect 20806 17008 20812 17060
rect 20864 17008 20870 17060
rect 23198 17048 23204 17060
rect 23124 17020 23204 17048
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11664 16952 11713 16980
rect 11664 16940 11670 16952
rect 11701 16949 11713 16952
rect 11747 16980 11759 16983
rect 12158 16980 12164 16992
rect 11747 16952 12164 16980
rect 11747 16949 11759 16952
rect 11701 16943 11759 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12342 16980 12348 16992
rect 12303 16952 12348 16980
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 14461 16983 14519 16989
rect 14461 16949 14473 16983
rect 14507 16980 14519 16983
rect 14550 16980 14556 16992
rect 14507 16952 14556 16980
rect 14507 16949 14519 16952
rect 14461 16943 14519 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 21266 16980 21272 16992
rect 19116 16952 21272 16980
rect 19116 16940 19122 16952
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 23124 16989 23152 17020
rect 23198 17008 23204 17020
rect 23256 17008 23262 17060
rect 23109 16983 23167 16989
rect 23109 16949 23121 16983
rect 23155 16949 23167 16983
rect 23290 16980 23296 16992
rect 23251 16952 23296 16980
rect 23109 16943 23167 16949
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 23750 16980 23756 16992
rect 23711 16952 23756 16980
rect 23750 16940 23756 16952
rect 23808 16940 23814 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 11885 16779 11943 16785
rect 11885 16745 11897 16779
rect 11931 16776 11943 16779
rect 12066 16776 12072 16788
rect 11931 16748 12072 16776
rect 11931 16745 11943 16748
rect 11885 16739 11943 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 16945 16779 17003 16785
rect 16945 16745 16957 16779
rect 16991 16776 17003 16779
rect 17770 16776 17776 16788
rect 16991 16748 17776 16776
rect 16991 16745 17003 16748
rect 16945 16739 17003 16745
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 19484 16748 19533 16776
rect 19484 16736 19490 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 47026 16776 47032 16788
rect 19521 16739 19579 16745
rect 19628 16748 47032 16776
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 13538 16708 13544 16720
rect 12032 16680 13544 16708
rect 12032 16668 12038 16680
rect 13538 16668 13544 16680
rect 13596 16708 13602 16720
rect 13596 16680 14412 16708
rect 13596 16668 13602 16680
rect 12342 16640 12348 16652
rect 11900 16612 12348 16640
rect 11900 16581 11928 16612
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12618 16640 12624 16652
rect 12452 16612 12624 16640
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16574 11943 16575
rect 12069 16575 12127 16581
rect 11931 16546 11965 16574
rect 11931 16541 11943 16546
rect 11885 16535 11943 16541
rect 12069 16541 12081 16575
rect 12115 16572 12127 16575
rect 12452 16572 12480 16612
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 14384 16649 14412 16680
rect 15930 16668 15936 16720
rect 15988 16708 15994 16720
rect 19628 16708 19656 16748
rect 47026 16736 47032 16748
rect 47084 16736 47090 16788
rect 15988 16680 19656 16708
rect 15988 16668 15994 16680
rect 20622 16668 20628 16720
rect 20680 16708 20686 16720
rect 21082 16708 21088 16720
rect 20680 16680 21088 16708
rect 20680 16668 20686 16680
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 23290 16708 23296 16720
rect 22112 16680 23296 16708
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16609 14427 16643
rect 14550 16640 14556 16652
rect 14511 16612 14556 16640
rect 14369 16603 14427 16609
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 19058 16640 19064 16652
rect 18524 16612 19064 16640
rect 16758 16572 16764 16584
rect 12115 16544 12480 16572
rect 16719 16544 16764 16572
rect 12115 16541 12127 16544
rect 12069 16535 12127 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 18524 16581 18552 16612
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 22112 16649 22140 16680
rect 23290 16668 23296 16680
rect 23348 16708 23354 16720
rect 23348 16680 23888 16708
rect 23348 16668 23354 16680
rect 22097 16643 22155 16649
rect 22097 16609 22109 16643
rect 22143 16609 22155 16643
rect 22370 16640 22376 16652
rect 22331 16612 22376 16640
rect 22097 16603 22155 16609
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23750 16640 23756 16652
rect 23492 16612 23756 16640
rect 17497 16575 17555 16581
rect 17497 16572 17509 16575
rect 17000 16544 17509 16572
rect 17000 16532 17006 16544
rect 17497 16541 17509 16544
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 18656 16544 18701 16572
rect 18656 16532 18662 16544
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19337 16575 19395 16581
rect 19337 16572 19349 16575
rect 19300 16544 19349 16572
rect 19300 16532 19306 16544
rect 19337 16541 19349 16544
rect 19383 16541 19395 16575
rect 19337 16535 19395 16541
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20312 16544 20361 16572
rect 20312 16532 20318 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16572 20499 16575
rect 20714 16572 20720 16584
rect 20487 16544 20720 16572
rect 20487 16541 20499 16544
rect 20441 16535 20499 16541
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 21174 16572 21180 16584
rect 21135 16544 21180 16572
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16572 22063 16575
rect 22186 16572 22192 16584
rect 22051 16544 22192 16572
rect 22051 16541 22063 16544
rect 22005 16535 22063 16541
rect 22186 16532 22192 16544
rect 22244 16572 22250 16584
rect 22646 16572 22652 16584
rect 22244 16544 22652 16572
rect 22244 16532 22250 16544
rect 22646 16532 22652 16544
rect 22704 16532 22710 16584
rect 22830 16581 22836 16584
rect 22825 16572 22836 16581
rect 22791 16544 22836 16572
rect 22825 16535 22836 16544
rect 22830 16532 22836 16535
rect 22888 16532 22894 16584
rect 23492 16581 23520 16612
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 23860 16572 23888 16680
rect 23934 16600 23940 16652
rect 23992 16640 23998 16652
rect 24670 16640 24676 16652
rect 23992 16612 24676 16640
rect 23992 16600 23998 16612
rect 24670 16600 24676 16612
rect 24728 16640 24734 16652
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 24728 16612 25881 16640
rect 24728 16600 24734 16612
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 27522 16640 27528 16652
rect 27483 16612 27528 16640
rect 25869 16603 25927 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 46293 16643 46351 16649
rect 28684 16612 28856 16640
rect 28684 16600 28690 16612
rect 23707 16544 23888 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 24302 16532 24308 16584
rect 24360 16572 24366 16584
rect 28828 16581 28856 16612
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 24360 16544 24409 16572
rect 24360 16532 24366 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16541 28871 16575
rect 29546 16572 29552 16584
rect 29507 16544 29552 16572
rect 28813 16535 28871 16541
rect 29546 16532 29552 16544
rect 29604 16532 29610 16584
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 38654 16572 38660 16584
rect 31435 16544 38660 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 38654 16532 38660 16544
rect 38712 16532 38718 16584
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 26050 16504 26056 16516
rect 16255 16476 25912 16504
rect 26011 16476 26056 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 17586 16436 17592 16448
rect 17547 16408 17592 16436
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16436 21327 16439
rect 22830 16436 22836 16448
rect 21315 16408 22836 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 23566 16436 23572 16448
rect 22980 16408 23025 16436
rect 23527 16408 23572 16436
rect 22980 16396 22986 16408
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 24486 16436 24492 16448
rect 24447 16408 24492 16436
rect 24486 16396 24492 16408
rect 24544 16396 24550 16448
rect 25884 16436 25912 16476
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 28905 16507 28963 16513
rect 28905 16473 28917 16507
rect 28951 16504 28963 16507
rect 29733 16507 29791 16513
rect 29733 16504 29745 16507
rect 28951 16476 29745 16504
rect 28951 16473 28963 16476
rect 28905 16467 28963 16473
rect 29733 16473 29745 16476
rect 29779 16473 29791 16507
rect 45554 16504 45560 16516
rect 29733 16467 29791 16473
rect 31726 16476 45560 16504
rect 31726 16436 31754 16476
rect 45554 16464 45560 16476
rect 45612 16464 45618 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 46842 16504 46848 16516
rect 46523 16476 46848 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 46842 16464 46848 16476
rect 46900 16464 46906 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 25884 16408 31754 16436
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 16942 16232 16948 16244
rect 16040 16204 16948 16232
rect 11698 16096 11704 16108
rect 11659 16068 11704 16096
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 13170 16096 13176 16108
rect 12299 16068 13176 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 14642 16096 14648 16108
rect 14603 16068 14648 16096
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16040 16096 16068 16204
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 25314 16232 25320 16244
rect 18472 16204 24624 16232
rect 18472 16192 18478 16204
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16592 16136 16865 16164
rect 16592 16108 16620 16136
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 24486 16164 24492 16176
rect 24334 16136 24492 16164
rect 16853 16127 16911 16133
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 24596 16164 24624 16204
rect 24780 16204 25320 16232
rect 24780 16164 24808 16204
rect 25314 16192 25320 16204
rect 25372 16232 25378 16244
rect 46842 16232 46848 16244
rect 25372 16204 41414 16232
rect 46803 16204 46848 16232
rect 25372 16192 25378 16204
rect 38194 16164 38200 16176
rect 24596 16136 24808 16164
rect 25332 16136 38200 16164
rect 15979 16068 16068 16096
rect 16117 16099 16175 16105
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16574 16096 16580 16108
rect 16163 16068 16580 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 16942 16096 16948 16108
rect 16715 16068 16948 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 17083 16068 17693 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 17911 16068 18521 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 19058 16096 19064 16108
rect 19019 16068 19064 16096
rect 18509 16059 18567 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 19300 16068 20913 16096
rect 19300 16056 19306 16068
rect 20901 16065 20913 16068
rect 20947 16096 20959 16099
rect 21174 16096 21180 16108
rect 20947 16068 21180 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 22830 16096 22836 16108
rect 22791 16068 22836 16096
rect 22830 16056 22836 16068
rect 22888 16056 22894 16108
rect 25222 16096 25228 16108
rect 25183 16068 25228 16096
rect 25222 16056 25228 16068
rect 25280 16096 25286 16108
rect 25332 16096 25360 16136
rect 38194 16124 38200 16136
rect 38252 16124 38258 16176
rect 25958 16096 25964 16108
rect 25280 16068 25360 16096
rect 25919 16068 25964 16096
rect 25280 16056 25286 16068
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 26050 16056 26056 16108
rect 26108 16096 26114 16108
rect 28166 16096 28172 16108
rect 26108 16068 26153 16096
rect 28127 16068 28172 16096
rect 26108 16056 26114 16068
rect 28166 16056 28172 16068
rect 28224 16056 28230 16108
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16096 30067 16099
rect 30466 16096 30472 16108
rect 30055 16068 30472 16096
rect 30055 16065 30067 16068
rect 30009 16059 30067 16065
rect 30466 16056 30472 16068
rect 30524 16056 30530 16108
rect 41386 16096 41414 16204
rect 46842 16192 46848 16204
rect 46900 16192 46906 16244
rect 46753 16099 46811 16105
rect 46753 16096 46765 16099
rect 41386 16068 46765 16096
rect 46753 16065 46765 16068
rect 46799 16065 46811 16099
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 46753 16059 46811 16065
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 16028 16083 16031
rect 17126 16028 17132 16040
rect 16071 16000 17132 16028
rect 16071 15997 16083 16000
rect 16025 15991 16083 15997
rect 17126 15988 17132 16000
rect 17184 16028 17190 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17184 16000 17509 16028
rect 17184 15988 17190 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 23109 16031 23167 16037
rect 23109 15997 23121 16031
rect 23155 16028 23167 16031
rect 23566 16028 23572 16040
rect 23155 16000 23572 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 23566 15988 23572 16000
rect 23624 15988 23630 16040
rect 24581 16031 24639 16037
rect 24581 15997 24593 16031
rect 24627 16028 24639 16031
rect 24670 16028 24676 16040
rect 24627 16000 24676 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 28353 16031 28411 16037
rect 28353 15997 28365 16031
rect 28399 16028 28411 16031
rect 28442 16028 28448 16040
rect 28399 16000 28448 16028
rect 28399 15997 28411 16000
rect 28353 15991 28411 15997
rect 28442 15988 28448 16000
rect 28500 15988 28506 16040
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 19242 15960 19248 15972
rect 16816 15932 19248 15960
rect 16816 15920 16822 15932
rect 19242 15920 19248 15932
rect 19300 15920 19306 15972
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11112 15864 11529 15892
rect 11112 15852 11118 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 12342 15892 12348 15904
rect 12303 15864 12348 15892
rect 11517 15855 11575 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14737 15895 14795 15901
rect 14737 15892 14749 15895
rect 14056 15864 14749 15892
rect 14056 15852 14062 15864
rect 14737 15861 14749 15864
rect 14783 15861 14795 15895
rect 14737 15855 14795 15861
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 18414 15892 18420 15904
rect 16448 15864 18420 15892
rect 16448 15852 16454 15864
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 19153 15895 19211 15901
rect 19153 15861 19165 15895
rect 19199 15892 19211 15895
rect 19334 15892 19340 15904
rect 19199 15864 19340 15892
rect 19199 15861 19211 15864
rect 19153 15855 19211 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 21082 15892 21088 15904
rect 21043 15864 21088 15892
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 25314 15892 25320 15904
rect 25275 15864 25320 15892
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 12710 15688 12716 15700
rect 10336 15660 12716 15688
rect 10336 15561 10364 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 17586 15648 17592 15700
rect 17644 15688 17650 15700
rect 17644 15660 22600 15688
rect 17644 15648 17650 15660
rect 10597 15623 10655 15629
rect 10597 15589 10609 15623
rect 10643 15620 10655 15623
rect 22572 15620 22600 15660
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 22833 15691 22891 15697
rect 22833 15688 22845 15691
rect 22704 15660 22845 15688
rect 22704 15648 22710 15660
rect 22833 15657 22845 15660
rect 22879 15657 22891 15691
rect 22833 15651 22891 15657
rect 29546 15620 29552 15632
rect 10643 15592 11192 15620
rect 22572 15592 29552 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15521 10379 15555
rect 11054 15552 11060 15564
rect 11015 15524 11060 15552
rect 10321 15515 10379 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 11164 15552 11192 15592
rect 29546 15580 29552 15592
rect 29604 15580 29610 15632
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 11164 15524 11345 15552
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 12066 15552 12072 15564
rect 11848 15524 12072 15552
rect 11848 15512 11854 15524
rect 12066 15512 12072 15524
rect 12124 15552 12130 15564
rect 13081 15555 13139 15561
rect 13081 15552 13093 15555
rect 12124 15524 13093 15552
rect 12124 15512 12130 15524
rect 13081 15521 13093 15524
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 16942 15552 16948 15564
rect 15703 15524 16948 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17126 15552 17132 15564
rect 17087 15524 17132 15552
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 21082 15552 21088 15564
rect 21043 15524 21088 15552
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 21361 15555 21419 15561
rect 21361 15521 21373 15555
rect 21407 15552 21419 15555
rect 22370 15552 22376 15564
rect 21407 15524 22376 15552
rect 21407 15521 21419 15524
rect 21361 15515 21419 15521
rect 22370 15512 22376 15524
rect 22428 15512 22434 15564
rect 22922 15552 22928 15564
rect 22480 15524 22928 15552
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10244 15348 10272 15447
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 12400 15456 12466 15484
rect 12400 15444 12406 15456
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 15252 15456 15393 15484
rect 15252 15444 15258 15456
rect 15381 15453 15393 15456
rect 15427 15484 15439 15487
rect 15746 15484 15752 15496
rect 15427 15456 15752 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15416 14611 15419
rect 16758 15416 16764 15428
rect 14599 15388 16764 15416
rect 14599 15385 14611 15388
rect 14553 15379 14611 15385
rect 16758 15376 16764 15388
rect 16816 15376 16822 15428
rect 17034 15376 17040 15428
rect 17092 15416 17098 15428
rect 17236 15416 17264 15447
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17828 15456 18061 15484
rect 17828 15444 17834 15456
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 22480 15470 22508 15524
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 25314 15552 25320 15564
rect 25275 15524 25320 15552
rect 25314 15512 25320 15524
rect 25372 15512 25378 15564
rect 26694 15552 26700 15564
rect 26655 15524 26700 15552
rect 26694 15512 26700 15524
rect 26752 15512 26758 15564
rect 25133 15487 25191 15493
rect 25133 15484 25145 15487
rect 18049 15447 18107 15453
rect 22756 15456 25145 15484
rect 17092 15388 20024 15416
rect 17092 15376 17098 15388
rect 19996 15360 20024 15388
rect 12066 15348 12072 15360
rect 10244 15320 12072 15348
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 14826 15348 14832 15360
rect 14787 15320 14832 15348
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 17589 15351 17647 15357
rect 17589 15317 17601 15351
rect 17635 15348 17647 15351
rect 17954 15348 17960 15360
rect 17635 15320 17960 15348
rect 17635 15317 17647 15320
rect 17589 15311 17647 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18046 15308 18052 15360
rect 18104 15348 18110 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18104 15320 18245 15348
rect 18104 15308 18110 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 22756 15348 22784 15456
rect 25133 15453 25145 15456
rect 25179 15453 25191 15487
rect 25133 15447 25191 15453
rect 20036 15320 22784 15348
rect 20036 15308 20042 15320
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 18506 15144 18512 15156
rect 15059 15116 18512 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15105 15079 15163 15085
rect 15105 15045 15117 15079
rect 15151 15076 15163 15079
rect 15286 15076 15292 15088
rect 15151 15048 15292 15076
rect 15151 15045 15163 15048
rect 15105 15039 15163 15045
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 11698 15008 11704 15020
rect 11611 14980 11704 15008
rect 11698 14968 11704 14980
rect 11756 15008 11762 15020
rect 12250 15008 12256 15020
rect 11756 14980 12256 15008
rect 11756 14968 11762 14980
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12894 15008 12900 15020
rect 12575 14980 12900 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13170 15008 13176 15020
rect 13131 14980 13176 15008
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 16132 15017 16160 15116
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 19797 15147 19855 15153
rect 19797 15113 19809 15147
rect 19843 15144 19855 15147
rect 19978 15144 19984 15156
rect 19843 15116 19984 15144
rect 19843 15113 19855 15116
rect 19797 15107 19855 15113
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 16942 15076 16948 15088
rect 16868 15048 16948 15076
rect 16868 15017 16896 15048
rect 16942 15036 16948 15048
rect 17000 15036 17006 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18325 15079 18383 15085
rect 18325 15076 18337 15079
rect 18012 15048 18337 15076
rect 18012 15036 18018 15048
rect 18325 15045 18337 15048
rect 18371 15045 18383 15079
rect 18325 15039 18383 15045
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 16117 15011 16175 15017
rect 15252 14980 15297 15008
rect 15252 14968 15258 14980
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 16853 14971 16911 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 18046 15008 18052 15020
rect 18007 14980 18052 15008
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12912 14940 12940 14968
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 12912 14912 15393 14940
rect 12345 14903 12403 14909
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14909 17003 14943
rect 17126 14940 17132 14952
rect 17087 14912 17132 14940
rect 16945 14903 17003 14909
rect 12360 14872 12388 14903
rect 14829 14875 14887 14881
rect 12360 14844 14688 14872
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 11480 14776 11529 14804
rect 11480 14764 11486 14776
rect 11517 14773 11529 14776
rect 11563 14773 11575 14807
rect 12710 14804 12716 14816
rect 12671 14776 12716 14804
rect 11517 14767 11575 14773
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 14660 14804 14688 14844
rect 14829 14841 14841 14875
rect 14875 14872 14887 14875
rect 14918 14872 14924 14884
rect 14875 14844 14924 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 16574 14872 16580 14884
rect 16040 14844 16580 14872
rect 16040 14816 16068 14844
rect 16574 14832 16580 14844
rect 16632 14872 16638 14884
rect 16960 14872 16988 14903
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 16632 14844 16988 14872
rect 16632 14832 16638 14844
rect 15102 14804 15108 14816
rect 14660 14776 15108 14804
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15933 14807 15991 14813
rect 15933 14773 15945 14807
rect 15979 14804 15991 14807
rect 16022 14804 16028 14816
rect 15979 14776 16028 14804
rect 15979 14773 15991 14776
rect 15933 14767 15991 14773
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16669 14807 16727 14813
rect 16669 14773 16681 14807
rect 16715 14804 16727 14807
rect 17218 14804 17224 14816
rect 16715 14776 17224 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 17126 14600 17132 14612
rect 15948 14572 17132 14600
rect 6886 14504 11560 14532
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 6886 14396 6914 14504
rect 11422 14464 11428 14476
rect 11383 14436 11428 14464
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 11532 14464 11560 14504
rect 14918 14492 14924 14544
rect 14976 14532 14982 14544
rect 15948 14541 15976 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 15933 14535 15991 14541
rect 15933 14532 15945 14535
rect 14976 14504 15945 14532
rect 14976 14492 14982 14504
rect 15933 14501 15945 14504
rect 15979 14501 15991 14535
rect 15933 14495 15991 14501
rect 16114 14492 16120 14544
rect 16172 14532 16178 14544
rect 17034 14532 17040 14544
rect 16172 14504 17040 14532
rect 16172 14492 16178 14504
rect 17034 14492 17040 14504
rect 17092 14492 17098 14544
rect 17218 14532 17224 14544
rect 17179 14504 17224 14532
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 27706 14464 27712 14476
rect 11532 14436 27712 14464
rect 27706 14424 27712 14436
rect 27764 14424 27770 14476
rect 2188 14368 6914 14396
rect 15105 14399 15163 14405
rect 2188 14356 2194 14368
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 16022 14396 16028 14408
rect 15151 14368 16028 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 16022 14356 16028 14368
rect 16080 14396 16086 14408
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 16080 14368 16221 14396
rect 16080 14356 16086 14368
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16850 14396 16856 14408
rect 16347 14368 16856 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 18049 14399 18107 14405
rect 18049 14396 18061 14399
rect 17420 14368 18061 14396
rect 11698 14328 11704 14340
rect 11659 14300 11704 14328
rect 11698 14288 11704 14300
rect 11756 14288 11762 14340
rect 13262 14328 13268 14340
rect 12926 14300 13268 14328
rect 13262 14288 13268 14300
rect 13320 14288 13326 14340
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 14918 14328 14924 14340
rect 14332 14300 14924 14328
rect 14332 14288 14338 14300
rect 14918 14288 14924 14300
rect 14976 14288 14982 14340
rect 15286 14328 15292 14340
rect 15199 14300 15292 14328
rect 15286 14288 15292 14300
rect 15344 14328 15350 14340
rect 15838 14328 15844 14340
rect 15344 14300 15844 14328
rect 15344 14288 15350 14300
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 16114 14328 16120 14340
rect 16075 14300 16120 14328
rect 16114 14288 16120 14300
rect 16172 14288 16178 14340
rect 16945 14331 17003 14337
rect 16945 14297 16957 14331
rect 16991 14297 17003 14331
rect 16945 14291 17003 14297
rect 13170 14260 13176 14272
rect 13131 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15197 14263 15255 14269
rect 15197 14260 15209 14263
rect 15160 14232 15209 14260
rect 15160 14220 15166 14232
rect 15197 14229 15209 14232
rect 15243 14229 15255 14263
rect 15197 14223 15255 14229
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 15436 14232 15485 14260
rect 15436 14220 15442 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 16482 14260 16488 14272
rect 16443 14232 16488 14260
rect 15473 14223 15531 14229
rect 16482 14220 16488 14232
rect 16540 14260 16546 14272
rect 16960 14260 16988 14291
rect 17420 14269 17448 14368
rect 18049 14365 18061 14368
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14396 19395 14399
rect 20622 14396 20628 14408
rect 19383 14368 20628 14396
rect 19383 14365 19395 14368
rect 19337 14359 19395 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 16540 14232 16988 14260
rect 17405 14263 17463 14269
rect 16540 14220 16546 14232
rect 17405 14229 17417 14263
rect 17451 14229 17463 14263
rect 17862 14260 17868 14272
rect 17823 14232 17868 14260
rect 17405 14223 17463 14229
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 18472 14232 19533 14260
rect 18472 14220 18478 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 19521 14223 19579 14229
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11756 14028 11897 14056
rect 11756 14016 11762 14028
rect 11885 14025 11897 14028
rect 11931 14025 11943 14059
rect 11885 14019 11943 14025
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 15194 14056 15200 14068
rect 14139 14028 15200 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 17184 14028 19073 14056
rect 17184 14016 17190 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 12710 13988 12716 14000
rect 12084 13960 12716 13988
rect 12084 13929 12112 13960
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 13725 13991 13783 13997
rect 13725 13957 13737 13991
rect 13771 13957 13783 13991
rect 13725 13951 13783 13957
rect 13941 13991 13999 13997
rect 13941 13957 13953 13991
rect 13987 13988 13999 13991
rect 14550 13988 14556 14000
rect 13987 13960 14556 13988
rect 13987 13957 13999 13960
rect 13941 13951 13999 13957
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12434 13920 12440 13932
rect 12391 13892 12440 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 13170 13920 13176 13932
rect 12575 13892 13176 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12544 13852 12572 13883
rect 13170 13880 13176 13892
rect 13228 13920 13234 13932
rect 13740 13920 13768 13951
rect 14550 13948 14556 13960
rect 14608 13948 14614 14000
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 17862 13988 17868 14000
rect 17635 13960 17868 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 18598 13948 18604 14000
rect 18656 13948 18662 14000
rect 13228 13892 13768 13920
rect 13228 13880 13234 13892
rect 17310 13852 17316 13864
rect 11756 13824 12572 13852
rect 17271 13824 17316 13852
rect 11756 13812 11762 13824
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 15470 13784 15476 13796
rect 3476 13756 15476 13784
rect 3476 13744 3482 13756
rect 15470 13744 15476 13756
rect 15528 13744 15534 13796
rect 13906 13716 13912 13728
rect 13867 13688 13912 13716
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 12621 13515 12679 13521
rect 12621 13481 12633 13515
rect 12667 13512 12679 13515
rect 14550 13512 14556 13524
rect 12667 13484 14556 13512
rect 12667 13481 12679 13484
rect 12621 13475 12679 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 15746 13512 15752 13524
rect 15703 13484 15752 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 15838 13472 15844 13524
rect 15896 13512 15902 13524
rect 15896 13484 15941 13512
rect 15896 13472 15902 13484
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17368 13484 17417 13512
rect 17368 13472 17374 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 18509 13515 18567 13521
rect 18509 13481 18521 13515
rect 18555 13512 18567 13515
rect 18598 13512 18604 13524
rect 18555 13484 18604 13512
rect 18555 13481 18567 13484
rect 18509 13475 18567 13481
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 12492 13416 12817 13444
rect 12492 13404 12498 13416
rect 12805 13413 12817 13416
rect 12851 13413 12863 13447
rect 12805 13407 12863 13413
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16623 13280 17233 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 17770 13308 17776 13320
rect 17267 13280 17776 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18414 13308 18420 13320
rect 18375 13280 18420 13308
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 13906 13240 13912 13252
rect 12483 13212 13912 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 15470 13240 15476 13252
rect 15431 13212 15476 13240
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 15689 13243 15747 13249
rect 15689 13209 15701 13243
rect 15735 13240 15747 13243
rect 16114 13240 16120 13252
rect 15735 13212 16120 13240
rect 15735 13209 15747 13212
rect 15689 13203 15747 13209
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 12618 13172 12624 13184
rect 12676 13181 12682 13184
rect 12676 13175 12705 13181
rect 12557 13144 12624 13172
rect 12618 13132 12624 13144
rect 12693 13172 12705 13175
rect 15378 13172 15384 13184
rect 12693 13144 15384 13172
rect 12693 13141 12705 13144
rect 12676 13135 12705 13141
rect 12676 13132 12682 13135
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 16666 13172 16672 13184
rect 16627 13144 16672 13172
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 27614 12968 27620 12980
rect 1627 12940 27620 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 11992 12696 12020 12795
rect 14182 12792 14188 12844
rect 14240 12792 14246 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15286 12832 15292 12844
rect 15243 12804 15292 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15436 12804 15481 12832
rect 15436 12792 15442 12804
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12618 12764 12624 12776
rect 12115 12736 12624 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12912 12736 13093 12764
rect 12345 12699 12403 12705
rect 11992 12668 12112 12696
rect 12084 12628 12112 12668
rect 12345 12665 12357 12699
rect 12391 12696 12403 12699
rect 12912 12696 12940 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 12391 12668 12940 12696
rect 12391 12665 12403 12668
rect 12345 12659 12403 12665
rect 14550 12628 14556 12640
rect 12084 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12628 14614 12640
rect 15010 12628 15016 12640
rect 14608 12600 15016 12628
rect 14608 12588 14614 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 15194 12628 15200 12640
rect 15155 12600 15200 12628
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 47762 12628 47768 12640
rect 47723 12600 47768 12628
rect 47762 12588 47768 12600
rect 47820 12588 47826 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12424 12771 12427
rect 12802 12424 12808 12436
rect 12759 12396 12808 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 14182 12424 14188 12436
rect 14143 12396 14188 12424
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 16301 12359 16359 12365
rect 16301 12325 16313 12359
rect 16347 12356 16359 12359
rect 16347 12328 16896 12356
rect 16347 12325 16359 12328
rect 16301 12319 16359 12325
rect 12728 12260 14872 12288
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 12728 12229 12756 12260
rect 14844 12232 14872 12260
rect 15838 12248 15844 12300
rect 15896 12288 15902 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 15896 12260 16037 12288
rect 15896 12248 15902 12260
rect 16025 12257 16037 12260
rect 16071 12288 16083 12291
rect 16482 12288 16488 12300
rect 16071 12260 16488 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16724 12260 16773 12288
rect 16724 12248 16730 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 16868 12288 16896 12328
rect 17037 12291 17095 12297
rect 17037 12288 17049 12291
rect 16868 12260 17049 12288
rect 16761 12251 16819 12257
rect 17037 12257 17049 12260
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12288 46351 12291
rect 47762 12288 47768 12300
rect 46339 12260 47768 12288
rect 46339 12257 46351 12260
rect 46293 12251 46351 12257
rect 47762 12248 47768 12260
rect 47820 12248 47826 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12308 12192 12725 12220
rect 12308 12180 12314 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 12713 12183 12771 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14826 12220 14832 12232
rect 14787 12192 14832 12220
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 15746 12220 15752 12232
rect 15436 12192 15752 12220
rect 15436 12180 15442 12192
rect 15746 12180 15752 12192
rect 15804 12220 15810 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15804 12192 15945 12220
rect 15804 12180 15810 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 14918 12084 14924 12096
rect 14879 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15948 12084 15976 12183
rect 18046 12112 18052 12164
rect 18104 12112 18110 12164
rect 46477 12155 46535 12161
rect 46477 12121 46489 12155
rect 46523 12152 46535 12155
rect 47670 12152 47676 12164
rect 46523 12124 47676 12152
rect 46523 12121 46535 12124
rect 46477 12115 46535 12121
rect 47670 12112 47676 12124
rect 47728 12112 47734 12164
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 15948 12056 18521 12084
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11880 18015 11883
rect 18046 11880 18052 11892
rect 18003 11852 18052 11880
rect 18003 11849 18015 11852
rect 17957 11843 18015 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 47670 11880 47676 11892
rect 47631 11852 47676 11880
rect 47670 11840 47676 11852
rect 47728 11840 47734 11892
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 15565 11815 15623 11821
rect 15565 11812 15577 11815
rect 15528 11784 15577 11812
rect 15528 11772 15534 11784
rect 15565 11781 15577 11784
rect 15611 11812 15623 11815
rect 16574 11812 16580 11824
rect 15611 11784 16580 11812
rect 15611 11781 15623 11784
rect 15565 11775 15623 11781
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 12250 11744 12256 11756
rect 12211 11716 12256 11744
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12676 11716 12817 11744
rect 12676 11704 12682 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 14090 11744 14096 11756
rect 13771 11716 14096 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13004 11676 13032 11707
rect 14090 11704 14096 11716
rect 14148 11744 14154 11756
rect 14148 11716 15148 11744
rect 14148 11704 14154 11716
rect 15010 11676 15016 11688
rect 13004 11648 15016 11676
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15120 11676 15148 11716
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 15436 11716 15761 11744
rect 15436 11704 15442 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15838 11704 15844 11756
rect 15896 11744 15902 11756
rect 16669 11747 16727 11753
rect 15896 11716 15941 11744
rect 15896 11704 15902 11716
rect 16669 11713 16681 11747
rect 16715 11744 16727 11747
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 16715 11716 17877 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 17865 11713 17877 11716
rect 17911 11744 17923 11747
rect 18414 11744 18420 11756
rect 17911 11716 18420 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 16684 11676 16712 11707
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 25958 11744 25964 11756
rect 25648 11716 25964 11744
rect 25648 11704 25654 11716
rect 25958 11704 25964 11716
rect 26016 11744 26022 11756
rect 46753 11747 46811 11753
rect 46753 11744 46765 11747
rect 26016 11716 46765 11744
rect 26016 11704 26022 11716
rect 46753 11713 46765 11716
rect 46799 11713 46811 11747
rect 46753 11707 46811 11713
rect 47581 11747 47639 11753
rect 47581 11713 47593 11747
rect 47627 11713 47639 11747
rect 47581 11707 47639 11713
rect 15120 11648 16712 11676
rect 28626 11636 28632 11688
rect 28684 11676 28690 11688
rect 47596 11676 47624 11707
rect 28684 11648 47624 11676
rect 28684 11636 28690 11648
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15565 11611 15623 11617
rect 15565 11608 15577 11611
rect 15344 11580 15577 11608
rect 15344 11568 15350 11580
rect 15565 11577 15577 11580
rect 15611 11577 15623 11611
rect 15565 11571 15623 11577
rect 12250 11540 12256 11552
rect 12211 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 16758 11540 16764 11552
rect 16719 11512 16764 11540
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 46474 11500 46480 11552
rect 46532 11540 46538 11552
rect 46845 11543 46903 11549
rect 46845 11540 46857 11543
rect 46532 11512 46857 11540
rect 46532 11500 46538 11512
rect 46845 11509 46857 11512
rect 46891 11509 46903 11543
rect 46845 11503 46903 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 12161 11203 12219 11209
rect 12161 11169 12173 11203
rect 12207 11200 12219 11203
rect 12894 11200 12900 11212
rect 12207 11172 12900 11200
rect 12207 11169 12219 11172
rect 12161 11163 12219 11169
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 14918 11200 14924 11212
rect 14879 11172 14924 11200
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15194 11200 15200 11212
rect 15155 11172 15200 11200
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16632 11172 16681 11200
rect 16632 11160 16638 11172
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 46474 11200 46480 11212
rect 46435 11172 46480 11200
rect 16669 11163 16727 11169
rect 46474 11160 46480 11172
rect 46532 11160 46538 11212
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 13906 11132 13912 11144
rect 12115 11104 13912 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 16758 11132 16764 11144
rect 16330 11104 16764 11132
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 46293 11135 46351 11141
rect 46293 11101 46305 11135
rect 46339 11101 46351 11135
rect 46293 11095 46351 11101
rect 46308 11064 46336 11095
rect 47762 11064 47768 11076
rect 46308 11036 47768 11064
rect 47762 11024 47768 11036
rect 47820 11024 47826 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 4798 10996 4804 11008
rect 3568 10968 4804 10996
rect 3568 10956 3574 10968
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12492 10968 12537 10996
rect 12492 10956 12498 10968
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 12434 10684 12440 10736
rect 12492 10724 12498 10736
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 12492 10696 12541 10724
rect 12492 10684 12498 10696
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 13814 10724 13820 10736
rect 13754 10696 13820 10724
rect 12529 10687 12587 10693
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 14700 10696 14933 10724
rect 14700 10684 14706 10696
rect 14921 10693 14933 10696
rect 14967 10693 14979 10727
rect 14921 10687 14979 10693
rect 12250 10656 12256 10668
rect 12211 10628 12256 10656
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 45189 10591 45247 10597
rect 45189 10557 45201 10591
rect 45235 10557 45247 10591
rect 45189 10551 45247 10557
rect 45373 10591 45431 10597
rect 45373 10557 45385 10591
rect 45419 10588 45431 10591
rect 46382 10588 46388 10600
rect 45419 10560 46388 10588
rect 45419 10557 45431 10560
rect 45373 10551 45431 10557
rect 15102 10520 15108 10532
rect 15063 10492 15108 10520
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 45204 10520 45232 10551
rect 46382 10548 46388 10560
rect 46440 10548 46446 10600
rect 46750 10588 46756 10600
rect 46711 10560 46756 10588
rect 46750 10548 46756 10560
rect 46808 10548 46814 10600
rect 45646 10520 45652 10532
rect 45204 10492 45652 10520
rect 45646 10480 45652 10492
rect 45704 10480 45710 10532
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13964 10424 14013 10452
rect 13964 10412 13970 10424
rect 14001 10421 14013 10424
rect 14047 10452 14059 10455
rect 14090 10452 14096 10464
rect 14047 10424 14096 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 15010 10112 15016 10124
rect 14971 10084 15016 10112
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 46293 10115 46351 10121
rect 46293 10081 46305 10115
rect 46339 10112 46351 10115
rect 47026 10112 47032 10124
rect 46339 10084 47032 10112
rect 46339 10081 46351 10084
rect 46293 10075 46351 10081
rect 47026 10072 47032 10084
rect 47084 10072 47090 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 13872 10016 14381 10044
rect 13872 10004 13878 10016
rect 14369 10013 14381 10016
rect 14415 10044 14427 10047
rect 14918 10044 14924 10056
rect 14415 10016 14924 10044
rect 14415 10013 14427 10016
rect 14369 10007 14427 10013
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15197 9979 15255 9985
rect 15197 9945 15209 9979
rect 15243 9976 15255 9979
rect 16758 9976 16764 9988
rect 15243 9948 16764 9976
rect 15243 9945 15255 9948
rect 15197 9939 15255 9945
rect 16758 9936 16764 9948
rect 16816 9936 16822 9988
rect 16853 9979 16911 9985
rect 16853 9945 16865 9979
rect 16899 9976 16911 9979
rect 25866 9976 25872 9988
rect 16899 9948 25872 9976
rect 16899 9945 16911 9948
rect 16853 9939 16911 9945
rect 25866 9936 25872 9948
rect 25924 9936 25930 9988
rect 46477 9979 46535 9985
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 14458 9908 14464 9920
rect 14419 9880 14464 9908
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 15378 9704 15384 9716
rect 14292 9676 14596 9704
rect 13998 9636 14004 9648
rect 13004 9608 14004 9636
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 13004 9577 13032 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 11848 9540 13001 9568
rect 11848 9528 11854 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9568 13691 9571
rect 13814 9568 13820 9580
rect 13679 9540 13820 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 14292 9577 14320 9676
rect 14458 9636 14464 9648
rect 14419 9608 14464 9636
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 14568 9636 14596 9676
rect 15028 9676 15384 9704
rect 15028 9636 15056 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 14568 9608 15056 9636
rect 15102 9596 15108 9648
rect 15160 9636 15166 9648
rect 16758 9636 16764 9648
rect 15160 9608 15700 9636
rect 16719 9608 16764 9636
rect 15160 9596 15166 9608
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9537 14335 9571
rect 15672 9568 15700 9608
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 47670 9636 47676 9648
rect 47631 9608 47676 9636
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 15672 9540 16681 9568
rect 14277 9531 14335 9537
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 47026 9568 47032 9580
rect 46987 9540 47032 9568
rect 16669 9531 16727 9537
rect 47026 9528 47032 9540
rect 47084 9528 47090 9580
rect 47486 9528 47492 9580
rect 47544 9568 47550 9580
rect 47581 9571 47639 9577
rect 47581 9568 47593 9571
rect 47544 9540 47593 9568
rect 47544 9528 47550 9540
rect 47581 9537 47593 9540
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 14737 9503 14795 9509
rect 14737 9469 14749 9503
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 14752 9432 14780 9463
rect 13688 9404 14780 9432
rect 13688 9392 13694 9404
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 13081 9367 13139 9373
rect 13081 9364 13093 9367
rect 11940 9336 13093 9364
rect 11940 9324 11946 9336
rect 13081 9333 13093 9336
rect 13127 9333 13139 9367
rect 13722 9364 13728 9376
rect 13683 9336 13728 9364
rect 13081 9327 13139 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 12066 9092 12072 9104
rect 11716 9064 12072 9092
rect 11716 9033 11744 9064
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 14108 9064 14780 9092
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 8993 11759 9027
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11701 8987 11759 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 13538 8888 13544 8900
rect 13499 8860 13544 8888
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 14108 8820 14136 9064
rect 14274 9024 14280 9036
rect 14235 8996 14280 9024
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 14752 9033 14780 9064
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 8993 14795 9027
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 14737 8987 14795 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 17954 9024 17960 9036
rect 17915 8996 17960 9024
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 46842 8984 46848 9036
rect 46900 9024 46906 9036
rect 47305 9027 47363 9033
rect 47305 9024 47317 9027
rect 46900 8996 47317 9024
rect 46900 8984 46906 8996
rect 47305 8993 47317 8996
rect 47351 8993 47363 9027
rect 47305 8987 47363 8993
rect 46382 8916 46388 8968
rect 46440 8956 46446 8968
rect 47581 8959 47639 8965
rect 47581 8956 47593 8959
rect 46440 8928 47593 8956
rect 46440 8916 46446 8928
rect 47581 8925 47593 8928
rect 47627 8925 47639 8959
rect 47581 8919 47639 8925
rect 14458 8888 14464 8900
rect 14419 8860 14464 8888
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 16758 8888 16764 8900
rect 16719 8860 16764 8888
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 3844 8792 14136 8820
rect 3844 8780 3850 8792
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 14277 8551 14335 8557
rect 14277 8548 14289 8551
rect 13780 8520 14289 8548
rect 13780 8508 13786 8520
rect 14277 8517 14289 8520
rect 14323 8517 14335 8551
rect 47762 8548 47768 8560
rect 47723 8520 47768 8548
rect 14277 8511 14335 8517
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 14090 8480 14096 8492
rect 14051 8452 14096 8480
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 11882 8412 11888 8424
rect 11843 8384 11888 8412
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 14826 8412 14832 8424
rect 14787 8384 14832 8412
rect 12437 8375 12495 8381
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 12452 8276 12480 8375
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 42702 8372 42708 8424
rect 42760 8412 42766 8424
rect 46934 8412 46940 8424
rect 42760 8384 46940 8412
rect 42760 8372 42766 8384
rect 46934 8372 46940 8384
rect 46992 8372 46998 8424
rect 24762 8304 24768 8356
rect 24820 8344 24826 8356
rect 47949 8347 48007 8353
rect 47949 8344 47961 8347
rect 24820 8316 47961 8344
rect 24820 8304 24826 8316
rect 47949 8313 47961 8316
rect 47995 8313 48007 8347
rect 47949 8307 48007 8313
rect 4120 8248 12480 8276
rect 4120 8236 4126 8248
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 45554 8276 45560 8288
rect 13596 8248 45560 8276
rect 13596 8236 13602 8248
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 11882 8072 11888 8084
rect 11839 8044 11888 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14516 8044 14565 8072
rect 14516 8032 14522 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 16758 8072 16764 8084
rect 15243 8044 16764 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 46293 7939 46351 7945
rect 46293 7905 46305 7939
rect 46339 7936 46351 7939
rect 46566 7936 46572 7948
rect 46339 7908 46572 7936
rect 46339 7905 46351 7908
rect 46293 7899 46351 7905
rect 46566 7896 46572 7908
rect 46624 7896 46630 7948
rect 46658 7896 46664 7948
rect 46716 7936 46722 7948
rect 46753 7939 46811 7945
rect 46753 7936 46765 7939
rect 46716 7908 46765 7936
rect 46716 7896 46722 7908
rect 46753 7905 46765 7908
rect 46799 7905 46811 7939
rect 46753 7899 46811 7905
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 10468 7840 11713 7868
rect 10468 7828 10474 7840
rect 11701 7837 11713 7840
rect 11747 7868 11759 7871
rect 11790 7868 11796 7880
rect 11747 7840 11796 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 13872 7840 14473 7868
rect 13872 7828 13878 7840
rect 14461 7837 14473 7840
rect 14507 7868 14519 7871
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14507 7840 15117 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 46477 7803 46535 7809
rect 46477 7769 46489 7803
rect 46523 7800 46535 7803
rect 47486 7800 47492 7812
rect 46523 7772 47492 7800
rect 46523 7769 46535 7772
rect 46477 7763 46535 7769
rect 47486 7760 47492 7772
rect 47544 7760 47550 7812
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 1670 7420 1676 7472
rect 1728 7460 1734 7472
rect 45005 7463 45063 7469
rect 45005 7460 45017 7463
rect 1728 7432 45017 7460
rect 1728 7420 1734 7432
rect 45005 7429 45017 7432
rect 45051 7429 45063 7463
rect 45005 7423 45063 7429
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 44913 7327 44971 7333
rect 44913 7293 44925 7327
rect 44959 7293 44971 7327
rect 45186 7324 45192 7336
rect 45147 7296 45192 7324
rect 44913 7287 44971 7293
rect 44928 7256 44956 7287
rect 45186 7284 45192 7296
rect 45244 7284 45250 7336
rect 47949 7259 48007 7265
rect 47949 7256 47961 7259
rect 44928 7228 47961 7256
rect 47949 7225 47961 7228
rect 47995 7225 48007 7259
rect 47949 7219 48007 7225
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 17954 6848 17960 6860
rect 4120 6820 17960 6848
rect 4120 6808 4126 6820
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47486 6808 47492 6860
rect 47544 6848 47550 6860
rect 47581 6851 47639 6857
rect 47581 6848 47593 6851
rect 47544 6820 47593 6848
rect 47544 6808 47550 6820
rect 47581 6817 47593 6820
rect 47627 6817 47639 6851
rect 47581 6811 47639 6817
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 48130 6304 48136 6316
rect 48091 6276 48136 6304
rect 48130 6264 48136 6276
rect 48188 6264 48194 6316
rect 14366 6128 14372 6180
rect 14424 6168 14430 6180
rect 32214 6168 32220 6180
rect 14424 6140 32220 6168
rect 14424 6128 14430 6140
rect 32214 6128 32220 6140
rect 32272 6128 32278 6180
rect 47946 6100 47952 6112
rect 47907 6072 47952 6100
rect 47946 6060 47952 6072
rect 48004 6060 48010 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 46842 5720 46848 5772
rect 46900 5760 46906 5772
rect 47305 5763 47363 5769
rect 47305 5760 47317 5763
rect 46900 5732 47317 5760
rect 46900 5720 46906 5732
rect 47305 5729 47317 5732
rect 47351 5729 47363 5763
rect 47305 5723 47363 5729
rect 46198 5652 46204 5704
rect 46256 5692 46262 5704
rect 47581 5695 47639 5701
rect 47581 5692 47593 5695
rect 46256 5664 47593 5692
rect 46256 5652 46262 5664
rect 47581 5661 47593 5664
rect 47627 5661 47639 5695
rect 47581 5655 47639 5661
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 45649 5287 45707 5293
rect 45649 5253 45661 5287
rect 45695 5284 45707 5287
rect 47946 5284 47952 5296
rect 45695 5256 47952 5284
rect 45695 5253 45707 5256
rect 45649 5247 45707 5253
rect 47946 5244 47952 5256
rect 48004 5244 48010 5296
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 18138 5216 18144 5228
rect 16715 5188 18144 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 20070 5216 20076 5228
rect 20031 5188 20076 5216
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5216 20775 5219
rect 21358 5216 21364 5228
rect 20763 5188 21364 5216
rect 20763 5185 20775 5188
rect 20717 5179 20775 5185
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 47854 5216 47860 5228
rect 47815 5188 47860 5216
rect 47854 5176 47860 5188
rect 47912 5176 47918 5228
rect 45557 5151 45615 5157
rect 45557 5117 45569 5151
rect 45603 5148 45615 5151
rect 45646 5148 45652 5160
rect 45603 5120 45652 5148
rect 45603 5117 45615 5120
rect 45557 5111 45615 5117
rect 45646 5108 45652 5120
rect 45704 5108 45710 5160
rect 45833 5151 45891 5157
rect 45833 5117 45845 5151
rect 45879 5117 45891 5151
rect 45833 5111 45891 5117
rect 45186 5040 45192 5092
rect 45244 5080 45250 5092
rect 45848 5080 45876 5111
rect 45244 5052 45876 5080
rect 45244 5040 45250 5052
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 17586 5012 17592 5024
rect 16807 4984 17592 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 20165 5015 20223 5021
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20714 5012 20720 5024
rect 20211 4984 20720 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 20809 5015 20867 5021
rect 20809 4981 20821 5015
rect 20855 5012 20867 5015
rect 21910 5012 21916 5024
rect 20855 4984 21916 5012
rect 20855 4981 20867 4984
rect 20809 4975 20867 4981
rect 21910 4972 21916 4984
rect 21968 4972 21974 5024
rect 32766 4972 32772 5024
rect 32824 5012 32830 5024
rect 48041 5015 48099 5021
rect 48041 5012 48053 5015
rect 32824 4984 48053 5012
rect 32824 4972 32830 4984
rect 48041 4981 48053 4984
rect 48087 4981 48099 5015
rect 48041 4975 48099 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 20070 4768 20076 4820
rect 20128 4808 20134 4820
rect 20717 4811 20775 4817
rect 20717 4808 20729 4811
rect 20128 4780 20729 4808
rect 20128 4768 20134 4780
rect 20717 4777 20729 4780
rect 20763 4777 20775 4811
rect 21358 4808 21364 4820
rect 21319 4780 21364 4808
rect 20717 4771 20775 4777
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 31478 4768 31484 4820
rect 31536 4808 31542 4820
rect 45094 4808 45100 4820
rect 31536 4780 45100 4808
rect 31536 4768 31542 4780
rect 45094 4768 45100 4780
rect 45152 4768 45158 4820
rect 45830 4768 45836 4820
rect 45888 4808 45894 4820
rect 45888 4780 46336 4808
rect 45888 4768 45894 4780
rect 46308 4684 46336 4780
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 6972 4644 15301 4672
rect 6972 4632 6978 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 20898 4672 20904 4684
rect 15289 4635 15347 4641
rect 19996 4644 20904 4672
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9456 4576 9597 4604
rect 9456 4564 9462 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 9585 4567 9643 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4604 19395 4607
rect 19886 4604 19892 4616
rect 19383 4576 19892 4604
rect 19383 4573 19395 4576
rect 19337 4567 19395 4573
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 19996 4613 20024 4644
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 45646 4632 45652 4684
rect 45704 4672 45710 4684
rect 45833 4675 45891 4681
rect 45833 4672 45845 4675
rect 45704 4644 45845 4672
rect 45704 4632 45710 4644
rect 45833 4641 45845 4644
rect 45879 4641 45891 4675
rect 46290 4672 46296 4684
rect 46251 4644 46296 4672
rect 45833 4635 45891 4641
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 19981 4607 20039 4613
rect 19981 4573 19993 4607
rect 20027 4573 20039 4607
rect 19981 4567 20039 4573
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20119 4576 20637 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20625 4573 20637 4576
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 20772 4576 21281 4604
rect 20772 4564 20778 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 21910 4604 21916 4616
rect 21871 4576 21916 4604
rect 21269 4567 21327 4573
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 42886 4604 42892 4616
rect 42847 4576 42892 4604
rect 42886 4564 42892 4576
rect 42944 4564 42950 4616
rect 45186 4564 45192 4616
rect 45244 4604 45250 4616
rect 45373 4607 45431 4613
rect 45373 4604 45385 4607
rect 45244 4576 45385 4604
rect 45244 4564 45250 4576
rect 45373 4573 45385 4576
rect 45419 4573 45431 4607
rect 45373 4567 45431 4573
rect 15473 4539 15531 4545
rect 15473 4505 15485 4539
rect 15519 4536 15531 4539
rect 15562 4536 15568 4548
rect 15519 4508 15568 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 17129 4539 17187 4545
rect 17129 4505 17141 4539
rect 17175 4536 17187 4539
rect 43990 4536 43996 4548
rect 17175 4508 43996 4536
rect 17175 4505 17187 4508
rect 17129 4499 17187 4505
rect 43990 4496 43996 4508
rect 44048 4496 44054 4548
rect 46014 4536 46020 4548
rect 45975 4508 46020 4536
rect 46014 4496 46020 4508
rect 46072 4496 46078 4548
rect 17034 4428 17040 4480
rect 17092 4468 17098 4480
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17092 4440 17693 4468
rect 17092 4428 17098 4440
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 17681 4431 17739 4437
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4468 19487 4471
rect 20714 4468 20720 4480
rect 19475 4440 20720 4468
rect 19475 4437 19487 4440
rect 19429 4431 19487 4437
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 23014 4468 23020 4480
rect 22051 4440 23020 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 18230 4264 18236 4276
rect 11572 4236 18236 4264
rect 11572 4224 11578 4236
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 41322 4224 41328 4276
rect 41380 4264 41386 4276
rect 41380 4236 43300 4264
rect 41380 4224 41386 4236
rect 16666 4196 16672 4208
rect 15856 4168 16672 4196
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4097 9459 4131
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 9401 4091 9459 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3142 4060 3148 4072
rect 2363 4032 3148 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2148 3992 2176 4023
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 7098 4060 7104 4072
rect 3292 4032 3337 4060
rect 7059 4032 7104 4060
rect 3292 4020 3298 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 8202 4060 8208 4072
rect 7331 4032 8208 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4029 8355 4063
rect 9416 4060 9444 4091
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 13725 4131 13783 4137
rect 11572 4100 11617 4128
rect 11572 4088 11578 4100
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 15856 4128 15884 4168
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 42702 4196 42708 4208
rect 22756 4168 23244 4196
rect 13771 4100 15884 4128
rect 15933 4131 15991 4137
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 15933 4097 15945 4131
rect 15979 4128 15991 4131
rect 16850 4128 16856 4140
rect 15979 4100 16856 4128
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 17034 4128 17040 4140
rect 16995 4100 17040 4128
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4128 17739 4131
rect 17770 4128 17776 4140
rect 17727 4100 17776 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 18506 4128 18512 4140
rect 18371 4100 18512 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19334 4128 19340 4140
rect 19015 4100 19340 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4097 19671 4131
rect 20806 4128 20812 4140
rect 20767 4100 20812 4128
rect 19613 4091 19671 4097
rect 15654 4060 15660 4072
rect 9416 4032 15660 4060
rect 8297 4023 8355 4029
rect 3878 3992 3884 4004
rect 2148 3964 3884 3992
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 8312 3992 8340 4023
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 19628 4060 19656 4091
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 22756 4128 22784 4168
rect 22235 4100 22784 4128
rect 22833 4131 22891 4137
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22833 4097 22845 4131
rect 22879 4128 22891 4131
rect 23106 4128 23112 4140
rect 22879 4100 23112 4128
rect 22879 4097 22891 4100
rect 22833 4091 22891 4097
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23216 4128 23244 4168
rect 42628 4168 42708 4196
rect 25590 4128 25596 4140
rect 23216 4100 25596 4128
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 25685 4131 25743 4137
rect 25685 4097 25697 4131
rect 25731 4128 25743 4131
rect 25774 4128 25780 4140
rect 25731 4100 25780 4128
rect 25731 4097 25743 4100
rect 25685 4091 25743 4097
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 30926 4088 30932 4140
rect 30984 4128 30990 4140
rect 33137 4131 33195 4137
rect 33137 4128 33149 4131
rect 30984 4100 33149 4128
rect 30984 4088 30990 4100
rect 33137 4097 33149 4100
rect 33183 4097 33195 4131
rect 39758 4128 39764 4140
rect 39719 4100 39764 4128
rect 33137 4091 33195 4097
rect 39758 4088 39764 4100
rect 39816 4088 39822 4140
rect 42628 4137 42656 4168
rect 42702 4156 42708 4168
rect 42760 4156 42766 4208
rect 43272 4196 43300 4236
rect 45646 4196 45652 4208
rect 43272 4168 45652 4196
rect 43272 4137 43300 4168
rect 45646 4156 45652 4168
rect 45704 4156 45710 4208
rect 42613 4131 42671 4137
rect 42613 4097 42625 4131
rect 42659 4097 42671 4131
rect 42613 4091 42671 4097
rect 43257 4131 43315 4137
rect 43257 4097 43269 4131
rect 43303 4097 43315 4131
rect 46106 4128 46112 4140
rect 46067 4100 46112 4128
rect 43257 4091 43315 4097
rect 46106 4088 46112 4100
rect 46164 4088 46170 4140
rect 46658 4088 46664 4140
rect 46716 4128 46722 4140
rect 46753 4131 46811 4137
rect 46753 4128 46765 4131
rect 46716 4100 46765 4128
rect 46716 4088 46722 4100
rect 46753 4097 46765 4100
rect 46799 4097 46811 4131
rect 46753 4091 46811 4097
rect 46842 4088 46848 4140
rect 46900 4128 46906 4140
rect 47857 4131 47915 4137
rect 47857 4128 47869 4131
rect 46900 4100 47869 4128
rect 46900 4088 46906 4100
rect 47857 4097 47869 4100
rect 47903 4097 47915 4131
rect 47857 4091 47915 4097
rect 29549 4063 29607 4069
rect 29549 4060 29561 4063
rect 19300 4032 19656 4060
rect 22066 4032 29561 4060
rect 19300 4020 19306 4032
rect 10042 3992 10048 4004
rect 7248 3964 8340 3992
rect 8404 3964 10048 3992
rect 7248 3952 7254 3964
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 8404 3924 8432 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 17218 3952 17224 4004
rect 17276 3992 17282 4004
rect 22066 3992 22094 4032
rect 29549 4029 29561 4032
rect 29595 4029 29607 4063
rect 29549 4023 29607 4029
rect 29733 4063 29791 4069
rect 29733 4029 29745 4063
rect 29779 4060 29791 4063
rect 30006 4060 30012 4072
rect 29779 4032 30012 4060
rect 29779 4029 29791 4032
rect 29733 4023 29791 4029
rect 30006 4020 30012 4032
rect 30064 4020 30070 4072
rect 31386 4060 31392 4072
rect 31347 4032 31392 4060
rect 31386 4020 31392 4032
rect 31444 4020 31450 4072
rect 36170 4020 36176 4072
rect 36228 4060 36234 4072
rect 43441 4063 43499 4069
rect 36228 4032 43208 4060
rect 36228 4020 36234 4032
rect 17276 3964 22094 3992
rect 17276 3952 17282 3964
rect 22738 3952 22744 4004
rect 22796 3992 22802 4004
rect 36538 3992 36544 4004
rect 22796 3964 36544 3992
rect 22796 3952 22802 3964
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 37826 3952 37832 4004
rect 37884 3992 37890 4004
rect 43180 3992 43208 4032
rect 43441 4029 43453 4063
rect 43487 4060 43499 4063
rect 43898 4060 43904 4072
rect 43487 4032 43904 4060
rect 43487 4029 43499 4032
rect 43441 4023 43499 4029
rect 43898 4020 43904 4032
rect 43956 4020 43962 4072
rect 43990 4020 43996 4072
rect 44048 4060 44054 4072
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 44048 4032 44189 4060
rect 44048 4020 44054 4032
rect 44177 4029 44189 4032
rect 44223 4029 44235 4063
rect 44177 4023 44235 4029
rect 46937 3995 46995 4001
rect 46937 3992 46949 3995
rect 37884 3964 42932 3992
rect 43180 3964 46949 3992
rect 37884 3952 37890 3964
rect 9490 3924 9496 3936
rect 4028 3896 8432 3924
rect 9451 3896 9496 3924
rect 4028 3884 4034 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 9640 3896 10517 3924
rect 9640 3884 9646 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 11698 3924 11704 3936
rect 11655 3896 11704 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 16025 3927 16083 3933
rect 16025 3893 16037 3927
rect 16071 3924 16083 3927
rect 16942 3924 16948 3936
rect 16071 3896 16948 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17129 3927 17187 3933
rect 17129 3893 17141 3927
rect 17175 3924 17187 3927
rect 17678 3924 17684 3936
rect 17175 3896 17684 3924
rect 17175 3893 17187 3896
rect 17129 3887 17187 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 18322 3924 18328 3936
rect 17819 3896 18328 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 19058 3924 19064 3936
rect 18472 3896 18517 3924
rect 19019 3896 19064 3924
rect 18472 3884 18478 3896
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 19705 3927 19763 3933
rect 19705 3924 19717 3927
rect 19484 3896 19717 3924
rect 19484 3884 19490 3896
rect 19705 3893 19717 3896
rect 19751 3893 19763 3927
rect 19705 3887 19763 3893
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20312 3896 20913 3924
rect 20312 3884 20318 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 20901 3887 20959 3893
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 22925 3927 22983 3933
rect 22925 3893 22937 3927
rect 22971 3924 22983 3927
rect 23658 3924 23664 3936
rect 22971 3896 23664 3924
rect 22971 3893 22983 3896
rect 22925 3887 22983 3893
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 25777 3927 25835 3933
rect 25777 3924 25789 3927
rect 25372 3896 25789 3924
rect 25372 3884 25378 3896
rect 25777 3893 25789 3896
rect 25823 3893 25835 3927
rect 25777 3887 25835 3893
rect 25866 3884 25872 3936
rect 25924 3924 25930 3936
rect 30834 3924 30840 3936
rect 25924 3896 30840 3924
rect 25924 3884 25930 3896
rect 30834 3884 30840 3896
rect 30892 3884 30898 3936
rect 33226 3924 33232 3936
rect 33187 3896 33232 3924
rect 33226 3884 33232 3896
rect 33284 3884 33290 3936
rect 39850 3924 39856 3936
rect 39811 3896 39856 3924
rect 39850 3884 39856 3896
rect 39908 3884 39914 3936
rect 42705 3927 42763 3933
rect 42705 3893 42717 3927
rect 42751 3924 42763 3927
rect 42794 3924 42800 3936
rect 42751 3896 42800 3924
rect 42751 3893 42763 3896
rect 42705 3887 42763 3893
rect 42794 3884 42800 3896
rect 42852 3884 42858 3936
rect 42904 3924 42932 3964
rect 46937 3961 46949 3964
rect 46983 3961 46995 3995
rect 46937 3955 46995 3961
rect 43530 3924 43536 3936
rect 42904 3896 43536 3924
rect 43530 3884 43536 3896
rect 43588 3884 43594 3936
rect 46201 3927 46259 3933
rect 46201 3893 46213 3927
rect 46247 3924 46259 3927
rect 46474 3924 46480 3936
rect 46247 3896 46480 3924
rect 46247 3893 46259 3896
rect 46201 3887 46259 3893
rect 46474 3884 46480 3896
rect 46532 3884 46538 3936
rect 48038 3924 48044 3936
rect 47999 3896 48044 3924
rect 48038 3884 48044 3896
rect 48096 3884 48102 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3936 3692 3985 3720
rect 3936 3680 3942 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 8202 3720 8208 3732
rect 8163 3692 8208 3720
rect 3973 3683 4031 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8312 3692 9996 3720
rect 8312 3652 8340 3692
rect 5184 3624 8340 3652
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 5184 3525 5212 3624
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 9968 3652 9996 3692
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 17218 3720 17224 3732
rect 10100 3692 17224 3720
rect 10100 3680 10106 3692
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17770 3720 17776 3732
rect 17731 3692 17776 3720
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18417 3723 18475 3729
rect 18417 3689 18429 3723
rect 18463 3720 18475 3723
rect 18506 3720 18512 3732
rect 18463 3692 18512 3720
rect 18463 3689 18475 3692
rect 18417 3683 18475 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 33962 3720 33968 3732
rect 20220 3692 33968 3720
rect 20220 3680 20226 3692
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 36538 3680 36544 3732
rect 36596 3720 36602 3732
rect 41230 3720 41236 3732
rect 36596 3692 41236 3720
rect 36596 3680 36602 3692
rect 41230 3680 41236 3692
rect 41288 3680 41294 3732
rect 42610 3720 42616 3732
rect 41386 3692 42616 3720
rect 15102 3652 15108 3664
rect 9088 3624 9904 3652
rect 9968 3624 15108 3652
rect 9088 3612 9094 3624
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 9398 3584 9404 3596
rect 9359 3556 9404 3584
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9582 3584 9588 3596
rect 9543 3556 9588 3584
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9876 3593 9904 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 41386 3652 41414 3692
rect 42610 3680 42616 3692
rect 42668 3680 42674 3732
rect 42886 3652 42892 3664
rect 15212 3624 19380 3652
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 3099 3488 5181 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5810 3516 5816 3528
rect 5771 3488 5816 3516
rect 5169 3479 5227 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11572 3488 11897 3516
rect 11572 3476 11578 3488
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 5997 3451 6055 3457
rect 5997 3448 6009 3451
rect 5307 3420 6009 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 5997 3417 6009 3420
rect 6043 3417 6055 3451
rect 13630 3448 13636 3460
rect 5997 3411 6055 3417
rect 7116 3420 13636 3448
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2004 3352 2237 3380
rect 2004 3340 2010 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 7116 3380 7144 3420
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 4120 3352 7144 3380
rect 4120 3340 4126 3352
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 15212 3380 15240 3624
rect 15378 3584 15384 3596
rect 15339 3556 15384 3584
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3553 15899 3587
rect 15841 3547 15899 3553
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15856 3516 15884 3547
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 15856 3488 16313 3516
rect 15473 3479 15531 3485
rect 16301 3485 16313 3488
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 15488 3448 15516 3479
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16816 3488 16957 3516
rect 16816 3476 16822 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 17678 3516 17684 3528
rect 17639 3488 17684 3516
rect 16945 3479 17003 3485
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18472 3488 19257 3516
rect 18472 3476 18478 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19352 3516 19380 3624
rect 19628 3624 41414 3652
rect 42628 3624 42892 3652
rect 19628 3516 19656 3624
rect 20254 3584 20260 3596
rect 20215 3556 20260 3584
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 20346 3544 20352 3596
rect 20404 3584 20410 3596
rect 20533 3587 20591 3593
rect 20533 3584 20545 3587
rect 20404 3556 20545 3584
rect 20404 3544 20410 3556
rect 20533 3553 20545 3556
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 25314 3584 25320 3596
rect 20864 3556 23980 3584
rect 25275 3556 25320 3584
rect 20864 3544 20870 3556
rect 20070 3516 20076 3528
rect 19352 3488 19656 3516
rect 20031 3488 20076 3516
rect 19245 3479 19303 3485
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22152 3488 22569 3516
rect 22152 3476 22158 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 22557 3479 22615 3485
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23658 3516 23664 3528
rect 23164 3488 23209 3516
rect 23619 3488 23664 3516
rect 23164 3476 23170 3488
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 21082 3448 21088 3460
rect 15488 3420 21088 3448
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 21174 3408 21180 3460
rect 21232 3448 21238 3460
rect 23952 3448 23980 3556
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 25406 3544 25412 3596
rect 25464 3584 25470 3596
rect 25593 3587 25651 3593
rect 25593 3584 25605 3587
rect 25464 3556 25605 3584
rect 25464 3544 25470 3556
rect 25593 3553 25605 3556
rect 25639 3553 25651 3587
rect 25593 3547 25651 3553
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 42518 3584 42524 3596
rect 27580 3556 42524 3584
rect 27580 3544 27586 3556
rect 42518 3544 42524 3556
rect 42576 3544 42582 3596
rect 42628 3593 42656 3624
rect 42886 3612 42892 3624
rect 42944 3612 42950 3664
rect 45646 3612 45652 3664
rect 45704 3652 45710 3664
rect 47394 3652 47400 3664
rect 45704 3624 47400 3652
rect 45704 3612 45710 3624
rect 47394 3612 47400 3624
rect 47452 3612 47458 3664
rect 42613 3587 42671 3593
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 42794 3584 42800 3596
rect 42755 3556 42800 3584
rect 42613 3547 42671 3553
rect 42794 3544 42800 3556
rect 42852 3544 42858 3596
rect 43162 3584 43168 3596
rect 43123 3556 43168 3584
rect 43162 3544 43168 3556
rect 43220 3544 43226 3596
rect 45189 3587 45247 3593
rect 45189 3553 45201 3587
rect 45235 3584 45247 3587
rect 46474 3584 46480 3596
rect 45235 3556 45968 3584
rect 46435 3556 46480 3584
rect 45235 3553 45247 3556
rect 45189 3547 45247 3553
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3516 24731 3519
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 24719 3488 25145 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 25133 3485 25145 3488
rect 25179 3485 25191 3519
rect 25133 3479 25191 3485
rect 33042 3476 33048 3528
rect 33100 3516 33106 3528
rect 33321 3519 33379 3525
rect 33321 3516 33333 3519
rect 33100 3488 33333 3516
rect 33100 3476 33106 3488
rect 33321 3485 33333 3488
rect 33367 3485 33379 3519
rect 35986 3516 35992 3528
rect 35947 3488 35992 3516
rect 33321 3479 33379 3485
rect 35986 3476 35992 3488
rect 36044 3476 36050 3528
rect 37826 3516 37832 3528
rect 37787 3488 37832 3516
rect 37826 3476 37832 3488
rect 37884 3476 37890 3528
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40310 3516 40316 3528
rect 40271 3488 40316 3516
rect 40037 3479 40095 3485
rect 40310 3476 40316 3488
rect 40368 3476 40374 3528
rect 40402 3476 40408 3528
rect 40460 3516 40466 3528
rect 41322 3516 41328 3528
rect 40460 3488 41328 3516
rect 40460 3476 40466 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41506 3516 41512 3528
rect 41467 3488 41512 3516
rect 41506 3476 41512 3488
rect 41564 3476 41570 3528
rect 45646 3516 45652 3528
rect 45607 3488 45652 3516
rect 45646 3476 45652 3488
rect 45704 3476 45710 3528
rect 45940 3516 45968 3556
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 45940 3488 46305 3516
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 28626 3448 28632 3460
rect 21232 3420 23888 3448
rect 23952 3420 28632 3448
rect 21232 3408 21238 3420
rect 7340 3352 15240 3380
rect 16393 3383 16451 3389
rect 7340 3340 7346 3352
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 16666 3380 16672 3392
rect 16439 3352 16672 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17037 3383 17095 3389
rect 17037 3349 17049 3383
rect 17083 3380 17095 3383
rect 17310 3380 17316 3392
rect 17083 3352 17316 3380
rect 17083 3349 17095 3352
rect 17037 3343 17095 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 21266 3380 21272 3392
rect 19392 3352 21272 3380
rect 19392 3340 19398 3352
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 23750 3380 23756 3392
rect 23711 3352 23756 3380
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 23860 3380 23888 3420
rect 28626 3408 28632 3420
rect 28684 3408 28690 3460
rect 36170 3448 36176 3460
rect 36131 3420 36176 3448
rect 36170 3408 36176 3420
rect 36228 3408 36234 3460
rect 36446 3408 36452 3460
rect 36504 3448 36510 3460
rect 48038 3448 48044 3460
rect 36504 3420 40356 3448
rect 36504 3408 36510 3420
rect 30926 3380 30932 3392
rect 23860 3352 30932 3380
rect 30926 3340 30932 3352
rect 30984 3340 30990 3392
rect 31386 3340 31392 3392
rect 31444 3380 31450 3392
rect 36538 3380 36544 3392
rect 31444 3352 36544 3380
rect 31444 3340 31450 3352
rect 36538 3340 36544 3352
rect 36596 3340 36602 3392
rect 37734 3340 37740 3392
rect 37792 3380 37798 3392
rect 39209 3383 39267 3389
rect 39209 3380 39221 3383
rect 37792 3352 39221 3380
rect 37792 3340 37798 3352
rect 39209 3349 39221 3352
rect 39255 3349 39267 3383
rect 40328 3380 40356 3420
rect 41386 3420 48044 3448
rect 41386 3380 41414 3420
rect 48038 3408 48044 3420
rect 48096 3408 48102 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 40328 3352 41414 3380
rect 41969 3383 42027 3389
rect 39209 3343 39267 3349
rect 41969 3349 41981 3383
rect 42015 3380 42027 3383
rect 42426 3380 42432 3392
rect 42015 3352 42432 3380
rect 42015 3349 42027 3352
rect 41969 3343 42027 3349
rect 42426 3340 42432 3352
rect 42484 3340 42490 3392
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 7282 3176 7288 3188
rect 3936 3148 7288 3176
rect 3936 3136 3942 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 16758 3176 16764 3188
rect 16719 3148 16764 3176
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 16908 3148 17417 3176
rect 16908 3136 16914 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 19153 3179 19211 3185
rect 19153 3145 19165 3179
rect 19199 3176 19211 3179
rect 19242 3176 19248 3188
rect 19199 3148 19248 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 20898 3176 20904 3188
rect 20855 3148 20904 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21082 3136 21088 3188
rect 21140 3176 21146 3188
rect 30190 3176 30196 3188
rect 21140 3148 30196 3176
rect 21140 3136 21146 3148
rect 30190 3136 30196 3148
rect 30248 3136 30254 3188
rect 36446 3176 36452 3188
rect 30300 3148 36452 3176
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 8205 3111 8263 3117
rect 8205 3077 8217 3111
rect 8251 3108 8263 3111
rect 9490 3108 9496 3120
rect 8251 3080 9496 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 16390 3068 16396 3120
rect 16448 3108 16454 3120
rect 21174 3108 21180 3120
rect 16448 3080 21180 3108
rect 16448 3068 16454 3080
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 22278 3108 22284 3120
rect 22239 3080 22284 3108
rect 22278 3068 22284 3080
rect 22336 3068 22342 3120
rect 26510 3108 26516 3120
rect 23492 3080 26516 3108
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5868 3012 6561 3040
rect 5868 3000 5874 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7156 3012 7389 3040
rect 7156 3000 7162 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 7377 3003 7435 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17954 3040 17960 3052
rect 17915 3012 17960 3040
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 19058 3040 19064 3052
rect 19019 3012 19064 3040
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20128 3012 20269 3040
rect 20128 3000 20134 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20257 3003 20315 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 22094 3040 22100 3052
rect 22055 3012 22100 3040
rect 22094 3000 22100 3012
rect 22152 3000 22158 3052
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 2225 2935 2283 2941
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8496 2904 8524 2935
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11020 2944 11989 2972
rect 11020 2932 11026 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 20162 2972 20168 2984
rect 17460 2944 20168 2972
rect 17460 2932 17466 2944
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 7800 2876 8524 2904
rect 7800 2864 7806 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 23492 2904 23520 3080
rect 26510 3068 26516 3080
rect 26568 3068 26574 3120
rect 28902 3108 28908 3120
rect 28552 3080 28908 3108
rect 28552 3049 28580 3080
rect 28902 3068 28908 3080
rect 28960 3068 28966 3120
rect 28537 3043 28595 3049
rect 28537 3009 28549 3043
rect 28583 3009 28595 3043
rect 28537 3003 28595 3009
rect 24394 2972 24400 2984
rect 24355 2944 24400 2972
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2941 24639 2975
rect 26142 2972 26148 2984
rect 26103 2944 26148 2972
rect 24581 2935 24639 2941
rect 15160 2876 23520 2904
rect 24596 2904 24624 2935
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 28721 2975 28779 2981
rect 28721 2941 28733 2975
rect 28767 2972 28779 2975
rect 30300 2972 30328 3148
rect 36446 3136 36452 3148
rect 36504 3136 36510 3188
rect 36538 3136 36544 3188
rect 36596 3176 36602 3188
rect 46290 3176 46296 3188
rect 36596 3148 46296 3176
rect 36596 3136 36602 3148
rect 46290 3136 46296 3148
rect 46348 3136 46354 3188
rect 33226 3108 33232 3120
rect 33187 3080 33232 3108
rect 33226 3068 33232 3080
rect 33284 3068 33290 3120
rect 39025 3111 39083 3117
rect 39025 3077 39037 3111
rect 39071 3108 39083 3111
rect 39758 3108 39764 3120
rect 39071 3080 39764 3108
rect 39071 3077 39083 3080
rect 39025 3071 39083 3077
rect 39758 3068 39764 3080
rect 39816 3068 39822 3120
rect 41598 3068 41604 3120
rect 41656 3108 41662 3120
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 41656 3080 42625 3108
rect 41656 3068 41662 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 42613 3071 42671 3077
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 47762 3108 47768 3120
rect 47723 3080 47768 3108
rect 47762 3068 47768 3080
rect 47820 3068 47826 3120
rect 33042 3040 33048 3052
rect 33003 3012 33048 3040
rect 33042 3000 33048 3012
rect 33100 3000 33106 3052
rect 37734 3040 37740 3052
rect 37695 3012 37740 3040
rect 37734 3000 37740 3012
rect 37792 3000 37798 3052
rect 37829 3043 37887 3049
rect 37829 3009 37841 3043
rect 37875 3040 37887 3043
rect 39485 3043 39543 3049
rect 39485 3040 39497 3043
rect 37875 3012 39497 3040
rect 37875 3009 37887 3012
rect 37829 3003 37887 3009
rect 39485 3009 39497 3012
rect 39531 3009 39543 3043
rect 39485 3003 39543 3009
rect 41230 3000 41236 3052
rect 41288 3040 41294 3052
rect 42426 3040 42432 3052
rect 41288 3012 41828 3040
rect 42387 3012 42432 3040
rect 41288 3000 41294 3012
rect 28767 2944 30328 2972
rect 28767 2941 28779 2944
rect 28721 2935 28779 2941
rect 30374 2932 30380 2984
rect 30432 2972 30438 2984
rect 33502 2972 33508 2984
rect 30432 2944 30477 2972
rect 33463 2944 33508 2972
rect 30432 2932 30438 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 35986 2932 35992 2984
rect 36044 2972 36050 2984
rect 38381 2975 38439 2981
rect 38381 2972 38393 2975
rect 36044 2944 38393 2972
rect 36044 2932 36050 2944
rect 38381 2941 38393 2944
rect 38427 2941 38439 2975
rect 38381 2935 38439 2941
rect 38565 2975 38623 2981
rect 38565 2941 38577 2975
rect 38611 2972 38623 2975
rect 39669 2975 39727 2981
rect 39669 2972 39681 2975
rect 38611 2944 39681 2972
rect 38611 2941 38623 2944
rect 38565 2935 38623 2941
rect 39669 2941 39681 2944
rect 39715 2972 39727 2975
rect 40310 2972 40316 2984
rect 39715 2944 40316 2972
rect 39715 2941 39727 2944
rect 39669 2935 39727 2941
rect 35710 2904 35716 2916
rect 24596 2876 35716 2904
rect 15160 2864 15166 2876
rect 35710 2864 35716 2876
rect 35768 2864 35774 2916
rect 38396 2904 38424 2935
rect 40310 2932 40316 2944
rect 40368 2932 40374 2984
rect 41322 2972 41328 2984
rect 41283 2944 41328 2972
rect 41322 2932 41328 2944
rect 41380 2932 41386 2984
rect 40402 2904 40408 2916
rect 38396 2876 40408 2904
rect 40402 2864 40408 2876
rect 40460 2864 40466 2916
rect 41340 2904 41368 2932
rect 40512 2876 41368 2904
rect 41800 2904 41828 3012
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 44266 2972 44272 2984
rect 44179 2944 44272 2972
rect 44266 2932 44272 2944
rect 44324 2972 44330 2984
rect 46566 2972 46572 2984
rect 44324 2944 46572 2972
rect 44324 2932 44330 2944
rect 46566 2932 46572 2944
rect 46624 2932 46630 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 47949 2907 48007 2913
rect 47949 2904 47961 2907
rect 41800 2876 47961 2904
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 28258 2836 28264 2848
rect 18288 2808 28264 2836
rect 18288 2796 18294 2808
rect 28258 2796 28264 2808
rect 28316 2796 28322 2848
rect 30374 2796 30380 2848
rect 30432 2836 30438 2848
rect 40512 2836 40540 2876
rect 47949 2873 47961 2876
rect 47995 2873 48007 2907
rect 47949 2867 48007 2873
rect 30432 2808 40540 2836
rect 30432 2796 30438 2808
rect 40586 2796 40592 2848
rect 40644 2836 40650 2848
rect 42886 2836 42892 2848
rect 40644 2808 42892 2836
rect 40644 2796 40650 2808
rect 42886 2796 42892 2808
rect 42944 2796 42950 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 17310 2632 17316 2644
rect 6886 2604 17316 2632
rect 2133 2567 2191 2573
rect 2133 2533 2145 2567
rect 2179 2564 2191 2567
rect 6886 2564 6914 2604
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17954 2632 17960 2644
rect 17543 2604 17960 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 19978 2632 19984 2644
rect 19751 2604 19984 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20438 2632 20444 2644
rect 20399 2604 20444 2632
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 21818 2592 21824 2644
rect 21876 2632 21882 2644
rect 21913 2635 21971 2641
rect 21913 2632 21925 2635
rect 21876 2604 21925 2632
rect 21876 2592 21882 2604
rect 21913 2601 21925 2604
rect 21959 2601 21971 2635
rect 21913 2595 21971 2601
rect 23661 2635 23719 2641
rect 23661 2601 23673 2635
rect 23707 2632 23719 2635
rect 24394 2632 24400 2644
rect 23707 2604 24400 2632
rect 23707 2601 23719 2604
rect 23661 2595 23719 2601
rect 24394 2592 24400 2604
rect 24452 2592 24458 2644
rect 24486 2592 24492 2644
rect 24544 2632 24550 2644
rect 24949 2635 25007 2641
rect 24949 2632 24961 2635
rect 24544 2604 24961 2632
rect 24544 2592 24550 2604
rect 24949 2601 24961 2604
rect 24995 2601 25007 2635
rect 30650 2632 30656 2644
rect 24949 2595 25007 2601
rect 26206 2604 30656 2632
rect 2179 2536 6914 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 8018 2524 8024 2576
rect 8076 2564 8082 2576
rect 8205 2567 8263 2573
rect 8205 2564 8217 2567
rect 8076 2536 8217 2564
rect 8076 2524 8082 2536
rect 8205 2533 8217 2536
rect 8251 2533 8263 2567
rect 8205 2527 8263 2533
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 24578 2564 24584 2576
rect 16899 2536 24584 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 24578 2524 24584 2536
rect 24636 2524 24642 2576
rect 15562 2496 15568 2508
rect 15523 2468 15568 2496
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 26206 2496 26234 2604
rect 30650 2592 30656 2604
rect 30708 2592 30714 2644
rect 35710 2632 35716 2644
rect 35671 2604 35716 2632
rect 35710 2592 35716 2604
rect 35768 2592 35774 2644
rect 35866 2604 36124 2632
rect 26421 2567 26479 2573
rect 26421 2533 26433 2567
rect 26467 2564 26479 2567
rect 28350 2564 28356 2576
rect 26467 2536 28356 2564
rect 26467 2533 26479 2536
rect 26421 2527 26479 2533
rect 28350 2524 28356 2536
rect 28408 2524 28414 2576
rect 28442 2524 28448 2576
rect 28500 2564 28506 2576
rect 35866 2564 35894 2604
rect 28500 2536 35894 2564
rect 36096 2564 36124 2604
rect 36170 2592 36176 2644
rect 36228 2632 36234 2644
rect 36265 2635 36323 2641
rect 36265 2632 36277 2635
rect 36228 2604 36277 2632
rect 36228 2592 36234 2604
rect 36265 2601 36277 2604
rect 36311 2601 36323 2635
rect 36265 2595 36323 2601
rect 39114 2592 39120 2644
rect 39172 2632 39178 2644
rect 39209 2635 39267 2641
rect 39209 2632 39221 2635
rect 39172 2604 39221 2632
rect 39172 2592 39178 2604
rect 39209 2601 39221 2604
rect 39255 2601 39267 2635
rect 39209 2595 39267 2601
rect 39298 2592 39304 2644
rect 39356 2632 39362 2644
rect 40405 2635 40463 2641
rect 40405 2632 40417 2635
rect 39356 2604 40417 2632
rect 39356 2592 39362 2604
rect 40405 2601 40417 2604
rect 40451 2601 40463 2635
rect 42978 2632 42984 2644
rect 42939 2604 42984 2632
rect 40405 2595 40463 2601
rect 42978 2592 42984 2604
rect 43036 2592 43042 2644
rect 47949 2567 48007 2573
rect 47949 2564 47961 2567
rect 36096 2536 47961 2564
rect 28500 2524 28506 2536
rect 47949 2533 47961 2536
rect 47995 2533 48007 2567
rect 47949 2527 48007 2533
rect 20272 2468 26234 2496
rect 27617 2499 27675 2505
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 17000 2400 17417 2428
rect 17000 2388 17006 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 18046 2428 18052 2440
rect 18007 2400 18052 2428
rect 17405 2391 17463 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19484 2400 19625 2428
rect 19484 2388 19490 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1360 2332 1869 2360
rect 1360 2320 1366 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2648 2332 2789 2360
rect 2648 2320 2654 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 20272 2360 20300 2468
rect 27617 2465 27629 2499
rect 27663 2496 27675 2499
rect 28994 2496 29000 2508
rect 27663 2468 29000 2496
rect 27663 2465 27675 2468
rect 27617 2459 27675 2465
rect 28994 2456 29000 2468
rect 29052 2456 29058 2508
rect 30006 2496 30012 2508
rect 29967 2468 30012 2496
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 32398 2456 32404 2508
rect 32456 2496 32462 2508
rect 38381 2499 38439 2505
rect 38381 2496 38393 2499
rect 32456 2468 38393 2496
rect 32456 2456 32462 2468
rect 38381 2465 38393 2468
rect 38427 2465 38439 2499
rect 38381 2459 38439 2465
rect 41325 2499 41383 2505
rect 41325 2465 41337 2499
rect 41371 2496 41383 2499
rect 41506 2496 41512 2508
rect 41371 2468 41512 2496
rect 41371 2465 41383 2468
rect 41325 2459 41383 2465
rect 41506 2456 41512 2468
rect 41564 2456 41570 2508
rect 43898 2496 43904 2508
rect 43859 2468 43904 2496
rect 43898 2456 43904 2468
rect 43956 2456 43962 2508
rect 46201 2499 46259 2505
rect 46201 2465 46213 2499
rect 46247 2496 46259 2499
rect 47026 2496 47032 2508
rect 46247 2468 47032 2496
rect 46247 2465 46259 2468
rect 46201 2459 46259 2465
rect 47026 2456 47032 2468
rect 47084 2456 47090 2508
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 21315 2400 21925 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 21913 2397 21925 2400
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2428 23075 2431
rect 23750 2428 23756 2440
rect 23063 2400 23756 2428
rect 23063 2397 23075 2400
rect 23017 2391 23075 2397
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 9815 2332 20300 2360
rect 20349 2363 20407 2369
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 20622 2360 20628 2372
rect 20395 2332 20628 2360
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21131 2332 21956 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21928 2304 21956 2332
rect 23198 2320 23204 2372
rect 23256 2360 23262 2372
rect 23860 2360 23888 2391
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 36136 2400 36461 2428
rect 36136 2388 36142 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 39117 2431 39175 2437
rect 39117 2397 39129 2431
rect 39163 2428 39175 2431
rect 39850 2428 39856 2440
rect 39163 2400 39856 2428
rect 39163 2397 39175 2400
rect 39117 2391 39175 2397
rect 39850 2388 39856 2400
rect 39908 2388 39914 2440
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41230 2428 41236 2440
rect 41095 2400 41236 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 42886 2428 42892 2440
rect 42847 2400 42892 2428
rect 42886 2388 42892 2400
rect 42944 2388 42950 2440
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 46014 2388 46020 2440
rect 46072 2428 46078 2440
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 46072 2400 46489 2428
rect 46072 2388 46078 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 46477 2391 46535 2397
rect 23256 2332 23888 2360
rect 23256 2320 23262 2332
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26237 2363 26295 2369
rect 26237 2329 26249 2363
rect 26283 2360 26295 2363
rect 26418 2360 26424 2372
rect 26283 2332 26424 2360
rect 26283 2329 26295 2332
rect 26237 2323 26295 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27120 2332 27445 2360
rect 27120 2320 27126 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 35434 2320 35440 2372
rect 35492 2360 35498 2372
rect 35621 2363 35679 2369
rect 35621 2360 35633 2363
rect 35492 2332 35633 2360
rect 35492 2320 35498 2332
rect 35621 2329 35633 2332
rect 35667 2329 35679 2363
rect 35621 2323 35679 2329
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39356 2332 40325 2360
rect 39356 2320 39362 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 45373 2363 45431 2369
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 47765 2363 47823 2369
rect 47765 2329 47777 2363
rect 47811 2360 47823 2363
rect 48314 2360 48320 2372
rect 47811 2332 48320 2360
rect 47811 2329 47823 2332
rect 47765 2323 47823 2329
rect 48314 2320 48320 2332
rect 48372 2320 48378 2372
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 5261 2295 5319 2301
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 15378 2292 15384 2304
rect 5307 2264 15384 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 19150 2252 19156 2304
rect 19208 2292 19214 2304
rect 21818 2292 21824 2304
rect 19208 2264 21824 2292
rect 19208 2252 19214 2264
rect 21818 2252 21824 2264
rect 21876 2252 21882 2304
rect 21910 2252 21916 2304
rect 21968 2252 21974 2304
rect 25038 2252 25044 2304
rect 25096 2292 25102 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 25096 2264 28641 2292
rect 25096 2252 25102 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 45462 2292 45468 2304
rect 45423 2264 45468 2292
rect 28629 2255 28687 2261
rect 45462 2252 45468 2264
rect 45520 2252 45526 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 17310 2048 17316 2100
rect 17368 2088 17374 2100
rect 25498 2088 25504 2100
rect 17368 2060 25504 2088
rect 17368 2048 17374 2060
rect 25498 2048 25504 2060
rect 25556 2048 25562 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 28074 2020 28080 2032
rect 3108 1992 28080 2020
rect 3108 1980 3114 1992
rect 28074 1980 28080 1992
rect 28132 1980 28138 2032
rect 20990 1912 20996 1964
rect 21048 1952 21054 1964
rect 45462 1952 45468 1964
rect 21048 1924 45468 1952
rect 21048 1912 21054 1924
rect 45462 1912 45468 1924
rect 45520 1912 45526 1964
rect 21818 1844 21824 1896
rect 21876 1884 21882 1896
rect 35986 1884 35992 1896
rect 21876 1856 35992 1884
rect 21876 1844 21882 1856
rect 35986 1844 35992 1856
rect 36044 1844 36050 1896
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19984 47200 20036 47252
rect 20260 47132 20312 47184
rect 29368 47132 29420 47184
rect 3056 47064 3108 47116
rect 20076 47107 20128 47116
rect 1952 46996 2004 47048
rect 2780 46996 2832 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7104 46996 7156 47048
rect 9036 46996 9088 47048
rect 11612 46996 11664 47048
rect 11980 47039 12032 47048
rect 11980 47005 11989 47039
rect 11989 47005 12023 47039
rect 12023 47005 12032 47039
rect 11980 46996 12032 47005
rect 12900 46996 12952 47048
rect 13820 46996 13872 47048
rect 16488 46996 16540 47048
rect 16948 47039 17000 47048
rect 16948 47005 16957 47039
rect 16957 47005 16991 47039
rect 16991 47005 17000 47039
rect 16948 46996 17000 47005
rect 18696 46996 18748 47048
rect 2320 46971 2372 46980
rect 2320 46937 2329 46971
rect 2329 46937 2363 46971
rect 2363 46937 2372 46971
rect 2320 46928 2372 46937
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 7840 46928 7892 46980
rect 3148 46903 3200 46912
rect 3148 46869 3157 46903
rect 3157 46869 3191 46903
rect 3191 46869 3200 46903
rect 3148 46860 3200 46869
rect 6920 46903 6972 46912
rect 6920 46869 6929 46903
rect 6929 46869 6963 46903
rect 6963 46869 6972 46903
rect 9312 46903 9364 46912
rect 6920 46860 6972 46869
rect 9312 46869 9321 46903
rect 9321 46869 9355 46903
rect 9355 46869 9364 46903
rect 9312 46860 9364 46869
rect 12256 46860 12308 46912
rect 14648 46928 14700 46980
rect 15384 46928 15436 46980
rect 20076 47073 20085 47107
rect 20085 47073 20119 47107
rect 20119 47073 20128 47107
rect 20076 47064 20128 47073
rect 26608 47064 26660 47116
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 20352 47039 20404 47048
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 24584 46996 24636 47048
rect 25412 47039 25464 47048
rect 25412 47005 25421 47039
rect 25421 47005 25455 47039
rect 25455 47005 25464 47039
rect 25412 46996 25464 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 31024 47039 31076 47048
rect 31024 47005 31033 47039
rect 31033 47005 31067 47039
rect 31067 47005 31076 47039
rect 31024 46996 31076 47005
rect 22192 46928 22244 46980
rect 26700 46928 26752 46980
rect 46756 47064 46808 47116
rect 48320 47064 48372 47116
rect 38108 46996 38160 47048
rect 41880 47039 41932 47048
rect 41880 47005 41889 47039
rect 41889 47005 41923 47039
rect 41923 47005 41932 47039
rect 41880 46996 41932 47005
rect 42616 47039 42668 47048
rect 42616 47005 42625 47039
rect 42625 47005 42659 47039
rect 42659 47005 42668 47039
rect 42616 46996 42668 47005
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 28264 46860 28316 46912
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 42800 46971 42852 46980
rect 42800 46937 42809 46971
rect 42809 46937 42843 46971
rect 42843 46937 42852 46971
rect 42800 46928 42852 46937
rect 45376 46971 45428 46980
rect 43168 46860 43220 46912
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 3148 46588 3200 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 24584 46563 24636 46572
rect 24584 46529 24593 46563
rect 24593 46529 24627 46563
rect 24627 46529 24636 46563
rect 24584 46520 24636 46529
rect 28264 46563 28316 46572
rect 28264 46529 28273 46563
rect 28273 46529 28307 46563
rect 28307 46529 28316 46563
rect 28264 46520 28316 46529
rect 3884 46452 3936 46504
rect 3976 46452 4028 46504
rect 11704 46495 11756 46504
rect 11704 46461 11713 46495
rect 11713 46461 11747 46495
rect 11747 46461 11756 46495
rect 11704 46452 11756 46461
rect 13820 46495 13872 46504
rect 13820 46461 13829 46495
rect 13829 46461 13863 46495
rect 13863 46461 13872 46495
rect 13820 46452 13872 46461
rect 14004 46495 14056 46504
rect 14004 46461 14013 46495
rect 14013 46461 14047 46495
rect 14047 46461 14056 46495
rect 14004 46452 14056 46461
rect 14188 46452 14240 46504
rect 19432 46495 19484 46504
rect 19432 46461 19441 46495
rect 19441 46461 19475 46495
rect 19475 46461 19484 46495
rect 19432 46452 19484 46461
rect 20168 46452 20220 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 32220 46384 32272 46436
rect 38384 46588 38436 46640
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 46756 46588 46808 46640
rect 41880 46520 41932 46572
rect 47860 46563 47912 46572
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 38292 46495 38344 46504
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 1676 46316 1728 46368
rect 1952 46316 2004 46368
rect 10968 46316 11020 46368
rect 20720 46316 20772 46368
rect 41328 46316 41380 46368
rect 42524 46384 42576 46436
rect 46296 46452 46348 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 47768 46384 47820 46436
rect 43536 46316 43588 46368
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3884 46155 3936 46164
rect 3884 46121 3893 46155
rect 3893 46121 3927 46155
rect 3927 46121 3936 46155
rect 3884 46112 3936 46121
rect 11704 46112 11756 46164
rect 13820 46112 13872 46164
rect 20168 46155 20220 46164
rect 20168 46121 20177 46155
rect 20177 46121 20211 46155
rect 20211 46121 20220 46155
rect 20168 46112 20220 46121
rect 24768 46112 24820 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 20720 46019 20772 46028
rect 20720 45985 20729 46019
rect 20729 45985 20763 46019
rect 20763 45985 20772 46019
rect 20720 45976 20772 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25412 45976 25464 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41972 46019 42024 46028
rect 41972 45985 41981 46019
rect 41981 45985 42015 46019
rect 42015 45985 42024 46019
rect 41972 45976 42024 45985
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 2872 45815 2924 45824
rect 2872 45781 2881 45815
rect 2881 45781 2915 45815
rect 2915 45781 2924 45815
rect 2872 45772 2924 45781
rect 14096 45908 14148 45960
rect 20076 45951 20128 45960
rect 20076 45917 20085 45951
rect 20085 45917 20119 45951
rect 20119 45917 20128 45951
rect 20076 45908 20128 45917
rect 24676 45908 24728 45960
rect 38200 45951 38252 45960
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 38384 45908 38436 45960
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 45836 45908 45888 45960
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 41512 45883 41564 45892
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 25320 45772 25372 45824
rect 33324 45772 33376 45824
rect 45560 45772 45612 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 14004 45568 14056 45620
rect 14096 45568 14148 45620
rect 20904 45611 20956 45620
rect 2872 45500 2924 45552
rect 20904 45577 20913 45611
rect 20913 45577 20947 45611
rect 20947 45577 20956 45611
rect 20904 45568 20956 45577
rect 25412 45568 25464 45620
rect 32312 45568 32364 45620
rect 41512 45568 41564 45620
rect 45100 45568 45152 45620
rect 45652 45568 45704 45620
rect 46388 45568 46440 45620
rect 1952 45475 2004 45484
rect 1952 45441 1961 45475
rect 1961 45441 1995 45475
rect 1995 45441 2004 45475
rect 1952 45432 2004 45441
rect 13728 45475 13780 45484
rect 13728 45441 13737 45475
rect 13737 45441 13771 45475
rect 13771 45441 13780 45475
rect 13728 45432 13780 45441
rect 19432 45432 19484 45484
rect 24676 45500 24728 45552
rect 25320 45432 25372 45484
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 20076 45364 20128 45416
rect 40684 45500 40736 45552
rect 42800 45543 42852 45552
rect 42800 45509 42809 45543
rect 42809 45509 42843 45543
rect 42843 45509 42852 45543
rect 42800 45500 42852 45509
rect 45376 45500 45428 45552
rect 32220 45432 32272 45484
rect 44180 45432 44232 45484
rect 47584 45432 47636 45484
rect 44456 45364 44508 45416
rect 45100 45364 45152 45416
rect 45652 45407 45704 45416
rect 45652 45373 45661 45407
rect 45661 45373 45695 45407
rect 45695 45373 45704 45407
rect 45652 45364 45704 45373
rect 47400 45364 47452 45416
rect 43996 45271 44048 45280
rect 43996 45237 44005 45271
rect 44005 45237 44039 45271
rect 44039 45237 44048 45271
rect 43996 45228 44048 45237
rect 45468 45228 45520 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 42616 45024 42668 45076
rect 44456 45067 44508 45076
rect 44456 45033 44465 45067
rect 44465 45033 44499 45067
rect 44499 45033 44508 45067
rect 44456 45024 44508 45033
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 46480 45024 46532 45076
rect 40684 44956 40736 45008
rect 47584 44956 47636 45008
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 44916 44820 44968 44872
rect 45652 44863 45704 44872
rect 45652 44829 45661 44863
rect 45661 44829 45695 44863
rect 45695 44829 45704 44863
rect 45652 44820 45704 44829
rect 46940 44752 46992 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 46296 44523 46348 44532
rect 46296 44489 46305 44523
rect 46305 44489 46339 44523
rect 46339 44489 46348 44523
rect 46296 44480 46348 44489
rect 46940 44523 46992 44532
rect 46940 44489 46949 44523
rect 46949 44489 46983 44523
rect 46983 44489 46992 44523
rect 46940 44480 46992 44489
rect 46020 44412 46072 44464
rect 45192 44344 45244 44396
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 45652 44276 45704 44328
rect 47676 44183 47728 44192
rect 47676 44149 47685 44183
rect 47685 44149 47719 44183
rect 47719 44149 47728 44183
rect 47676 44140 47728 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 47676 43800 47728 43852
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 47768 43299 47820 43308
rect 47768 43265 47777 43299
rect 47777 43265 47811 43299
rect 47811 43265 47820 43299
rect 47768 43256 47820 43265
rect 1492 43188 1544 43240
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 46296 42168 46348 42220
rect 47400 42168 47452 42220
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46480 41216 46532 41268
rect 2412 41080 2464 41132
rect 46756 41123 46808 41132
rect 46756 41089 46765 41123
rect 46765 41089 46799 41123
rect 46799 41089 46808 41123
rect 46756 41080 46808 41089
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 43444 40876 43496 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 2044 40443 2096 40452
rect 2044 40409 2053 40443
rect 2053 40409 2087 40443
rect 2087 40409 2096 40443
rect 2044 40400 2096 40409
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 46940 39312 46992 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 46940 39083 46992 39092
rect 46940 39049 46949 39083
rect 46949 39049 46983 39083
rect 46983 39049 46992 39083
rect 46940 39040 46992 39049
rect 3516 38972 3568 39024
rect 7564 38972 7616 39024
rect 46756 38904 46808 38956
rect 47676 38947 47728 38956
rect 47676 38913 47685 38947
rect 47685 38913 47719 38947
rect 47719 38913 47728 38947
rect 47676 38904 47728 38913
rect 47860 38879 47912 38888
rect 47860 38845 47869 38879
rect 47869 38845 47903 38879
rect 47903 38845 47912 38879
rect 47860 38836 47912 38845
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 26608 38539 26660 38548
rect 26608 38505 26617 38539
rect 26617 38505 26651 38539
rect 26651 38505 26660 38539
rect 26608 38496 26660 38505
rect 22652 38335 22704 38344
rect 22652 38301 22661 38335
rect 22661 38301 22695 38335
rect 22695 38301 22704 38335
rect 22652 38292 22704 38301
rect 27528 38403 27580 38412
rect 27528 38369 27537 38403
rect 27537 38369 27571 38403
rect 27571 38369 27580 38403
rect 27528 38360 27580 38369
rect 22836 38156 22888 38208
rect 26148 38199 26200 38208
rect 26148 38165 26157 38199
rect 26157 38165 26191 38199
rect 26191 38165 26200 38199
rect 26148 38156 26200 38165
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 47676 38224 47728 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 27436 38199 27488 38208
rect 27436 38165 27445 38199
rect 27445 38165 27479 38199
rect 27479 38165 27488 38199
rect 27436 38156 27488 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 47676 37995 47728 38004
rect 47676 37961 47685 37995
rect 47685 37961 47719 37995
rect 47719 37961 47728 37995
rect 47676 37952 47728 37961
rect 22836 37927 22888 37936
rect 22836 37893 22845 37927
rect 22845 37893 22879 37927
rect 22879 37893 22888 37927
rect 22836 37884 22888 37893
rect 23848 37884 23900 37936
rect 26148 37884 26200 37936
rect 27988 37884 28040 37936
rect 32220 37816 32272 37868
rect 24216 37612 24268 37664
rect 24308 37655 24360 37664
rect 24308 37621 24317 37655
rect 24317 37621 24351 37655
rect 24351 37621 24360 37655
rect 27252 37748 27304 37800
rect 24308 37612 24360 37621
rect 28540 37612 28592 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 22652 37408 22704 37460
rect 23480 37408 23532 37460
rect 27436 37408 27488 37460
rect 46296 37408 46348 37460
rect 23388 37340 23440 37392
rect 27528 37340 27580 37392
rect 24492 37315 24544 37324
rect 24492 37281 24501 37315
rect 24501 37281 24535 37315
rect 24535 37281 24544 37315
rect 24492 37272 24544 37281
rect 25228 37272 25280 37324
rect 11980 37136 12032 37188
rect 23480 37136 23532 37188
rect 23848 37204 23900 37256
rect 24308 37204 24360 37256
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25872 37204 25924 37256
rect 27252 37204 27304 37256
rect 27804 37204 27856 37256
rect 27988 37247 28040 37256
rect 27988 37213 27997 37247
rect 27997 37213 28031 37247
rect 28031 37213 28040 37247
rect 27988 37204 28040 37213
rect 25504 37111 25556 37120
rect 25504 37077 25513 37111
rect 25513 37077 25547 37111
rect 25547 37077 25556 37111
rect 25504 37068 25556 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 22560 36864 22612 36916
rect 45560 36864 45612 36916
rect 25504 36796 25556 36848
rect 29828 36796 29880 36848
rect 28540 36771 28592 36780
rect 28540 36737 28549 36771
rect 28549 36737 28583 36771
rect 28583 36737 28592 36771
rect 28540 36728 28592 36737
rect 24216 36660 24268 36712
rect 26148 36660 26200 36712
rect 28816 36703 28868 36712
rect 28816 36669 28825 36703
rect 28825 36669 28859 36703
rect 28859 36669 28868 36703
rect 28816 36660 28868 36669
rect 25504 36524 25556 36576
rect 28264 36592 28316 36644
rect 26332 36524 26384 36576
rect 30288 36567 30340 36576
rect 30288 36533 30297 36567
rect 30297 36533 30331 36567
rect 30331 36533 30340 36567
rect 30288 36524 30340 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2044 36320 2096 36372
rect 24492 36363 24544 36372
rect 24492 36329 24501 36363
rect 24501 36329 24535 36363
rect 24535 36329 24544 36363
rect 24492 36320 24544 36329
rect 24584 36320 24636 36372
rect 26148 36363 26200 36372
rect 26148 36329 26157 36363
rect 26157 36329 26191 36363
rect 26191 36329 26200 36363
rect 26148 36320 26200 36329
rect 28724 36320 28776 36372
rect 29828 36320 29880 36372
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 22560 36184 22612 36236
rect 23204 36184 23256 36236
rect 26056 36252 26108 36304
rect 2228 36048 2280 36100
rect 20812 36023 20864 36032
rect 20812 35989 20821 36023
rect 20821 35989 20855 36023
rect 20855 35989 20864 36023
rect 20812 35980 20864 35989
rect 25044 36048 25096 36100
rect 22468 36023 22520 36032
rect 22468 35989 22477 36023
rect 22477 35989 22511 36023
rect 22511 35989 22520 36023
rect 25504 36116 25556 36168
rect 26148 36184 26200 36236
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 26332 36116 26384 36168
rect 26240 36048 26292 36100
rect 28172 36116 28224 36168
rect 29276 36116 29328 36168
rect 22468 35980 22520 35989
rect 26148 35980 26200 36032
rect 27804 36048 27856 36100
rect 26608 36023 26660 36032
rect 26608 35989 26617 36023
rect 26617 35989 26651 36023
rect 26651 35989 26660 36023
rect 26608 35980 26660 35989
rect 28080 35980 28132 36032
rect 34520 35980 34572 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 25228 35819 25280 35828
rect 25228 35785 25237 35819
rect 25237 35785 25271 35819
rect 25271 35785 25280 35819
rect 25228 35776 25280 35785
rect 26240 35819 26292 35828
rect 26240 35785 26249 35819
rect 26249 35785 26283 35819
rect 26283 35785 26292 35819
rect 26240 35776 26292 35785
rect 27712 35776 27764 35828
rect 28816 35819 28868 35828
rect 28816 35785 28825 35819
rect 28825 35785 28859 35819
rect 28859 35785 28868 35819
rect 28816 35776 28868 35785
rect 29276 35819 29328 35828
rect 29276 35785 29285 35819
rect 29285 35785 29319 35819
rect 29319 35785 29328 35819
rect 29276 35776 29328 35785
rect 20260 35708 20312 35760
rect 27160 35751 27212 35760
rect 27160 35717 27169 35751
rect 27169 35717 27203 35751
rect 27203 35717 27212 35751
rect 27160 35708 27212 35717
rect 27252 35708 27304 35760
rect 1400 35640 1452 35692
rect 19156 35572 19208 35624
rect 20812 35572 20864 35624
rect 23112 35640 23164 35692
rect 24860 35683 24912 35692
rect 24860 35649 24869 35683
rect 24869 35649 24903 35683
rect 24903 35649 24912 35683
rect 24860 35640 24912 35649
rect 25688 35683 25740 35692
rect 25688 35649 25697 35683
rect 25697 35649 25731 35683
rect 25731 35649 25740 35683
rect 25688 35640 25740 35649
rect 26608 35640 26660 35692
rect 28080 35683 28132 35692
rect 28080 35649 28089 35683
rect 28089 35649 28123 35683
rect 28123 35649 28132 35683
rect 28080 35640 28132 35649
rect 28264 35683 28316 35692
rect 28264 35649 28273 35683
rect 28273 35649 28307 35683
rect 28307 35649 28316 35683
rect 28264 35640 28316 35649
rect 28632 35683 28684 35692
rect 21364 35572 21416 35624
rect 22468 35572 22520 35624
rect 23296 35572 23348 35624
rect 25964 35572 26016 35624
rect 27344 35615 27396 35624
rect 27344 35581 27353 35615
rect 27353 35581 27387 35615
rect 27387 35581 27396 35615
rect 28632 35649 28641 35683
rect 28641 35649 28675 35683
rect 28675 35649 28684 35683
rect 28632 35640 28684 35649
rect 30288 35640 30340 35692
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 31392 35640 31444 35649
rect 27344 35572 27396 35581
rect 31208 35572 31260 35624
rect 32128 35615 32180 35624
rect 32128 35581 32137 35615
rect 32137 35581 32171 35615
rect 32171 35581 32180 35615
rect 32128 35572 32180 35581
rect 32864 35572 32916 35624
rect 19892 35436 19944 35488
rect 25044 35479 25096 35488
rect 25044 35445 25053 35479
rect 25053 35445 25087 35479
rect 25087 35445 25096 35479
rect 25044 35436 25096 35445
rect 25412 35436 25464 35488
rect 25780 35479 25832 35488
rect 25780 35445 25789 35479
rect 25789 35445 25823 35479
rect 25823 35445 25832 35479
rect 25780 35436 25832 35445
rect 25964 35436 26016 35488
rect 27252 35436 27304 35488
rect 27712 35436 27764 35488
rect 28632 35436 28684 35488
rect 31944 35436 31996 35488
rect 33140 35436 33192 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 2044 35164 2096 35216
rect 19892 35232 19944 35284
rect 20260 35232 20312 35284
rect 28356 35232 28408 35284
rect 32864 35275 32916 35284
rect 32864 35241 32873 35275
rect 32873 35241 32907 35275
rect 32907 35241 32916 35275
rect 32864 35232 32916 35241
rect 25688 35164 25740 35216
rect 27620 35164 27672 35216
rect 24860 35096 24912 35148
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 2136 35071 2188 35080
rect 2136 35037 2145 35071
rect 2145 35037 2179 35071
rect 2179 35037 2188 35071
rect 2136 35028 2188 35037
rect 19248 35028 19300 35080
rect 23296 35071 23348 35080
rect 23296 35037 23305 35071
rect 23305 35037 23339 35071
rect 23339 35037 23348 35071
rect 23296 35028 23348 35037
rect 23940 35028 23992 35080
rect 25780 35028 25832 35080
rect 26056 35071 26108 35080
rect 26056 35037 26065 35071
rect 26065 35037 26099 35071
rect 26099 35037 26108 35071
rect 26056 35028 26108 35037
rect 26332 35028 26384 35080
rect 27160 35028 27212 35080
rect 27344 35028 27396 35080
rect 28540 35096 28592 35148
rect 32128 35164 32180 35216
rect 32956 35164 33008 35216
rect 34520 35164 34572 35216
rect 31944 35139 31996 35148
rect 31944 35105 31953 35139
rect 31953 35105 31987 35139
rect 31987 35105 31996 35139
rect 31944 35096 31996 35105
rect 32772 35096 32824 35148
rect 1492 34892 1544 34944
rect 23480 34892 23532 34944
rect 24768 34892 24820 34944
rect 26792 34892 26844 34944
rect 27712 34960 27764 35012
rect 31208 35028 31260 35080
rect 29920 35003 29972 35012
rect 29920 34969 29929 35003
rect 29929 34969 29963 35003
rect 29963 34969 29972 35003
rect 29920 34960 29972 34969
rect 30932 34960 30984 35012
rect 32864 35028 32916 35080
rect 35348 35096 35400 35148
rect 33140 34960 33192 35012
rect 28172 34892 28224 34944
rect 28540 34892 28592 34944
rect 35440 35028 35492 35080
rect 35808 35028 35860 35080
rect 47308 35071 47360 35080
rect 47308 35037 47317 35071
rect 47317 35037 47351 35071
rect 47351 35037 47360 35071
rect 47308 35028 47360 35037
rect 47492 35028 47544 35080
rect 35532 34960 35584 35012
rect 34520 34892 34572 34944
rect 35716 34935 35768 34944
rect 35716 34901 35725 34935
rect 35725 34901 35759 34935
rect 35759 34901 35768 34935
rect 35716 34892 35768 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 25964 34731 26016 34740
rect 25964 34697 25973 34731
rect 25973 34697 26007 34731
rect 26007 34697 26016 34731
rect 25964 34688 26016 34697
rect 26148 34688 26200 34740
rect 23296 34663 23348 34672
rect 23296 34629 23305 34663
rect 23305 34629 23339 34663
rect 23339 34629 23348 34663
rect 23296 34620 23348 34629
rect 23664 34620 23716 34672
rect 25780 34620 25832 34672
rect 27252 34663 27304 34672
rect 27252 34629 27261 34663
rect 27261 34629 27295 34663
rect 27295 34629 27304 34663
rect 27252 34620 27304 34629
rect 19984 34552 20036 34604
rect 25872 34552 25924 34604
rect 27712 34552 27764 34604
rect 28540 34620 28592 34672
rect 29920 34688 29972 34740
rect 30932 34731 30984 34740
rect 30932 34697 30941 34731
rect 30941 34697 30975 34731
rect 30975 34697 30984 34731
rect 30932 34688 30984 34697
rect 32864 34731 32916 34740
rect 32864 34697 32873 34731
rect 32873 34697 32907 34731
rect 32907 34697 32916 34731
rect 32864 34688 32916 34697
rect 24216 34527 24268 34536
rect 24216 34493 24225 34527
rect 24225 34493 24259 34527
rect 24259 34493 24268 34527
rect 24216 34484 24268 34493
rect 26792 34484 26844 34536
rect 28448 34552 28500 34604
rect 31392 34620 31444 34672
rect 33048 34595 33100 34604
rect 28356 34484 28408 34536
rect 29828 34484 29880 34536
rect 30472 34484 30524 34536
rect 33048 34561 33057 34595
rect 33057 34561 33091 34595
rect 33091 34561 33100 34595
rect 33048 34552 33100 34561
rect 33140 34595 33192 34604
rect 33140 34561 33149 34595
rect 33149 34561 33183 34595
rect 33183 34561 33192 34595
rect 33140 34552 33192 34561
rect 33416 34595 33468 34604
rect 33416 34561 33425 34595
rect 33425 34561 33459 34595
rect 33459 34561 33468 34595
rect 36268 34688 36320 34740
rect 34520 34620 34572 34672
rect 35716 34620 35768 34672
rect 48136 34595 48188 34604
rect 33416 34552 33468 34561
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 32956 34484 33008 34536
rect 33324 34459 33376 34468
rect 19248 34348 19300 34400
rect 23020 34348 23072 34400
rect 23388 34348 23440 34400
rect 23572 34348 23624 34400
rect 23848 34348 23900 34400
rect 33324 34425 33333 34459
rect 33333 34425 33367 34459
rect 33367 34425 33376 34459
rect 33324 34416 33376 34425
rect 29920 34391 29972 34400
rect 29920 34357 29929 34391
rect 29929 34357 29963 34391
rect 29963 34357 29972 34391
rect 29920 34348 29972 34357
rect 35716 34391 35768 34400
rect 35716 34357 35725 34391
rect 35725 34357 35759 34391
rect 35759 34357 35768 34391
rect 35716 34348 35768 34357
rect 47952 34391 48004 34400
rect 47952 34357 47961 34391
rect 47961 34357 47995 34391
rect 47995 34357 48004 34391
rect 47952 34348 48004 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14648 34144 14700 34196
rect 20352 34076 20404 34128
rect 21088 34076 21140 34128
rect 19248 33940 19300 33992
rect 19432 33847 19484 33856
rect 19432 33813 19441 33847
rect 19441 33813 19475 33847
rect 19475 33813 19484 33847
rect 19432 33804 19484 33813
rect 20720 33983 20772 33992
rect 20720 33949 20730 33983
rect 20730 33949 20764 33983
rect 20764 33949 20772 33983
rect 20720 33940 20772 33949
rect 20904 33983 20956 33992
rect 20904 33949 20913 33983
rect 20913 33949 20947 33983
rect 20947 33949 20956 33983
rect 20904 33940 20956 33949
rect 21088 33983 21140 33992
rect 21088 33949 21102 33983
rect 21102 33949 21136 33983
rect 21136 33949 21140 33983
rect 21088 33940 21140 33949
rect 20904 33804 20956 33856
rect 21272 33847 21324 33856
rect 21272 33813 21281 33847
rect 21281 33813 21315 33847
rect 21315 33813 21324 33847
rect 21272 33804 21324 33813
rect 21916 33983 21968 33992
rect 21916 33949 21923 33983
rect 21923 33949 21968 33983
rect 21916 33940 21968 33949
rect 22008 33915 22060 33924
rect 22008 33881 22017 33915
rect 22017 33881 22051 33915
rect 22051 33881 22060 33915
rect 22008 33872 22060 33881
rect 22376 34187 22428 34196
rect 22376 34153 22385 34187
rect 22385 34153 22419 34187
rect 22419 34153 22428 34187
rect 22376 34144 22428 34153
rect 23296 34144 23348 34196
rect 25780 34187 25832 34196
rect 23572 34076 23624 34128
rect 25780 34153 25789 34187
rect 25789 34153 25823 34187
rect 25823 34153 25832 34187
rect 25780 34144 25832 34153
rect 27620 34076 27672 34128
rect 23388 33983 23440 33992
rect 23388 33949 23395 33983
rect 23395 33949 23440 33983
rect 23388 33940 23440 33949
rect 24032 34008 24084 34060
rect 24952 34008 25004 34060
rect 27804 34008 27856 34060
rect 29920 34076 29972 34128
rect 35348 34144 35400 34196
rect 35532 34144 35584 34196
rect 47860 34076 47912 34128
rect 34796 34051 34848 34060
rect 34796 34017 34805 34051
rect 34805 34017 34839 34051
rect 34839 34017 34848 34051
rect 34796 34008 34848 34017
rect 24492 33940 24544 33992
rect 26240 33940 26292 33992
rect 26792 33983 26844 33992
rect 26792 33949 26801 33983
rect 26801 33949 26835 33983
rect 26835 33949 26844 33983
rect 26792 33940 26844 33949
rect 28356 33940 28408 33992
rect 34520 33940 34572 33992
rect 35716 34008 35768 34060
rect 36176 34051 36228 34060
rect 35900 33983 35952 33992
rect 35900 33949 35909 33983
rect 35909 33949 35943 33983
rect 35943 33949 35952 33983
rect 35900 33940 35952 33949
rect 36176 34017 36185 34051
rect 36185 34017 36219 34051
rect 36219 34017 36228 34051
rect 36176 34008 36228 34017
rect 47952 34008 48004 34060
rect 36268 33983 36320 33992
rect 36268 33949 36277 33983
rect 36277 33949 36311 33983
rect 36311 33949 36320 33983
rect 36268 33940 36320 33949
rect 24308 33872 24360 33924
rect 24860 33872 24912 33924
rect 47492 33872 47544 33924
rect 22652 33804 22704 33856
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 46204 33804 46256 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 19156 33600 19208 33652
rect 19432 33532 19484 33584
rect 18512 33507 18564 33516
rect 18512 33473 18521 33507
rect 18521 33473 18555 33507
rect 18555 33473 18564 33507
rect 18512 33464 18564 33473
rect 21732 33532 21784 33584
rect 22284 33600 22336 33652
rect 24216 33600 24268 33652
rect 24584 33643 24636 33652
rect 24584 33609 24593 33643
rect 24593 33609 24627 33643
rect 24627 33609 24636 33643
rect 24584 33600 24636 33609
rect 28632 33643 28684 33652
rect 28632 33609 28641 33643
rect 28641 33609 28675 33643
rect 28675 33609 28684 33643
rect 28632 33600 28684 33609
rect 47860 33600 47912 33652
rect 22376 33532 22428 33584
rect 22744 33532 22796 33584
rect 26148 33532 26200 33584
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1676 33439 1728 33448
rect 1676 33405 1685 33439
rect 1685 33405 1719 33439
rect 1719 33405 1728 33439
rect 1676 33396 1728 33405
rect 21272 33396 21324 33448
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 26056 33507 26108 33516
rect 24308 33439 24360 33448
rect 24308 33405 24317 33439
rect 24317 33405 24351 33439
rect 24351 33405 24360 33439
rect 24308 33396 24360 33405
rect 20536 33260 20588 33312
rect 21180 33260 21232 33312
rect 21364 33260 21416 33312
rect 23112 33328 23164 33380
rect 26056 33473 26065 33507
rect 26065 33473 26099 33507
rect 26099 33473 26108 33507
rect 26056 33464 26108 33473
rect 28356 33532 28408 33584
rect 27620 33507 27672 33516
rect 27620 33473 27629 33507
rect 27629 33473 27663 33507
rect 27663 33473 27672 33507
rect 27620 33464 27672 33473
rect 34520 33464 34572 33516
rect 47860 33507 47912 33516
rect 47860 33473 47869 33507
rect 47869 33473 47903 33507
rect 47903 33473 47912 33507
rect 47860 33464 47912 33473
rect 27712 33396 27764 33448
rect 34612 33396 34664 33448
rect 26332 33328 26384 33380
rect 34796 33371 34848 33380
rect 34796 33337 34805 33371
rect 34805 33337 34839 33371
rect 34839 33337 34848 33371
rect 34796 33328 34848 33337
rect 35348 33328 35400 33380
rect 22468 33260 22520 33312
rect 23296 33260 23348 33312
rect 23572 33303 23624 33312
rect 23572 33269 23581 33303
rect 23581 33269 23615 33303
rect 23615 33269 23624 33303
rect 23572 33260 23624 33269
rect 25044 33260 25096 33312
rect 27988 33260 28040 33312
rect 28356 33303 28408 33312
rect 28356 33269 28365 33303
rect 28365 33269 28399 33303
rect 28399 33269 28408 33303
rect 28356 33260 28408 33269
rect 28816 33260 28868 33312
rect 29828 33260 29880 33312
rect 31760 33260 31812 33312
rect 32772 33260 32824 33312
rect 35532 33260 35584 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 20904 33056 20956 33108
rect 22652 33099 22704 33108
rect 22652 33065 22661 33099
rect 22661 33065 22695 33099
rect 22695 33065 22704 33099
rect 22652 33056 22704 33065
rect 25596 33056 25648 33108
rect 26056 33056 26108 33108
rect 28448 33099 28500 33108
rect 1492 32988 1544 33040
rect 17960 32920 18012 32972
rect 18512 32920 18564 32972
rect 19156 32852 19208 32904
rect 20536 32895 20588 32904
rect 1400 32784 1452 32836
rect 3792 32784 3844 32836
rect 17224 32827 17276 32836
rect 17224 32793 17233 32827
rect 17233 32793 17267 32827
rect 17267 32793 17276 32827
rect 17224 32784 17276 32793
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 21364 32988 21416 33040
rect 21548 32988 21600 33040
rect 22836 32988 22888 33040
rect 25228 32988 25280 33040
rect 25872 32988 25924 33040
rect 28448 33065 28457 33099
rect 28457 33065 28491 33099
rect 28491 33065 28500 33099
rect 28448 33056 28500 33065
rect 27252 32988 27304 33040
rect 30564 33056 30616 33108
rect 31576 33056 31628 33108
rect 33048 33056 33100 33108
rect 35900 33056 35952 33108
rect 23664 32920 23716 32972
rect 24400 32920 24452 32972
rect 25136 32963 25188 32972
rect 25136 32929 25145 32963
rect 25145 32929 25179 32963
rect 25179 32929 25188 32963
rect 25136 32920 25188 32929
rect 26148 32920 26200 32972
rect 29828 33031 29880 33040
rect 29828 32997 29837 33031
rect 29837 32997 29871 33031
rect 29871 32997 29880 33031
rect 29828 32988 29880 32997
rect 30012 32988 30064 33040
rect 20996 32784 21048 32836
rect 18052 32716 18104 32768
rect 20352 32716 20404 32768
rect 20720 32716 20772 32768
rect 21548 32784 21600 32836
rect 22652 32852 22704 32904
rect 23020 32852 23072 32904
rect 23572 32852 23624 32904
rect 25044 32852 25096 32904
rect 24308 32784 24360 32836
rect 25504 32784 25556 32836
rect 26056 32852 26108 32904
rect 28080 32920 28132 32972
rect 30656 32920 30708 32972
rect 27988 32895 28040 32904
rect 27988 32861 27997 32895
rect 27997 32861 28031 32895
rect 28031 32861 28040 32895
rect 27988 32852 28040 32861
rect 28172 32852 28224 32904
rect 28816 32852 28868 32904
rect 29000 32895 29052 32904
rect 29000 32861 29009 32895
rect 29009 32861 29043 32895
rect 29043 32861 29052 32895
rect 29000 32852 29052 32861
rect 30012 32852 30064 32904
rect 30472 32895 30524 32904
rect 30472 32861 30481 32895
rect 30481 32861 30515 32895
rect 30515 32861 30524 32895
rect 30472 32852 30524 32861
rect 30564 32895 30616 32904
rect 30564 32861 30573 32895
rect 30573 32861 30607 32895
rect 30607 32861 30616 32895
rect 33416 32988 33468 33040
rect 31760 32963 31812 32972
rect 31760 32929 31769 32963
rect 31769 32929 31803 32963
rect 31803 32929 31812 32963
rect 31760 32920 31812 32929
rect 35716 32920 35768 32972
rect 30564 32852 30616 32861
rect 31668 32895 31720 32904
rect 29552 32784 29604 32836
rect 31668 32861 31677 32895
rect 31677 32861 31711 32895
rect 31711 32861 31720 32895
rect 31668 32852 31720 32861
rect 32220 32895 32272 32904
rect 32220 32861 32229 32895
rect 32229 32861 32263 32895
rect 32263 32861 32272 32895
rect 32220 32852 32272 32861
rect 34796 32852 34848 32904
rect 35440 32852 35492 32904
rect 35808 32895 35860 32904
rect 35808 32861 35817 32895
rect 35817 32861 35851 32895
rect 35851 32861 35860 32895
rect 35808 32852 35860 32861
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 23020 32716 23072 32768
rect 25872 32716 25924 32768
rect 26148 32716 26200 32768
rect 28540 32716 28592 32768
rect 30380 32716 30432 32768
rect 31392 32716 31444 32768
rect 35624 32784 35676 32836
rect 47676 32784 47728 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 32588 32716 32640 32768
rect 35072 32716 35124 32768
rect 36084 32716 36136 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 17224 32512 17276 32564
rect 20536 32512 20588 32564
rect 21548 32512 21600 32564
rect 22284 32555 22336 32564
rect 22284 32521 22293 32555
rect 22293 32521 22327 32555
rect 22327 32521 22336 32555
rect 22284 32512 22336 32521
rect 22376 32512 22428 32564
rect 24124 32512 24176 32564
rect 24768 32512 24820 32564
rect 26240 32555 26292 32564
rect 1676 32444 1728 32496
rect 16948 32444 17000 32496
rect 18144 32444 18196 32496
rect 23756 32444 23808 32496
rect 24584 32487 24636 32496
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 1952 32351 2004 32360
rect 1952 32317 1961 32351
rect 1961 32317 1995 32351
rect 1995 32317 2004 32351
rect 1952 32308 2004 32317
rect 3792 32351 3844 32360
rect 3792 32317 3801 32351
rect 3801 32317 3835 32351
rect 3835 32317 3844 32351
rect 3792 32308 3844 32317
rect 18328 32419 18380 32428
rect 18328 32385 18337 32419
rect 18337 32385 18371 32419
rect 18371 32385 18380 32419
rect 18328 32376 18380 32385
rect 22652 32376 22704 32428
rect 18052 32351 18104 32360
rect 18052 32317 18061 32351
rect 18061 32317 18095 32351
rect 18095 32317 18104 32351
rect 18052 32308 18104 32317
rect 18144 32351 18196 32360
rect 18144 32317 18153 32351
rect 18153 32317 18187 32351
rect 18187 32317 18196 32351
rect 23572 32376 23624 32428
rect 23848 32419 23900 32428
rect 23848 32385 23857 32419
rect 23857 32385 23891 32419
rect 23891 32385 23900 32419
rect 23848 32376 23900 32385
rect 24584 32453 24593 32487
rect 24593 32453 24627 32487
rect 24627 32453 24636 32487
rect 24584 32444 24636 32453
rect 26240 32521 26249 32555
rect 26249 32521 26283 32555
rect 26283 32521 26292 32555
rect 26240 32512 26292 32521
rect 28264 32512 28316 32564
rect 26056 32376 26108 32428
rect 26148 32376 26200 32428
rect 28172 32444 28224 32496
rect 28816 32444 28868 32496
rect 29000 32444 29052 32496
rect 28448 32376 28500 32428
rect 28724 32419 28776 32428
rect 28724 32385 28733 32419
rect 28733 32385 28767 32419
rect 28767 32385 28776 32419
rect 28724 32376 28776 32385
rect 31852 32512 31904 32564
rect 32680 32512 32732 32564
rect 30380 32444 30432 32496
rect 31208 32376 31260 32428
rect 32404 32419 32456 32428
rect 32404 32385 32413 32419
rect 32413 32385 32447 32419
rect 32447 32385 32456 32419
rect 32404 32376 32456 32385
rect 47676 32555 47728 32564
rect 47676 32521 47685 32555
rect 47685 32521 47719 32555
rect 47719 32521 47728 32555
rect 47676 32512 47728 32521
rect 32956 32444 33008 32496
rect 35072 32487 35124 32496
rect 35072 32453 35081 32487
rect 35081 32453 35115 32487
rect 35115 32453 35124 32487
rect 35072 32444 35124 32453
rect 36084 32444 36136 32496
rect 18144 32308 18196 32317
rect 23480 32308 23532 32360
rect 24124 32351 24176 32360
rect 24124 32317 24133 32351
rect 24133 32317 24167 32351
rect 24167 32317 24176 32351
rect 24124 32308 24176 32317
rect 25136 32308 25188 32360
rect 25504 32308 25556 32360
rect 28264 32308 28316 32360
rect 29828 32351 29880 32360
rect 29828 32317 29837 32351
rect 29837 32317 29871 32351
rect 29871 32317 29880 32351
rect 29828 32308 29880 32317
rect 19340 32240 19392 32292
rect 23296 32240 23348 32292
rect 26332 32240 26384 32292
rect 31392 32308 31444 32360
rect 31576 32351 31628 32360
rect 31576 32317 31585 32351
rect 31585 32317 31619 32351
rect 31619 32317 31628 32351
rect 31576 32308 31628 32317
rect 32220 32308 32272 32360
rect 33416 32351 33468 32360
rect 23388 32172 23440 32224
rect 24584 32172 24636 32224
rect 24860 32172 24912 32224
rect 27988 32172 28040 32224
rect 28264 32172 28316 32224
rect 32036 32240 32088 32292
rect 33416 32317 33425 32351
rect 33425 32317 33459 32351
rect 33459 32317 33468 32351
rect 33416 32308 33468 32317
rect 46848 32376 46900 32428
rect 47584 32419 47636 32428
rect 47584 32385 47593 32419
rect 47593 32385 47627 32419
rect 47627 32385 47636 32419
rect 47584 32376 47636 32385
rect 34704 32308 34756 32360
rect 34796 32240 34848 32292
rect 32496 32215 32548 32224
rect 32496 32181 32505 32215
rect 32505 32181 32539 32215
rect 32539 32181 32548 32215
rect 32496 32172 32548 32181
rect 35808 32172 35860 32224
rect 46848 32215 46900 32224
rect 46848 32181 46857 32215
rect 46857 32181 46891 32215
rect 46891 32181 46900 32215
rect 46848 32172 46900 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1400 32011 1452 32020
rect 1400 31977 1409 32011
rect 1409 31977 1443 32011
rect 1443 31977 1452 32011
rect 1400 31968 1452 31977
rect 21916 31968 21968 32020
rect 23388 32011 23440 32020
rect 23388 31977 23397 32011
rect 23397 31977 23431 32011
rect 23431 31977 23440 32011
rect 23388 31968 23440 31977
rect 24124 31968 24176 32020
rect 24768 31968 24820 32020
rect 1768 31900 1820 31952
rect 2044 31900 2096 31952
rect 17776 31900 17828 31952
rect 21456 31900 21508 31952
rect 22376 31900 22428 31952
rect 23020 31900 23072 31952
rect 23572 31943 23624 31952
rect 23572 31909 23581 31943
rect 23581 31909 23615 31943
rect 23615 31909 23624 31943
rect 23572 31900 23624 31909
rect 28632 31968 28684 32020
rect 30380 31968 30432 32020
rect 31668 31968 31720 32020
rect 32220 31968 32272 32020
rect 32404 31968 32456 32020
rect 34336 31968 34388 32020
rect 34796 31968 34848 32020
rect 35624 31968 35676 32020
rect 46296 31968 46348 32020
rect 9312 31832 9364 31884
rect 22284 31832 22336 31884
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 2044 31764 2096 31816
rect 2964 31807 3016 31816
rect 2964 31773 2973 31807
rect 2973 31773 3007 31807
rect 3007 31773 3016 31807
rect 2964 31764 3016 31773
rect 19984 31764 20036 31816
rect 20260 31764 20312 31816
rect 25228 31900 25280 31952
rect 25872 31900 25924 31952
rect 28908 31900 28960 31952
rect 29828 31875 29880 31884
rect 29828 31841 29837 31875
rect 29837 31841 29871 31875
rect 29871 31841 29880 31875
rect 29828 31832 29880 31841
rect 23020 31807 23072 31816
rect 22100 31696 22152 31748
rect 3056 31671 3108 31680
rect 3056 31637 3065 31671
rect 3065 31637 3099 31671
rect 3099 31637 3108 31671
rect 3056 31628 3108 31637
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 23480 31764 23532 31816
rect 25228 31807 25280 31816
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 26332 31807 26384 31816
rect 26332 31773 26341 31807
rect 26341 31773 26375 31807
rect 26375 31773 26384 31807
rect 26332 31764 26384 31773
rect 28816 31764 28868 31816
rect 30288 31764 30340 31816
rect 31576 31764 31628 31816
rect 23664 31696 23716 31748
rect 27804 31696 27856 31748
rect 27988 31696 28040 31748
rect 30380 31696 30432 31748
rect 32036 31764 32088 31816
rect 32404 31807 32456 31816
rect 32404 31773 32413 31807
rect 32413 31773 32447 31807
rect 32447 31773 32456 31807
rect 32404 31764 32456 31773
rect 33416 31900 33468 31952
rect 33600 31900 33652 31952
rect 34612 31900 34664 31952
rect 32864 31764 32916 31816
rect 32588 31696 32640 31748
rect 34704 31832 34756 31884
rect 34888 31832 34940 31884
rect 35808 31832 35860 31884
rect 33600 31807 33652 31816
rect 33600 31773 33609 31807
rect 33609 31773 33643 31807
rect 33643 31773 33652 31807
rect 33600 31764 33652 31773
rect 34336 31764 34388 31816
rect 34428 31764 34480 31816
rect 46848 31832 46900 31884
rect 36268 31807 36320 31816
rect 34520 31696 34572 31748
rect 34796 31696 34848 31748
rect 36268 31773 36277 31807
rect 36277 31773 36311 31807
rect 36311 31773 36320 31807
rect 36268 31764 36320 31773
rect 22836 31628 22888 31680
rect 27712 31628 27764 31680
rect 28448 31628 28500 31680
rect 32956 31671 33008 31680
rect 32956 31637 32965 31671
rect 32965 31637 32999 31671
rect 32999 31637 33008 31671
rect 32956 31628 33008 31637
rect 35900 31628 35952 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 3056 31356 3108 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 17960 31424 18012 31476
rect 18604 31356 18656 31408
rect 19156 31288 19208 31340
rect 20904 31424 20956 31476
rect 22560 31424 22612 31476
rect 22744 31424 22796 31476
rect 23664 31424 23716 31476
rect 23940 31424 23992 31476
rect 27804 31424 27856 31476
rect 31208 31467 31260 31476
rect 31208 31433 31217 31467
rect 31217 31433 31251 31467
rect 31251 31433 31260 31467
rect 31208 31424 31260 31433
rect 34336 31467 34388 31476
rect 34336 31433 34345 31467
rect 34345 31433 34379 31467
rect 34379 31433 34388 31467
rect 34336 31424 34388 31433
rect 34704 31424 34756 31476
rect 35716 31467 35768 31476
rect 20996 31356 21048 31408
rect 20904 31331 20956 31340
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 19248 31220 19300 31272
rect 20904 31297 20913 31331
rect 20913 31297 20947 31331
rect 20947 31297 20956 31331
rect 20904 31288 20956 31297
rect 21088 31331 21140 31340
rect 21088 31297 21097 31331
rect 21097 31297 21131 31331
rect 21131 31297 21140 31331
rect 22192 31356 22244 31408
rect 23020 31356 23072 31408
rect 28172 31356 28224 31408
rect 21088 31288 21140 31297
rect 22284 31288 22336 31340
rect 19064 31127 19116 31136
rect 19064 31093 19073 31127
rect 19073 31093 19107 31127
rect 19107 31093 19116 31127
rect 19064 31084 19116 31093
rect 19432 31084 19484 31136
rect 24952 31288 25004 31340
rect 25228 31288 25280 31340
rect 27252 31331 27304 31340
rect 27252 31297 27268 31331
rect 27268 31297 27302 31331
rect 27302 31297 27304 31331
rect 27252 31288 27304 31297
rect 27528 31331 27580 31340
rect 25504 31263 25556 31272
rect 25504 31229 25513 31263
rect 25513 31229 25547 31263
rect 25547 31229 25556 31263
rect 25504 31220 25556 31229
rect 26240 31220 26292 31272
rect 27528 31297 27537 31331
rect 27537 31297 27571 31331
rect 27571 31297 27580 31331
rect 27528 31288 27580 31297
rect 27620 31331 27672 31340
rect 27620 31297 27629 31331
rect 27629 31297 27663 31331
rect 27663 31297 27672 31331
rect 27620 31288 27672 31297
rect 28264 31288 28316 31340
rect 29276 31356 29328 31408
rect 32956 31356 33008 31408
rect 33508 31356 33560 31408
rect 29184 31331 29236 31340
rect 29184 31297 29193 31331
rect 29193 31297 29227 31331
rect 29227 31297 29236 31331
rect 29184 31288 29236 31297
rect 28448 31220 28500 31272
rect 31852 31288 31904 31340
rect 35348 31356 35400 31408
rect 35716 31433 35725 31467
rect 35725 31433 35759 31467
rect 35759 31433 35768 31467
rect 35716 31424 35768 31433
rect 34888 31331 34940 31340
rect 34888 31297 34897 31331
rect 34897 31297 34931 31331
rect 34931 31297 34940 31331
rect 34888 31288 34940 31297
rect 35532 31288 35584 31340
rect 33416 31220 33468 31272
rect 30380 31152 30432 31204
rect 30748 31152 30800 31204
rect 21824 31127 21876 31136
rect 21824 31093 21833 31127
rect 21833 31093 21867 31127
rect 21867 31093 21876 31127
rect 21824 31084 21876 31093
rect 24032 31127 24084 31136
rect 24032 31093 24041 31127
rect 24041 31093 24075 31127
rect 24075 31093 24084 31127
rect 24032 31084 24084 31093
rect 24584 31084 24636 31136
rect 26792 31084 26844 31136
rect 34796 31127 34848 31136
rect 34796 31093 34805 31127
rect 34805 31093 34839 31127
rect 34839 31093 34848 31127
rect 34796 31084 34848 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 18604 30880 18656 30932
rect 19248 30923 19300 30932
rect 19248 30889 19257 30923
rect 19257 30889 19291 30923
rect 19291 30889 19300 30923
rect 19248 30880 19300 30889
rect 20536 30880 20588 30932
rect 27896 30880 27948 30932
rect 28448 30880 28500 30932
rect 33508 30923 33560 30932
rect 33508 30889 33517 30923
rect 33517 30889 33551 30923
rect 33551 30889 33560 30923
rect 33508 30880 33560 30889
rect 19340 30812 19392 30864
rect 20628 30812 20680 30864
rect 19064 30744 19116 30796
rect 19156 30676 19208 30728
rect 20352 30676 20404 30728
rect 20904 30812 20956 30864
rect 24308 30812 24360 30864
rect 21824 30744 21876 30796
rect 22284 30787 22336 30796
rect 22284 30753 22293 30787
rect 22293 30753 22327 30787
rect 22327 30753 22336 30787
rect 22284 30744 22336 30753
rect 23388 30744 23440 30796
rect 21088 30676 21140 30728
rect 21364 30719 21416 30728
rect 21364 30685 21373 30719
rect 21373 30685 21407 30719
rect 21407 30685 21416 30719
rect 22560 30719 22612 30728
rect 21364 30676 21416 30685
rect 22560 30685 22569 30719
rect 22569 30685 22603 30719
rect 22603 30685 22612 30719
rect 22560 30676 22612 30685
rect 20628 30608 20680 30660
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 26240 30744 26292 30796
rect 26792 30676 26844 30728
rect 28724 30676 28776 30728
rect 32496 30744 32548 30796
rect 20444 30540 20496 30592
rect 21640 30583 21692 30592
rect 21640 30549 21649 30583
rect 21649 30549 21683 30583
rect 21683 30549 21692 30583
rect 21640 30540 21692 30549
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 23848 30540 23900 30592
rect 25964 30651 26016 30660
rect 25964 30617 25973 30651
rect 25973 30617 26007 30651
rect 26007 30617 26016 30651
rect 25964 30608 26016 30617
rect 29184 30608 29236 30660
rect 30472 30676 30524 30728
rect 32312 30719 32364 30728
rect 32312 30685 32321 30719
rect 32321 30685 32355 30719
rect 32355 30685 32364 30719
rect 32312 30676 32364 30685
rect 32588 30719 32640 30728
rect 31392 30608 31444 30660
rect 32588 30685 32597 30719
rect 32597 30685 32631 30719
rect 32631 30685 32640 30719
rect 32588 30676 32640 30685
rect 33416 30719 33468 30728
rect 33416 30685 33425 30719
rect 33425 30685 33459 30719
rect 33459 30685 33468 30719
rect 33416 30676 33468 30685
rect 32496 30608 32548 30660
rect 29276 30540 29328 30592
rect 32404 30540 32456 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19432 30268 19484 30320
rect 20812 30336 20864 30388
rect 46848 30336 46900 30388
rect 20536 30243 20588 30252
rect 20536 30209 20545 30243
rect 20545 30209 20579 30243
rect 20579 30209 20588 30243
rect 20536 30200 20588 30209
rect 20628 30200 20680 30252
rect 21364 30268 21416 30320
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 24032 30268 24084 30320
rect 25872 30311 25924 30320
rect 25872 30277 25881 30311
rect 25881 30277 25915 30311
rect 25915 30277 25924 30311
rect 25872 30268 25924 30277
rect 28540 30268 28592 30320
rect 22192 30200 22244 30252
rect 23020 30200 23072 30252
rect 25044 30200 25096 30252
rect 26332 30200 26384 30252
rect 17868 30175 17920 30184
rect 17868 30141 17877 30175
rect 17877 30141 17911 30175
rect 17911 30141 17920 30175
rect 17868 30132 17920 30141
rect 20996 30132 21048 30184
rect 23204 30175 23256 30184
rect 23204 30141 23213 30175
rect 23213 30141 23247 30175
rect 23247 30141 23256 30175
rect 23204 30132 23256 30141
rect 23848 30132 23900 30184
rect 24952 30175 25004 30184
rect 24952 30141 24961 30175
rect 24961 30141 24995 30175
rect 24995 30141 25004 30175
rect 24952 30132 25004 30141
rect 28356 30200 28408 30252
rect 28724 30200 28776 30252
rect 29552 30268 29604 30320
rect 30288 30268 30340 30320
rect 29920 30200 29972 30252
rect 33416 30200 33468 30252
rect 30104 30132 30156 30184
rect 25504 30064 25556 30116
rect 20628 29996 20680 30048
rect 22652 30039 22704 30048
rect 22652 30005 22661 30039
rect 22661 30005 22695 30039
rect 22695 30005 22704 30039
rect 22652 29996 22704 30005
rect 22836 29996 22888 30048
rect 28540 29996 28592 30048
rect 28908 29996 28960 30048
rect 32772 30064 32824 30116
rect 33692 29996 33744 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 20720 29835 20772 29844
rect 20720 29801 20729 29835
rect 20729 29801 20763 29835
rect 20763 29801 20772 29835
rect 20720 29792 20772 29801
rect 26240 29792 26292 29844
rect 28356 29835 28408 29844
rect 28356 29801 28365 29835
rect 28365 29801 28399 29835
rect 28399 29801 28408 29835
rect 28356 29792 28408 29801
rect 20536 29724 20588 29776
rect 23848 29724 23900 29776
rect 25136 29724 25188 29776
rect 32496 29792 32548 29844
rect 34428 29792 34480 29844
rect 18328 29656 18380 29708
rect 19984 29656 20036 29708
rect 23572 29656 23624 29708
rect 24768 29656 24820 29708
rect 20628 29631 20680 29640
rect 20628 29597 20637 29631
rect 20637 29597 20671 29631
rect 20671 29597 20680 29631
rect 20628 29588 20680 29597
rect 21088 29588 21140 29640
rect 24400 29631 24452 29640
rect 24400 29597 24409 29631
rect 24409 29597 24443 29631
rect 24443 29597 24452 29631
rect 24400 29588 24452 29597
rect 24584 29631 24636 29640
rect 24584 29597 24593 29631
rect 24593 29597 24627 29631
rect 24627 29597 24636 29631
rect 24584 29588 24636 29597
rect 25412 29588 25464 29640
rect 26332 29588 26384 29640
rect 27620 29588 27672 29640
rect 28172 29563 28224 29572
rect 15384 29452 15436 29504
rect 20536 29452 20588 29504
rect 28172 29529 28181 29563
rect 28181 29529 28215 29563
rect 28215 29529 28224 29563
rect 28172 29520 28224 29529
rect 29645 29631 29697 29640
rect 29645 29597 29654 29631
rect 29654 29597 29688 29631
rect 29688 29597 29697 29631
rect 29645 29588 29697 29597
rect 30012 29724 30064 29776
rect 30748 29631 30800 29640
rect 30748 29597 30757 29631
rect 30757 29597 30791 29631
rect 30791 29597 30800 29631
rect 30748 29588 30800 29597
rect 45376 29656 45428 29708
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 31024 29520 31076 29572
rect 32680 29563 32732 29572
rect 32680 29529 32689 29563
rect 32689 29529 32723 29563
rect 32723 29529 32732 29563
rect 32680 29520 32732 29529
rect 33692 29520 33744 29572
rect 30196 29495 30248 29504
rect 30196 29461 30205 29495
rect 30205 29461 30239 29495
rect 30239 29461 30248 29495
rect 30196 29452 30248 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 17960 29248 18012 29300
rect 18972 29248 19024 29300
rect 18328 29180 18380 29232
rect 20444 29248 20496 29300
rect 22652 29248 22704 29300
rect 21640 29180 21692 29232
rect 23756 29180 23808 29232
rect 25412 29248 25464 29300
rect 25688 29248 25740 29300
rect 26332 29248 26384 29300
rect 29644 29248 29696 29300
rect 43996 29248 44048 29300
rect 19892 29112 19944 29164
rect 14280 29087 14332 29096
rect 14280 29053 14289 29087
rect 14289 29053 14323 29087
rect 14323 29053 14332 29087
rect 14280 29044 14332 29053
rect 14464 29087 14516 29096
rect 14464 29053 14473 29087
rect 14473 29053 14507 29087
rect 14507 29053 14516 29087
rect 14464 29044 14516 29053
rect 17316 29087 17368 29096
rect 8300 28976 8352 29028
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 20536 29112 20588 29164
rect 22560 29112 22612 29164
rect 22928 29112 22980 29164
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 23940 29112 23992 29164
rect 24860 29112 24912 29164
rect 25504 29112 25556 29164
rect 20904 29044 20956 29096
rect 21088 29044 21140 29096
rect 24584 29044 24636 29096
rect 30012 29180 30064 29232
rect 30196 29180 30248 29232
rect 32680 29180 32732 29232
rect 27436 29155 27488 29164
rect 27436 29121 27445 29155
rect 27445 29121 27479 29155
rect 27479 29121 27488 29155
rect 27436 29112 27488 29121
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 28172 29112 28224 29164
rect 28540 29112 28592 29164
rect 29828 29155 29880 29164
rect 27620 29044 27672 29096
rect 28724 29087 28776 29096
rect 28724 29053 28733 29087
rect 28733 29053 28767 29087
rect 28767 29053 28776 29087
rect 28724 29044 28776 29053
rect 18972 28976 19024 29028
rect 23296 28976 23348 29028
rect 23480 28976 23532 29028
rect 23848 28976 23900 29028
rect 25596 29019 25648 29028
rect 25596 28985 25605 29019
rect 25605 28985 25639 29019
rect 25639 28985 25648 29019
rect 29828 29121 29837 29155
rect 29837 29121 29871 29155
rect 29871 29121 29880 29155
rect 29828 29112 29880 29121
rect 31208 29112 31260 29164
rect 32404 29155 32456 29164
rect 32404 29121 32413 29155
rect 32413 29121 32447 29155
rect 32447 29121 32456 29155
rect 32404 29112 32456 29121
rect 32588 29155 32640 29164
rect 32588 29121 32597 29155
rect 32597 29121 32631 29155
rect 32631 29121 32640 29155
rect 32588 29112 32640 29121
rect 32864 29112 32916 29164
rect 32496 29044 32548 29096
rect 32772 29087 32824 29096
rect 32772 29053 32781 29087
rect 32781 29053 32815 29087
rect 32815 29053 32824 29087
rect 32772 29044 32824 29053
rect 25596 28976 25648 28985
rect 18788 28951 18840 28960
rect 18788 28917 18797 28951
rect 18797 28917 18831 28951
rect 18831 28917 18840 28951
rect 18788 28908 18840 28917
rect 20536 28908 20588 28960
rect 22008 28908 22060 28960
rect 26608 28908 26660 28960
rect 29092 28908 29144 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1860 28704 1912 28756
rect 14464 28704 14516 28756
rect 17316 28704 17368 28756
rect 20444 28704 20496 28756
rect 21088 28704 21140 28756
rect 25504 28704 25556 28756
rect 31208 28704 31260 28756
rect 19984 28636 20036 28688
rect 3148 28432 3200 28484
rect 18788 28568 18840 28620
rect 20444 28568 20496 28620
rect 14648 28543 14700 28552
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 17684 28543 17736 28552
rect 17684 28509 17693 28543
rect 17693 28509 17727 28543
rect 17727 28509 17736 28543
rect 17684 28500 17736 28509
rect 17868 28543 17920 28552
rect 17868 28509 17877 28543
rect 17877 28509 17911 28543
rect 17911 28509 17920 28543
rect 17868 28500 17920 28509
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 19892 28500 19944 28552
rect 20628 28500 20680 28552
rect 20720 28500 20772 28552
rect 22008 28543 22060 28552
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 23480 28568 23532 28620
rect 24308 28568 24360 28620
rect 26240 28636 26292 28688
rect 26792 28679 26844 28688
rect 26792 28645 26801 28679
rect 26801 28645 26835 28679
rect 26835 28645 26844 28679
rect 26792 28636 26844 28645
rect 15568 28475 15620 28484
rect 15568 28441 15577 28475
rect 15577 28441 15611 28475
rect 15611 28441 15620 28475
rect 15568 28432 15620 28441
rect 7840 28364 7892 28416
rect 18144 28432 18196 28484
rect 19340 28432 19392 28484
rect 23572 28500 23624 28552
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 25412 28568 25464 28620
rect 25688 28543 25740 28552
rect 25688 28509 25697 28543
rect 25697 28509 25731 28543
rect 25731 28509 25740 28543
rect 25688 28500 25740 28509
rect 27436 28568 27488 28620
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 26884 28543 26936 28552
rect 26884 28509 26893 28543
rect 26893 28509 26927 28543
rect 26927 28509 26936 28543
rect 26884 28500 26936 28509
rect 27712 28500 27764 28552
rect 28724 28500 28776 28552
rect 30932 28500 30984 28552
rect 20904 28407 20956 28416
rect 20904 28373 20913 28407
rect 20913 28373 20947 28407
rect 20947 28373 20956 28407
rect 20904 28364 20956 28373
rect 21824 28407 21876 28416
rect 21824 28373 21833 28407
rect 21833 28373 21867 28407
rect 21867 28373 21876 28407
rect 21824 28364 21876 28373
rect 23480 28364 23532 28416
rect 23572 28407 23624 28416
rect 23572 28373 23581 28407
rect 23581 28373 23615 28407
rect 23615 28373 23624 28407
rect 23572 28364 23624 28373
rect 24216 28364 24268 28416
rect 27160 28432 27212 28484
rect 28172 28475 28224 28484
rect 28172 28441 28181 28475
rect 28181 28441 28215 28475
rect 28215 28441 28224 28475
rect 28172 28432 28224 28441
rect 26424 28407 26476 28416
rect 26424 28373 26433 28407
rect 26433 28373 26467 28407
rect 26467 28373 26476 28407
rect 26424 28364 26476 28373
rect 28448 28364 28500 28416
rect 32496 28364 32548 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 15568 28203 15620 28212
rect 15568 28169 15577 28203
rect 15577 28169 15611 28203
rect 15611 28169 15620 28203
rect 15568 28160 15620 28169
rect 14188 28092 14240 28144
rect 14648 28092 14700 28144
rect 18144 28092 18196 28144
rect 21824 28160 21876 28212
rect 19340 28092 19392 28144
rect 22928 28135 22980 28144
rect 18972 28067 19024 28076
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 22652 28067 22704 28076
rect 22652 28033 22661 28067
rect 22661 28033 22695 28067
rect 22695 28033 22704 28067
rect 22652 28024 22704 28033
rect 22928 28101 22937 28135
rect 22937 28101 22971 28135
rect 22971 28101 22980 28135
rect 22928 28092 22980 28101
rect 24032 28092 24084 28144
rect 28172 28160 28224 28212
rect 29092 28160 29144 28212
rect 28632 28092 28684 28144
rect 30288 28135 30340 28144
rect 23756 28024 23808 28076
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 24584 28024 24636 28076
rect 24768 28024 24820 28076
rect 26516 28024 26568 28076
rect 26976 28067 27028 28076
rect 26976 28033 26985 28067
rect 26985 28033 27019 28067
rect 27019 28033 27028 28067
rect 26976 28024 27028 28033
rect 27620 28024 27672 28076
rect 27712 28067 27764 28076
rect 27712 28033 27721 28067
rect 27721 28033 27755 28067
rect 27755 28033 27764 28067
rect 28540 28067 28592 28076
rect 27712 28024 27764 28033
rect 28540 28033 28549 28067
rect 28549 28033 28583 28067
rect 28583 28033 28592 28067
rect 28540 28024 28592 28033
rect 30288 28101 30297 28135
rect 30297 28101 30331 28135
rect 30331 28101 30340 28135
rect 30288 28092 30340 28101
rect 12256 27999 12308 28008
rect 12256 27965 12265 27999
rect 12265 27965 12299 27999
rect 12299 27965 12308 27999
rect 12256 27956 12308 27965
rect 12532 27999 12584 28008
rect 12532 27965 12541 27999
rect 12541 27965 12575 27999
rect 12575 27965 12584 27999
rect 12532 27956 12584 27965
rect 14556 27956 14608 28008
rect 16856 27999 16908 28008
rect 16856 27965 16865 27999
rect 16865 27965 16899 27999
rect 16899 27965 16908 27999
rect 16856 27956 16908 27965
rect 16580 27888 16632 27940
rect 17684 27956 17736 28008
rect 20628 27956 20680 28008
rect 22744 27931 22796 27940
rect 22744 27897 22753 27931
rect 22753 27897 22787 27931
rect 22787 27897 22796 27931
rect 22744 27888 22796 27897
rect 26884 27956 26936 28008
rect 28908 27956 28960 28008
rect 30564 28067 30616 28076
rect 30564 28033 30573 28067
rect 30573 28033 30607 28067
rect 30607 28033 30616 28067
rect 30564 28024 30616 28033
rect 30380 27956 30432 28008
rect 32496 28067 32548 28076
rect 32496 28033 32505 28067
rect 32505 28033 32539 28067
rect 32539 28033 32548 28067
rect 32496 28024 32548 28033
rect 45928 28024 45980 28076
rect 23664 27888 23716 27940
rect 20904 27820 20956 27872
rect 22836 27863 22888 27872
rect 22836 27829 22845 27863
rect 22845 27829 22879 27863
rect 22879 27829 22888 27863
rect 22836 27820 22888 27829
rect 26332 27863 26384 27872
rect 26332 27829 26341 27863
rect 26341 27829 26375 27863
rect 26375 27829 26384 27863
rect 26332 27820 26384 27829
rect 27528 27888 27580 27940
rect 29920 27888 29972 27940
rect 31392 27956 31444 28008
rect 32220 27956 32272 28008
rect 27896 27863 27948 27872
rect 27896 27829 27905 27863
rect 27905 27829 27939 27863
rect 27939 27829 27948 27863
rect 27896 27820 27948 27829
rect 28540 27820 28592 27872
rect 28908 27820 28960 27872
rect 29736 27820 29788 27872
rect 31024 27863 31076 27872
rect 31024 27829 31033 27863
rect 31033 27829 31067 27863
rect 31067 27829 31076 27863
rect 31024 27820 31076 27829
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 46480 27820 46532 27872
rect 47032 27820 47084 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 12256 27616 12308 27668
rect 12532 27659 12584 27668
rect 12532 27625 12541 27659
rect 12541 27625 12575 27659
rect 12575 27625 12584 27659
rect 12532 27616 12584 27625
rect 16856 27616 16908 27668
rect 26424 27616 26476 27668
rect 26884 27616 26936 27668
rect 29920 27659 29972 27668
rect 14188 27591 14240 27600
rect 14188 27557 14197 27591
rect 14197 27557 14231 27591
rect 14231 27557 14240 27591
rect 14188 27548 14240 27557
rect 18328 27548 18380 27600
rect 19340 27591 19392 27600
rect 19340 27557 19349 27591
rect 19349 27557 19383 27591
rect 19383 27557 19392 27591
rect 19340 27548 19392 27557
rect 21640 27548 21692 27600
rect 21916 27591 21968 27600
rect 21916 27557 21925 27591
rect 21925 27557 21959 27591
rect 21959 27557 21968 27591
rect 21916 27548 21968 27557
rect 22744 27548 22796 27600
rect 27620 27548 27672 27600
rect 16488 27523 16540 27532
rect 16488 27489 16497 27523
rect 16497 27489 16531 27523
rect 16531 27489 16540 27523
rect 16488 27480 16540 27489
rect 11428 27455 11480 27464
rect 11428 27421 11437 27455
rect 11437 27421 11471 27455
rect 11471 27421 11480 27455
rect 11428 27412 11480 27421
rect 12348 27344 12400 27396
rect 13268 27455 13320 27464
rect 13268 27421 13277 27455
rect 13277 27421 13311 27455
rect 13311 27421 13320 27455
rect 14096 27455 14148 27464
rect 13268 27412 13320 27421
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 14096 27412 14148 27421
rect 14648 27412 14700 27464
rect 16948 27412 17000 27464
rect 19432 27412 19484 27464
rect 20628 27480 20680 27532
rect 22284 27480 22336 27532
rect 29920 27625 29929 27659
rect 29929 27625 29963 27659
rect 29963 27625 29972 27659
rect 29920 27616 29972 27625
rect 31024 27616 31076 27668
rect 21088 27412 21140 27464
rect 22192 27412 22244 27464
rect 22652 27412 22704 27464
rect 23296 27412 23348 27464
rect 13360 27344 13412 27396
rect 15016 27387 15068 27396
rect 15016 27353 15025 27387
rect 15025 27353 15059 27387
rect 15059 27353 15068 27387
rect 15016 27344 15068 27353
rect 20536 27344 20588 27396
rect 22008 27344 22060 27396
rect 26332 27344 26384 27396
rect 27804 27455 27856 27464
rect 27804 27421 27813 27455
rect 27813 27421 27847 27455
rect 27847 27421 27856 27455
rect 28632 27455 28684 27464
rect 27804 27412 27856 27421
rect 28632 27421 28641 27455
rect 28641 27421 28675 27455
rect 28675 27421 28684 27455
rect 28632 27412 28684 27421
rect 27896 27344 27948 27396
rect 7564 27276 7616 27328
rect 8208 27276 8260 27328
rect 21180 27276 21232 27328
rect 26516 27276 26568 27328
rect 30932 27548 30984 27600
rect 29736 27480 29788 27532
rect 31392 27480 31444 27532
rect 47032 27548 47084 27600
rect 46480 27523 46532 27532
rect 46480 27489 46489 27523
rect 46489 27489 46523 27523
rect 46523 27489 46532 27523
rect 46480 27480 46532 27489
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 28908 27344 28960 27396
rect 29460 27344 29512 27396
rect 30196 27412 30248 27464
rect 30564 27344 30616 27396
rect 32312 27344 32364 27396
rect 29000 27276 29052 27328
rect 30380 27276 30432 27328
rect 32220 27276 32272 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 15016 27115 15068 27124
rect 15016 27081 15025 27115
rect 15025 27081 15059 27115
rect 15059 27081 15068 27115
rect 15016 27072 15068 27081
rect 12900 27004 12952 27056
rect 21180 27004 21232 27056
rect 11152 26936 11204 26988
rect 12532 26979 12584 26988
rect 12532 26945 12541 26979
rect 12541 26945 12575 26979
rect 12575 26945 12584 26979
rect 12532 26936 12584 26945
rect 13820 26936 13872 26988
rect 15016 26936 15068 26988
rect 20444 26936 20496 26988
rect 21088 26936 21140 26988
rect 22284 27072 22336 27124
rect 22468 27072 22520 27124
rect 23940 27072 23992 27124
rect 26516 27072 26568 27124
rect 29000 27072 29052 27124
rect 30012 27072 30064 27124
rect 46848 27072 46900 27124
rect 23572 27004 23624 27056
rect 21824 26936 21876 26988
rect 22284 26936 22336 26988
rect 22468 26979 22520 26988
rect 22468 26945 22477 26979
rect 22477 26945 22511 26979
rect 22511 26945 22520 26979
rect 22468 26936 22520 26945
rect 23020 26936 23072 26988
rect 26976 27004 27028 27056
rect 24768 26979 24820 26988
rect 24768 26945 24777 26979
rect 24777 26945 24811 26979
rect 24811 26945 24820 26979
rect 24768 26936 24820 26945
rect 26056 26979 26108 26988
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 31116 27004 31168 27056
rect 32312 27004 32364 27056
rect 8116 26868 8168 26920
rect 8208 26868 8260 26920
rect 22008 26868 22060 26920
rect 23112 26868 23164 26920
rect 9312 26800 9364 26852
rect 10324 26800 10376 26852
rect 28816 26800 28868 26852
rect 9680 26732 9732 26784
rect 12440 26732 12492 26784
rect 12624 26732 12676 26784
rect 15016 26732 15068 26784
rect 17960 26732 18012 26784
rect 21916 26732 21968 26784
rect 29184 26979 29236 26988
rect 29184 26945 29193 26979
rect 29193 26945 29227 26979
rect 29227 26945 29236 26979
rect 29184 26936 29236 26945
rect 31392 26936 31444 26988
rect 29828 26911 29880 26920
rect 29828 26877 29837 26911
rect 29837 26877 29871 26911
rect 29871 26877 29880 26911
rect 29828 26868 29880 26877
rect 30196 26868 30248 26920
rect 29092 26800 29144 26852
rect 29184 26800 29236 26852
rect 29460 26732 29512 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8116 26571 8168 26580
rect 8116 26537 8125 26571
rect 8125 26537 8159 26571
rect 8159 26537 8168 26571
rect 8116 26528 8168 26537
rect 12532 26571 12584 26580
rect 12532 26537 12541 26571
rect 12541 26537 12575 26571
rect 12575 26537 12584 26571
rect 12532 26528 12584 26537
rect 19432 26571 19484 26580
rect 19432 26537 19441 26571
rect 19441 26537 19475 26571
rect 19475 26537 19484 26571
rect 19432 26528 19484 26537
rect 22008 26571 22060 26580
rect 22008 26537 22017 26571
rect 22017 26537 22051 26571
rect 22051 26537 22060 26571
rect 22008 26528 22060 26537
rect 9680 26435 9732 26444
rect 9680 26401 9689 26435
rect 9689 26401 9723 26435
rect 9723 26401 9732 26435
rect 9680 26392 9732 26401
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 13268 26460 13320 26512
rect 14280 26503 14332 26512
rect 14280 26469 14289 26503
rect 14289 26469 14323 26503
rect 14323 26469 14332 26503
rect 14280 26460 14332 26469
rect 20628 26460 20680 26512
rect 23112 26528 23164 26580
rect 23204 26528 23256 26580
rect 31116 26571 31168 26580
rect 26516 26503 26568 26512
rect 11152 26392 11204 26401
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 9404 26367 9456 26376
rect 9404 26333 9413 26367
rect 9413 26333 9447 26367
rect 9447 26333 9456 26367
rect 9404 26324 9456 26333
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12164 26324 12216 26333
rect 12348 26435 12400 26444
rect 12348 26401 12357 26435
rect 12357 26401 12391 26435
rect 12391 26401 12400 26435
rect 12348 26392 12400 26401
rect 13452 26392 13504 26444
rect 21824 26392 21876 26444
rect 22284 26392 22336 26444
rect 22560 26392 22612 26444
rect 13268 26324 13320 26376
rect 13360 26367 13412 26376
rect 13360 26333 13369 26367
rect 13369 26333 13403 26367
rect 13403 26333 13412 26367
rect 13360 26324 13412 26333
rect 13820 26324 13872 26376
rect 14464 26324 14516 26376
rect 14648 26367 14700 26376
rect 14648 26333 14657 26367
rect 14657 26333 14691 26367
rect 14691 26333 14700 26367
rect 14648 26324 14700 26333
rect 20260 26324 20312 26376
rect 20536 26324 20588 26376
rect 22008 26324 22060 26376
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 23112 26392 23164 26444
rect 26516 26469 26525 26503
rect 26525 26469 26559 26503
rect 26559 26469 26568 26503
rect 26516 26460 26568 26469
rect 31116 26537 31125 26571
rect 31125 26537 31159 26571
rect 31159 26537 31168 26571
rect 31116 26528 31168 26537
rect 10416 26256 10468 26308
rect 13176 26299 13228 26308
rect 13176 26265 13185 26299
rect 13185 26265 13219 26299
rect 13219 26265 13228 26299
rect 13176 26256 13228 26265
rect 7472 26231 7524 26240
rect 7472 26197 7481 26231
rect 7481 26197 7515 26231
rect 7515 26197 7524 26231
rect 7472 26188 7524 26197
rect 14372 26256 14424 26308
rect 21548 26256 21600 26308
rect 22560 26256 22612 26308
rect 22744 26256 22796 26308
rect 23756 26324 23808 26376
rect 27712 26392 27764 26444
rect 46848 26392 46900 26444
rect 27252 26367 27304 26376
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 13452 26188 13504 26240
rect 14556 26231 14608 26240
rect 14556 26197 14565 26231
rect 14565 26197 14599 26231
rect 14599 26197 14608 26231
rect 14556 26188 14608 26197
rect 22008 26188 22060 26240
rect 23020 26188 23072 26240
rect 26792 26188 26844 26240
rect 30564 26324 30616 26376
rect 31392 26324 31444 26376
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 10416 25984 10468 26036
rect 14280 25984 14332 26036
rect 23572 25984 23624 26036
rect 7472 25916 7524 25968
rect 20260 25916 20312 25968
rect 9864 25848 9916 25900
rect 13084 25848 13136 25900
rect 15292 25848 15344 25900
rect 16120 25848 16172 25900
rect 17960 25848 18012 25900
rect 23020 25891 23072 25900
rect 23020 25857 23029 25891
rect 23029 25857 23063 25891
rect 23063 25857 23072 25891
rect 23020 25848 23072 25857
rect 23388 25891 23440 25900
rect 8300 25780 8352 25832
rect 3516 25712 3568 25764
rect 11612 25780 11664 25832
rect 12440 25780 12492 25832
rect 13912 25823 13964 25832
rect 13912 25789 13921 25823
rect 13921 25789 13955 25823
rect 13955 25789 13964 25823
rect 13912 25780 13964 25789
rect 14188 25823 14240 25832
rect 14188 25789 14197 25823
rect 14197 25789 14231 25823
rect 14231 25789 14240 25823
rect 14188 25780 14240 25789
rect 19432 25780 19484 25832
rect 13452 25687 13504 25696
rect 13452 25653 13461 25687
rect 13461 25653 13495 25687
rect 13495 25653 13504 25687
rect 13452 25644 13504 25653
rect 17132 25687 17184 25696
rect 17132 25653 17141 25687
rect 17141 25653 17175 25687
rect 17175 25653 17184 25687
rect 17132 25644 17184 25653
rect 21548 25644 21600 25696
rect 23112 25712 23164 25764
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 26516 25916 26568 25968
rect 27160 25959 27212 25968
rect 27160 25925 27169 25959
rect 27169 25925 27203 25959
rect 27203 25925 27212 25959
rect 27160 25916 27212 25925
rect 24400 25848 24452 25900
rect 26792 25848 26844 25900
rect 27344 25891 27396 25900
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 28908 25891 28960 25900
rect 27344 25848 27396 25857
rect 28908 25857 28917 25891
rect 28917 25857 28951 25891
rect 28951 25857 28960 25891
rect 28908 25848 28960 25857
rect 25780 25644 25832 25696
rect 26976 25712 27028 25764
rect 28448 25780 28500 25832
rect 29000 25780 29052 25832
rect 28632 25644 28684 25696
rect 46296 25644 46348 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 9404 25440 9456 25492
rect 11612 25483 11664 25492
rect 11612 25449 11621 25483
rect 11621 25449 11655 25483
rect 11655 25449 11664 25483
rect 11612 25440 11664 25449
rect 13084 25440 13136 25492
rect 14188 25440 14240 25492
rect 14464 25483 14516 25492
rect 14464 25449 14473 25483
rect 14473 25449 14507 25483
rect 14507 25449 14516 25483
rect 14464 25440 14516 25449
rect 15292 25440 15344 25492
rect 16120 25483 16172 25492
rect 16120 25449 16129 25483
rect 16129 25449 16163 25483
rect 16163 25449 16172 25483
rect 16120 25440 16172 25449
rect 20260 25440 20312 25492
rect 22652 25483 22704 25492
rect 22652 25449 22661 25483
rect 22661 25449 22695 25483
rect 22695 25449 22704 25483
rect 22652 25440 22704 25449
rect 27620 25483 27672 25492
rect 27620 25449 27629 25483
rect 27629 25449 27663 25483
rect 27663 25449 27672 25483
rect 27620 25440 27672 25449
rect 27804 25440 27856 25492
rect 28908 25440 28960 25492
rect 14280 25372 14332 25424
rect 19156 25372 19208 25424
rect 23204 25372 23256 25424
rect 30288 25372 30340 25424
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 8484 25236 8536 25288
rect 17132 25347 17184 25356
rect 17132 25313 17141 25347
rect 17141 25313 17175 25347
rect 17175 25313 17184 25347
rect 17132 25304 17184 25313
rect 18144 25304 18196 25356
rect 22008 25347 22060 25356
rect 10048 25279 10100 25288
rect 10048 25245 10057 25279
rect 10057 25245 10091 25279
rect 10091 25245 10100 25279
rect 10048 25236 10100 25245
rect 10324 25236 10376 25288
rect 11428 25236 11480 25288
rect 11888 25236 11940 25288
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 14004 25236 14056 25288
rect 15384 25236 15436 25288
rect 16396 25279 16448 25288
rect 14096 25168 14148 25220
rect 14832 25168 14884 25220
rect 16396 25245 16405 25279
rect 16405 25245 16439 25279
rect 16439 25245 16448 25279
rect 16396 25236 16448 25245
rect 16856 25279 16908 25288
rect 16856 25245 16865 25279
rect 16865 25245 16899 25279
rect 16899 25245 16908 25279
rect 16856 25236 16908 25245
rect 22008 25313 22017 25347
rect 22017 25313 22051 25347
rect 22051 25313 22060 25347
rect 22008 25304 22060 25313
rect 19524 25236 19576 25288
rect 19984 25236 20036 25288
rect 10140 25143 10192 25152
rect 10140 25109 10149 25143
rect 10149 25109 10183 25143
rect 10183 25109 10192 25143
rect 10140 25100 10192 25109
rect 13544 25100 13596 25152
rect 15844 25100 15896 25152
rect 16304 25143 16356 25152
rect 16304 25109 16313 25143
rect 16313 25109 16347 25143
rect 16347 25109 16356 25143
rect 16304 25100 16356 25109
rect 18420 25168 18472 25220
rect 22100 25168 22152 25220
rect 19340 25143 19392 25152
rect 19340 25109 19349 25143
rect 19349 25109 19383 25143
rect 19383 25109 19392 25143
rect 19340 25100 19392 25109
rect 21088 25100 21140 25152
rect 21364 25143 21416 25152
rect 21364 25109 21373 25143
rect 21373 25109 21407 25143
rect 21407 25109 21416 25143
rect 21364 25100 21416 25109
rect 21548 25100 21600 25152
rect 23388 25304 23440 25356
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 25780 25279 25832 25288
rect 22284 25236 22336 25245
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 26240 25236 26292 25288
rect 27252 25304 27304 25356
rect 29276 25304 29328 25356
rect 28448 25236 28500 25288
rect 28632 25279 28684 25288
rect 28632 25245 28641 25279
rect 28641 25245 28675 25279
rect 28675 25245 28684 25279
rect 28632 25236 28684 25245
rect 28724 25236 28776 25288
rect 40408 25304 40460 25356
rect 46296 25347 46348 25356
rect 46296 25313 46305 25347
rect 46305 25313 46339 25347
rect 46339 25313 46348 25347
rect 46296 25304 46348 25313
rect 29828 25279 29880 25288
rect 29828 25245 29837 25279
rect 29837 25245 29871 25279
rect 29871 25245 29880 25279
rect 30104 25279 30156 25288
rect 29828 25236 29880 25245
rect 22744 25168 22796 25220
rect 26792 25211 26844 25220
rect 26792 25177 26801 25211
rect 26801 25177 26835 25211
rect 26835 25177 26844 25211
rect 26792 25168 26844 25177
rect 27252 25168 27304 25220
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 30564 25279 30616 25288
rect 30564 25245 30573 25279
rect 30573 25245 30607 25279
rect 30607 25245 30616 25279
rect 30564 25236 30616 25245
rect 48136 25279 48188 25288
rect 48136 25245 48145 25279
rect 48145 25245 48179 25279
rect 48179 25245 48188 25279
rect 48136 25236 48188 25245
rect 47676 25168 47728 25220
rect 24952 25100 25004 25152
rect 27712 25100 27764 25152
rect 29460 25100 29512 25152
rect 30564 25100 30616 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 13912 24896 13964 24948
rect 15844 24939 15896 24948
rect 15844 24905 15853 24939
rect 15853 24905 15887 24939
rect 15887 24905 15896 24939
rect 15844 24896 15896 24905
rect 16304 24896 16356 24948
rect 16856 24939 16908 24948
rect 16856 24905 16865 24939
rect 16865 24905 16899 24939
rect 16899 24905 16908 24939
rect 16856 24896 16908 24905
rect 22100 24939 22152 24948
rect 22100 24905 22109 24939
rect 22109 24905 22143 24939
rect 22143 24905 22152 24939
rect 22100 24896 22152 24905
rect 29828 24896 29880 24948
rect 13268 24828 13320 24880
rect 46756 24828 46808 24880
rect 8484 24760 8536 24812
rect 10232 24760 10284 24812
rect 12808 24760 12860 24812
rect 13360 24760 13412 24812
rect 14372 24760 14424 24812
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 15384 24760 15436 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18420 24760 18472 24812
rect 10140 24692 10192 24744
rect 10324 24624 10376 24676
rect 12164 24624 12216 24676
rect 16396 24692 16448 24744
rect 18512 24692 18564 24744
rect 19340 24692 19392 24744
rect 22284 24692 22336 24744
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 24676 24760 24728 24812
rect 27620 24803 27672 24812
rect 27620 24769 27629 24803
rect 27629 24769 27663 24803
rect 27663 24769 27672 24803
rect 27620 24760 27672 24769
rect 30564 24760 30616 24812
rect 46572 24760 46624 24812
rect 47492 24760 47544 24812
rect 47676 24803 47728 24812
rect 47676 24769 47685 24803
rect 47685 24769 47719 24803
rect 47719 24769 47728 24803
rect 47676 24760 47728 24769
rect 20444 24624 20496 24676
rect 22928 24692 22980 24744
rect 23296 24735 23348 24744
rect 23296 24701 23305 24735
rect 23305 24701 23339 24735
rect 23339 24701 23348 24735
rect 23296 24692 23348 24701
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 26240 24692 26292 24744
rect 27712 24735 27764 24744
rect 27712 24701 27721 24735
rect 27721 24701 27755 24735
rect 27755 24701 27764 24735
rect 27712 24692 27764 24701
rect 28908 24692 28960 24744
rect 29184 24735 29236 24744
rect 29184 24701 29193 24735
rect 29193 24701 29227 24735
rect 29227 24701 29236 24735
rect 29184 24692 29236 24701
rect 29460 24735 29512 24744
rect 29460 24701 29469 24735
rect 29469 24701 29503 24735
rect 29503 24701 29512 24735
rect 29460 24692 29512 24701
rect 25964 24624 26016 24676
rect 9312 24556 9364 24608
rect 13912 24599 13964 24608
rect 13912 24565 13921 24599
rect 13921 24565 13955 24599
rect 13955 24565 13964 24599
rect 13912 24556 13964 24565
rect 14464 24556 14516 24608
rect 16672 24556 16724 24608
rect 22744 24556 22796 24608
rect 29000 24556 29052 24608
rect 46756 24692 46808 24744
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10232 24352 10284 24404
rect 15292 24352 15344 24404
rect 18512 24395 18564 24404
rect 18512 24361 18521 24395
rect 18521 24361 18555 24395
rect 18555 24361 18564 24395
rect 18512 24352 18564 24361
rect 20628 24352 20680 24404
rect 22008 24352 22060 24404
rect 22284 24352 22336 24404
rect 26792 24352 26844 24404
rect 27988 24352 28040 24404
rect 28724 24352 28776 24404
rect 28908 24395 28960 24404
rect 28908 24361 28917 24395
rect 28917 24361 28951 24395
rect 28951 24361 28960 24395
rect 29920 24395 29972 24404
rect 28908 24352 28960 24361
rect 29920 24361 29929 24395
rect 29929 24361 29963 24395
rect 29963 24361 29972 24395
rect 29920 24352 29972 24361
rect 46388 24352 46440 24404
rect 19432 24216 19484 24268
rect 23296 24216 23348 24268
rect 24952 24259 25004 24268
rect 24952 24225 24961 24259
rect 24961 24225 24995 24259
rect 24995 24225 25004 24259
rect 24952 24216 25004 24225
rect 27620 24216 27672 24268
rect 9864 24191 9916 24200
rect 9864 24157 9873 24191
rect 9873 24157 9907 24191
rect 9907 24157 9916 24191
rect 9864 24148 9916 24157
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 12900 24148 12952 24200
rect 15844 24191 15896 24200
rect 13360 24123 13412 24132
rect 13360 24089 13369 24123
rect 13369 24089 13403 24123
rect 13403 24089 13412 24123
rect 13360 24080 13412 24089
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 16396 24148 16448 24200
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 12532 24055 12584 24064
rect 12532 24021 12541 24055
rect 12541 24021 12575 24055
rect 12575 24021 12584 24055
rect 12532 24012 12584 24021
rect 16304 24012 16356 24064
rect 18328 24080 18380 24132
rect 20536 24080 20588 24132
rect 21088 24080 21140 24132
rect 25688 24080 25740 24132
rect 21364 24012 21416 24064
rect 27804 24191 27856 24200
rect 27804 24157 27813 24191
rect 27813 24157 27847 24191
rect 27847 24157 27856 24191
rect 27804 24148 27856 24157
rect 28448 24148 28500 24200
rect 28908 24216 28960 24268
rect 30288 24216 30340 24268
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 27988 24080 28040 24132
rect 30104 24148 30156 24200
rect 47768 24080 47820 24132
rect 29276 24012 29328 24064
rect 29552 24055 29604 24064
rect 29552 24021 29561 24055
rect 29561 24021 29595 24055
rect 29595 24021 29604 24055
rect 29552 24012 29604 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1768 23808 1820 23860
rect 12808 23851 12860 23860
rect 12808 23817 12817 23851
rect 12817 23817 12851 23851
rect 12851 23817 12860 23851
rect 12808 23808 12860 23817
rect 14372 23808 14424 23860
rect 16304 23808 16356 23860
rect 16764 23808 16816 23860
rect 18328 23851 18380 23860
rect 18328 23817 18337 23851
rect 18337 23817 18371 23851
rect 18371 23817 18380 23851
rect 18328 23808 18380 23817
rect 24676 23808 24728 23860
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 27896 23808 27948 23860
rect 28908 23808 28960 23860
rect 9312 23740 9364 23792
rect 12072 23740 12124 23792
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 8484 23715 8536 23724
rect 8484 23681 8493 23715
rect 8493 23681 8527 23715
rect 8527 23681 8536 23715
rect 8484 23672 8536 23681
rect 9128 23604 9180 23656
rect 9680 23715 9732 23724
rect 9680 23681 9689 23715
rect 9689 23681 9723 23715
rect 9723 23681 9732 23715
rect 9680 23672 9732 23681
rect 9864 23672 9916 23724
rect 15292 23783 15344 23792
rect 15292 23749 15301 23783
rect 15301 23749 15335 23783
rect 15335 23749 15344 23783
rect 15292 23740 15344 23749
rect 45376 23783 45428 23792
rect 45376 23749 45385 23783
rect 45385 23749 45419 23783
rect 45419 23749 45428 23783
rect 45376 23740 45428 23749
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 13544 23672 13596 23724
rect 10048 23536 10100 23588
rect 12532 23604 12584 23656
rect 15200 23672 15252 23724
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 16672 23715 16724 23724
rect 13820 23604 13872 23656
rect 15108 23604 15160 23656
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 18236 23715 18288 23724
rect 18236 23681 18245 23715
rect 18245 23681 18279 23715
rect 18279 23681 18288 23715
rect 18236 23672 18288 23681
rect 19984 23672 20036 23724
rect 24676 23672 24728 23724
rect 19432 23604 19484 23656
rect 13268 23536 13320 23588
rect 15200 23536 15252 23588
rect 15752 23536 15804 23588
rect 8392 23468 8444 23520
rect 10140 23468 10192 23520
rect 10416 23468 10468 23520
rect 15936 23468 15988 23520
rect 18972 23511 19024 23520
rect 18972 23477 18981 23511
rect 18981 23477 19015 23511
rect 19015 23477 19024 23511
rect 18972 23468 19024 23477
rect 28724 23672 28776 23724
rect 30012 23672 30064 23724
rect 47768 23715 47820 23724
rect 47768 23681 47777 23715
rect 47777 23681 47811 23715
rect 47811 23681 47820 23715
rect 47768 23672 47820 23681
rect 29552 23604 29604 23656
rect 45744 23604 45796 23656
rect 46756 23647 46808 23656
rect 46756 23613 46765 23647
rect 46765 23613 46799 23647
rect 46799 23613 46808 23647
rect 46756 23604 46808 23613
rect 29184 23468 29236 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8300 23264 8352 23316
rect 9588 23264 9640 23316
rect 10232 23307 10284 23316
rect 10232 23273 10241 23307
rect 10241 23273 10275 23307
rect 10275 23273 10284 23307
rect 10232 23264 10284 23273
rect 10416 23307 10468 23316
rect 10416 23273 10425 23307
rect 10425 23273 10459 23307
rect 10459 23273 10468 23307
rect 10416 23264 10468 23273
rect 11888 23307 11940 23316
rect 11888 23273 11897 23307
rect 11897 23273 11931 23307
rect 11931 23273 11940 23307
rect 11888 23264 11940 23273
rect 15844 23264 15896 23316
rect 19432 23307 19484 23316
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 2320 23196 2372 23248
rect 9128 23103 9180 23112
rect 9128 23069 9134 23103
rect 9134 23069 9168 23103
rect 9168 23069 9180 23103
rect 9128 23060 9180 23069
rect 8300 22924 8352 22976
rect 9680 23128 9732 23180
rect 9772 23060 9824 23112
rect 10600 23060 10652 23112
rect 10968 23035 11020 23044
rect 9588 22924 9640 22976
rect 10968 23001 10977 23035
rect 10977 23001 11011 23035
rect 11011 23001 11020 23035
rect 10968 22992 11020 23001
rect 13912 23128 13964 23180
rect 17960 23196 18012 23248
rect 22100 23264 22152 23316
rect 21088 23196 21140 23248
rect 45744 23128 45796 23180
rect 46848 23171 46900 23180
rect 46848 23137 46857 23171
rect 46857 23137 46891 23171
rect 46891 23137 46900 23171
rect 46848 23128 46900 23137
rect 13820 23060 13872 23112
rect 14464 23060 14516 23112
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 15292 23060 15344 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 20904 23060 20956 23112
rect 11244 22992 11296 23044
rect 11796 23035 11848 23044
rect 11796 23001 11805 23035
rect 11805 23001 11839 23035
rect 11839 23001 11848 23035
rect 11796 22992 11848 23001
rect 12624 22992 12676 23044
rect 13360 22992 13412 23044
rect 10232 22967 10284 22976
rect 10232 22933 10257 22967
rect 10257 22933 10284 22967
rect 10232 22924 10284 22933
rect 13636 22924 13688 22976
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14924 22967 14976 22976
rect 14924 22933 14933 22967
rect 14933 22933 14967 22967
rect 14967 22933 14976 22967
rect 14924 22924 14976 22933
rect 15476 22992 15528 23044
rect 16120 22992 16172 23044
rect 20812 22992 20864 23044
rect 22008 23035 22060 23044
rect 22008 23001 22017 23035
rect 22017 23001 22051 23035
rect 22051 23001 22060 23035
rect 22008 22992 22060 23001
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 27160 23103 27212 23112
rect 27160 23069 27169 23103
rect 27169 23069 27203 23103
rect 27203 23069 27212 23103
rect 27160 23060 27212 23069
rect 30380 22992 30432 23044
rect 45468 23060 45520 23112
rect 45836 23060 45888 23112
rect 46112 22992 46164 23044
rect 47676 22992 47728 23044
rect 19248 22924 19300 22976
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 22928 22924 22980 22976
rect 42800 22924 42852 22976
rect 45192 22924 45244 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9588 22720 9640 22772
rect 10968 22720 11020 22772
rect 8300 22695 8352 22704
rect 8300 22661 8309 22695
rect 8309 22661 8343 22695
rect 8343 22661 8352 22695
rect 8300 22652 8352 22661
rect 10140 22652 10192 22704
rect 10324 22652 10376 22704
rect 12900 22720 12952 22772
rect 13544 22720 13596 22772
rect 15108 22763 15160 22772
rect 15108 22729 15117 22763
rect 15117 22729 15151 22763
rect 15151 22729 15160 22763
rect 15108 22720 15160 22729
rect 22008 22720 22060 22772
rect 13636 22695 13688 22704
rect 13636 22661 13645 22695
rect 13645 22661 13679 22695
rect 13679 22661 13688 22695
rect 13636 22652 13688 22661
rect 14924 22652 14976 22704
rect 22928 22652 22980 22704
rect 12440 22584 12492 22636
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 16672 22584 16724 22636
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 19432 22584 19484 22636
rect 20904 22584 20956 22636
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 21088 22584 21140 22593
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 27068 22720 27120 22772
rect 47676 22763 47728 22772
rect 8392 22516 8444 22568
rect 14280 22516 14332 22568
rect 22836 22516 22888 22568
rect 24952 22516 25004 22568
rect 27160 22516 27212 22568
rect 10600 22491 10652 22500
rect 10600 22457 10609 22491
rect 10609 22457 10643 22491
rect 10643 22457 10652 22491
rect 10600 22448 10652 22457
rect 29276 22516 29328 22568
rect 47676 22729 47685 22763
rect 47685 22729 47719 22763
rect 47719 22729 47728 22763
rect 47676 22720 47728 22729
rect 44640 22627 44692 22636
rect 44640 22593 44649 22627
rect 44649 22593 44683 22627
rect 44683 22593 44692 22627
rect 44640 22584 44692 22593
rect 44916 22627 44968 22636
rect 44916 22593 44925 22627
rect 44925 22593 44959 22627
rect 44959 22593 44968 22627
rect 44916 22584 44968 22593
rect 40040 22516 40092 22568
rect 45376 22516 45428 22568
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 46204 22559 46256 22568
rect 46204 22525 46213 22559
rect 46213 22525 46247 22559
rect 46247 22525 46256 22559
rect 46204 22516 46256 22525
rect 10048 22380 10100 22432
rect 10232 22380 10284 22432
rect 12072 22380 12124 22432
rect 14832 22380 14884 22432
rect 15200 22380 15252 22432
rect 18696 22423 18748 22432
rect 18696 22389 18705 22423
rect 18705 22389 18739 22423
rect 18739 22389 18748 22423
rect 18696 22380 18748 22389
rect 19984 22380 20036 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14464 22176 14516 22228
rect 22192 22219 22244 22228
rect 22192 22185 22201 22219
rect 22201 22185 22235 22219
rect 22235 22185 22244 22219
rect 22192 22176 22244 22185
rect 22836 22219 22888 22228
rect 22836 22185 22845 22219
rect 22845 22185 22879 22219
rect 22879 22185 22888 22219
rect 22836 22176 22888 22185
rect 8116 22040 8168 22092
rect 11244 22040 11296 22092
rect 11888 22040 11940 22092
rect 15200 22083 15252 22092
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 15200 22049 15209 22083
rect 15209 22049 15243 22083
rect 15243 22049 15252 22083
rect 15200 22040 15252 22049
rect 15568 22040 15620 22092
rect 16488 22040 16540 22092
rect 17960 22083 18012 22092
rect 17960 22049 17969 22083
rect 17969 22049 18003 22083
rect 18003 22049 18012 22083
rect 17960 22040 18012 22049
rect 10876 21947 10928 21956
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 10876 21913 10885 21947
rect 10885 21913 10919 21947
rect 10919 21913 10928 21947
rect 10876 21904 10928 21913
rect 11336 21904 11388 21956
rect 10324 21836 10376 21888
rect 12624 21836 12676 21888
rect 15476 21947 15528 21956
rect 15476 21913 15485 21947
rect 15485 21913 15519 21947
rect 15519 21913 15528 21947
rect 15476 21904 15528 21913
rect 16764 21904 16816 21956
rect 17960 21836 18012 21888
rect 18696 21972 18748 22024
rect 19984 21904 20036 21956
rect 18236 21836 18288 21888
rect 22560 22040 22612 22092
rect 24952 22083 25004 22092
rect 24952 22049 24961 22083
rect 24961 22049 24995 22083
rect 24995 22049 25004 22083
rect 24952 22040 25004 22049
rect 27988 22040 28040 22092
rect 21272 21972 21324 22024
rect 22652 21972 22704 22024
rect 22008 21947 22060 21956
rect 22008 21913 22017 21947
rect 22017 21913 22051 21947
rect 22051 21913 22060 21947
rect 22008 21904 22060 21913
rect 25136 21972 25188 22024
rect 25504 22015 25556 22024
rect 25504 21981 25513 22015
rect 25513 21981 25547 22015
rect 25547 21981 25556 22015
rect 25504 21972 25556 21981
rect 29368 22040 29420 22092
rect 21916 21836 21968 21888
rect 26240 21904 26292 21956
rect 27528 21904 27580 21956
rect 29552 22015 29604 22024
rect 29552 21981 29561 22015
rect 29561 21981 29595 22015
rect 29595 21981 29604 22015
rect 29552 21972 29604 21981
rect 44916 22108 44968 22160
rect 46572 22040 46624 22092
rect 46664 22040 46716 22092
rect 37280 21972 37332 22024
rect 43444 22015 43496 22024
rect 43444 21981 43453 22015
rect 43453 21981 43487 22015
rect 43487 21981 43496 22015
rect 43444 21972 43496 21981
rect 43628 22015 43680 22024
rect 43628 21981 43637 22015
rect 43637 21981 43671 22015
rect 43671 21981 43680 22015
rect 43628 21972 43680 21981
rect 45284 22015 45336 22024
rect 45284 21981 45293 22015
rect 45293 21981 45327 22015
rect 45327 21981 45336 22015
rect 45284 21972 45336 21981
rect 22192 21879 22244 21888
rect 22192 21845 22217 21879
rect 22217 21845 22244 21879
rect 22192 21836 22244 21845
rect 22652 21836 22704 21888
rect 27988 21879 28040 21888
rect 27988 21845 27997 21879
rect 27997 21845 28031 21879
rect 28031 21845 28040 21879
rect 27988 21836 28040 21845
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 28908 21836 28960 21888
rect 39580 21904 39632 21956
rect 44456 21904 44508 21956
rect 45192 21904 45244 21956
rect 45652 21947 45704 21956
rect 45652 21913 45661 21947
rect 45661 21913 45695 21947
rect 45695 21913 45704 21947
rect 45652 21904 45704 21913
rect 47676 21904 47728 21956
rect 38568 21836 38620 21888
rect 45928 21836 45980 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11336 21632 11388 21684
rect 14832 21632 14884 21684
rect 16764 21675 16816 21684
rect 9772 21607 9824 21616
rect 9772 21573 9781 21607
rect 9781 21573 9815 21607
rect 9815 21573 9824 21607
rect 9772 21564 9824 21573
rect 15384 21564 15436 21616
rect 16764 21641 16773 21675
rect 16773 21641 16807 21675
rect 16807 21641 16816 21675
rect 16764 21632 16816 21641
rect 9864 21496 9916 21548
rect 9680 21360 9732 21412
rect 12440 21496 12492 21548
rect 1584 21292 1636 21344
rect 9956 21292 10008 21344
rect 10692 21292 10744 21344
rect 14280 21292 14332 21344
rect 15476 21428 15528 21480
rect 17960 21496 18012 21548
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 21916 21632 21968 21684
rect 22008 21632 22060 21684
rect 22560 21675 22612 21684
rect 22560 21641 22569 21675
rect 22569 21641 22603 21675
rect 22603 21641 22612 21675
rect 26240 21675 26292 21684
rect 22560 21632 22612 21641
rect 26240 21641 26249 21675
rect 26249 21641 26283 21675
rect 26283 21641 26292 21675
rect 26240 21632 26292 21641
rect 27436 21632 27488 21684
rect 28908 21632 28960 21684
rect 29276 21632 29328 21684
rect 44456 21632 44508 21684
rect 44640 21675 44692 21684
rect 44640 21641 44649 21675
rect 44649 21641 44683 21675
rect 44683 21641 44692 21675
rect 44640 21632 44692 21641
rect 27344 21564 27396 21616
rect 20260 21539 20312 21548
rect 15936 21360 15988 21412
rect 18144 21428 18196 21480
rect 18512 21403 18564 21412
rect 18512 21369 18521 21403
rect 18521 21369 18555 21403
rect 18555 21369 18564 21403
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 20904 21496 20956 21548
rect 19616 21428 19668 21480
rect 20168 21428 20220 21480
rect 21272 21428 21324 21480
rect 22100 21428 22152 21480
rect 25136 21496 25188 21548
rect 27528 21539 27580 21548
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 31392 21496 31444 21548
rect 24584 21428 24636 21480
rect 28448 21428 28500 21480
rect 22192 21403 22244 21412
rect 18512 21360 18564 21369
rect 22192 21369 22201 21403
rect 22201 21369 22235 21403
rect 22235 21369 22244 21403
rect 22192 21360 22244 21369
rect 38568 21360 38620 21412
rect 42800 21564 42852 21616
rect 39304 21471 39356 21480
rect 39304 21437 39313 21471
rect 39313 21437 39347 21471
rect 39347 21437 39356 21471
rect 39304 21428 39356 21437
rect 39580 21471 39632 21480
rect 39580 21437 39589 21471
rect 39589 21437 39623 21471
rect 39623 21437 39632 21471
rect 39580 21428 39632 21437
rect 45284 21564 45336 21616
rect 47952 21607 48004 21616
rect 47952 21573 47961 21607
rect 47961 21573 47995 21607
rect 47995 21573 48004 21607
rect 47952 21564 48004 21573
rect 44456 21539 44508 21548
rect 44456 21505 44465 21539
rect 44465 21505 44499 21539
rect 44499 21505 44508 21539
rect 44456 21496 44508 21505
rect 45652 21539 45704 21548
rect 45652 21505 45661 21539
rect 45661 21505 45695 21539
rect 45695 21505 45704 21539
rect 45652 21496 45704 21505
rect 17040 21292 17092 21344
rect 20168 21292 20220 21344
rect 20444 21292 20496 21344
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 22836 21292 22888 21344
rect 25780 21292 25832 21344
rect 46572 21292 46624 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9956 21088 10008 21140
rect 10600 21020 10652 21072
rect 22560 21020 22612 21072
rect 8116 20995 8168 21004
rect 8116 20961 8125 20995
rect 8125 20961 8159 20995
rect 8159 20961 8168 20995
rect 8116 20952 8168 20961
rect 13820 20952 13872 21004
rect 14280 20995 14332 21004
rect 14280 20961 14289 20995
rect 14289 20961 14323 20995
rect 14323 20961 14332 20995
rect 14280 20952 14332 20961
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 16488 20952 16540 21004
rect 17040 20995 17092 21004
rect 17040 20961 17049 20995
rect 17049 20961 17083 20995
rect 17083 20961 17092 20995
rect 17040 20952 17092 20961
rect 20168 20995 20220 21004
rect 20168 20961 20177 20995
rect 20177 20961 20211 20995
rect 20211 20961 20220 20995
rect 20168 20952 20220 20961
rect 20444 20995 20496 21004
rect 20444 20961 20453 20995
rect 20453 20961 20487 20995
rect 20487 20961 20496 20995
rect 20444 20952 20496 20961
rect 22008 20952 22060 21004
rect 25780 20995 25832 21004
rect 7564 20884 7616 20936
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 11980 20884 12032 20936
rect 19984 20884 20036 20936
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 25780 20961 25789 20995
rect 25789 20961 25823 20995
rect 25823 20961 25832 20995
rect 25780 20952 25832 20961
rect 28724 20952 28776 21004
rect 23664 20884 23716 20936
rect 24860 20884 24912 20936
rect 9956 20816 10008 20868
rect 18696 20859 18748 20868
rect 18696 20825 18705 20859
rect 18705 20825 18739 20859
rect 18739 20825 18748 20859
rect 18696 20816 18748 20825
rect 21180 20816 21232 20868
rect 22192 20816 22244 20868
rect 25504 20816 25556 20868
rect 26792 20816 26844 20868
rect 27528 20816 27580 20868
rect 28632 20816 28684 20868
rect 45284 21088 45336 21140
rect 30196 20952 30248 21004
rect 30472 20995 30524 21004
rect 30472 20961 30481 20995
rect 30481 20961 30515 20995
rect 30515 20961 30524 20995
rect 30472 20952 30524 20961
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 45468 20884 45520 20936
rect 46296 20927 46348 20936
rect 46296 20893 46305 20927
rect 46305 20893 46339 20927
rect 46339 20893 46348 20927
rect 46296 20884 46348 20893
rect 10048 20748 10100 20800
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 20260 20748 20312 20800
rect 23204 20748 23256 20800
rect 24492 20791 24544 20800
rect 24492 20757 24501 20791
rect 24501 20757 24535 20791
rect 24535 20757 24544 20791
rect 24492 20748 24544 20757
rect 45836 20816 45888 20868
rect 47308 20816 47360 20868
rect 32588 20748 32640 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3516 20544 3568 20596
rect 25228 20544 25280 20596
rect 25412 20544 25464 20596
rect 33784 20544 33836 20596
rect 44456 20544 44508 20596
rect 47676 20587 47728 20596
rect 3424 20476 3476 20528
rect 9956 20519 10008 20528
rect 7564 20451 7616 20460
rect 7564 20417 7573 20451
rect 7573 20417 7607 20451
rect 7607 20417 7616 20451
rect 7564 20408 7616 20417
rect 7932 20340 7984 20392
rect 9956 20485 9965 20519
rect 9965 20485 9999 20519
rect 9999 20485 10008 20519
rect 9956 20476 10008 20485
rect 15016 20476 15068 20528
rect 19340 20476 19392 20528
rect 24492 20476 24544 20528
rect 28816 20476 28868 20528
rect 45376 20519 45428 20528
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 10692 20451 10744 20460
rect 9864 20408 9916 20417
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12624 20451 12676 20460
rect 12624 20417 12633 20451
rect 12633 20417 12667 20451
rect 12667 20417 12676 20451
rect 12624 20408 12676 20417
rect 17408 20408 17460 20460
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 19984 20408 20036 20460
rect 22560 20451 22612 20460
rect 12808 20383 12860 20392
rect 4804 20204 4856 20256
rect 10876 20272 10928 20324
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 16580 20340 16632 20392
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 22836 20408 22888 20460
rect 23204 20451 23256 20460
rect 23204 20417 23213 20451
rect 23213 20417 23247 20451
rect 23247 20417 23256 20451
rect 23204 20408 23256 20417
rect 26792 20408 26844 20460
rect 27252 20408 27304 20460
rect 11980 20247 12032 20256
rect 11980 20213 11989 20247
rect 11989 20213 12023 20247
rect 12023 20213 12032 20247
rect 11980 20204 12032 20213
rect 16672 20204 16724 20256
rect 16948 20204 17000 20256
rect 19708 20204 19760 20256
rect 22468 20204 22520 20256
rect 25504 20340 25556 20392
rect 27712 20383 27764 20392
rect 27712 20349 27721 20383
rect 27721 20349 27755 20383
rect 27755 20349 27764 20383
rect 27712 20340 27764 20349
rect 25228 20272 25280 20324
rect 25136 20204 25188 20256
rect 26148 20247 26200 20256
rect 26148 20213 26157 20247
rect 26157 20213 26191 20247
rect 26191 20213 26200 20247
rect 26148 20204 26200 20213
rect 26792 20204 26844 20256
rect 27252 20204 27304 20256
rect 45376 20485 45385 20519
rect 45385 20485 45419 20519
rect 45419 20485 45428 20519
rect 45376 20476 45428 20485
rect 47676 20553 47685 20587
rect 47685 20553 47719 20587
rect 47719 20553 47728 20587
rect 47676 20544 47728 20553
rect 47860 20476 47912 20528
rect 43812 20451 43864 20460
rect 43812 20417 43821 20451
rect 43821 20417 43855 20451
rect 43855 20417 43864 20451
rect 43812 20408 43864 20417
rect 44180 20451 44232 20460
rect 44180 20417 44189 20451
rect 44189 20417 44223 20451
rect 44223 20417 44232 20451
rect 44180 20408 44232 20417
rect 45100 20408 45152 20460
rect 47584 20451 47636 20460
rect 33784 20340 33836 20392
rect 44456 20340 44508 20392
rect 44640 20383 44692 20392
rect 44640 20349 44649 20383
rect 44649 20349 44683 20383
rect 44683 20349 44692 20383
rect 44640 20340 44692 20349
rect 47584 20417 47593 20451
rect 47593 20417 47627 20451
rect 47627 20417 47636 20451
rect 47584 20408 47636 20417
rect 46664 20383 46716 20392
rect 46664 20349 46673 20383
rect 46673 20349 46707 20383
rect 46707 20349 46716 20383
rect 46664 20340 46716 20349
rect 40776 20272 40828 20324
rect 44272 20272 44324 20324
rect 44364 20272 44416 20324
rect 45376 20272 45428 20324
rect 40684 20204 40736 20256
rect 46020 20204 46072 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7932 20043 7984 20052
rect 7932 20009 7941 20043
rect 7941 20009 7975 20043
rect 7975 20009 7984 20043
rect 7932 20000 7984 20009
rect 8944 20043 8996 20052
rect 8944 20009 8953 20043
rect 8953 20009 8987 20043
rect 8987 20009 8996 20043
rect 8944 20000 8996 20009
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 3792 19932 3844 19984
rect 28540 20000 28592 20052
rect 44272 20000 44324 20052
rect 47584 20000 47636 20052
rect 18236 19932 18288 19984
rect 19432 19932 19484 19984
rect 1768 19796 1820 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 13728 19864 13780 19916
rect 16396 19907 16448 19916
rect 15016 19796 15068 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 20260 19932 20312 19984
rect 22468 19932 22520 19984
rect 25136 19975 25188 19984
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 18236 19771 18288 19780
rect 18236 19737 18245 19771
rect 18245 19737 18279 19771
rect 18279 19737 18288 19771
rect 18236 19728 18288 19737
rect 22652 19864 22704 19916
rect 23020 19864 23072 19916
rect 23388 19864 23440 19916
rect 25136 19941 25145 19975
rect 25145 19941 25179 19975
rect 25179 19941 25188 19975
rect 25136 19932 25188 19941
rect 26516 19932 26568 19984
rect 27988 19864 28040 19916
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 23664 19839 23716 19848
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 24308 19796 24360 19848
rect 25780 19796 25832 19848
rect 27252 19796 27304 19848
rect 28816 19839 28868 19848
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 23296 19728 23348 19780
rect 24860 19728 24912 19780
rect 26516 19771 26568 19780
rect 26516 19737 26525 19771
rect 26525 19737 26559 19771
rect 26559 19737 26568 19771
rect 26516 19728 26568 19737
rect 27804 19728 27856 19780
rect 17408 19660 17460 19712
rect 18144 19660 18196 19712
rect 19432 19660 19484 19712
rect 23112 19660 23164 19712
rect 23848 19660 23900 19712
rect 23940 19660 23992 19712
rect 27712 19660 27764 19712
rect 28908 19660 28960 19712
rect 40684 19728 40736 19780
rect 40960 19771 41012 19780
rect 40960 19737 40969 19771
rect 40969 19737 41003 19771
rect 41003 19737 41012 19771
rect 40960 19728 41012 19737
rect 42616 19771 42668 19780
rect 42616 19737 42625 19771
rect 42625 19737 42659 19771
rect 42659 19737 42668 19771
rect 42616 19728 42668 19737
rect 44640 19932 44692 19984
rect 45376 19975 45428 19984
rect 45376 19941 45385 19975
rect 45385 19941 45419 19975
rect 45419 19941 45428 19975
rect 45376 19932 45428 19941
rect 48044 19864 48096 19916
rect 43996 19796 44048 19848
rect 43444 19660 43496 19712
rect 43904 19728 43956 19780
rect 46664 19728 46716 19780
rect 45100 19660 45152 19712
rect 45560 19660 45612 19712
rect 47032 19660 47084 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 15200 19456 15252 19508
rect 23020 19456 23072 19508
rect 8300 19388 8352 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 8392 19252 8444 19304
rect 3056 19184 3108 19236
rect 8484 19184 8536 19236
rect 20 19116 72 19168
rect 9128 19252 9180 19304
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 12808 19320 12860 19372
rect 13452 19320 13504 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 18512 19388 18564 19440
rect 19156 19388 19208 19440
rect 19432 19388 19484 19440
rect 26148 19456 26200 19508
rect 40960 19456 41012 19508
rect 43812 19456 43864 19508
rect 23388 19431 23440 19440
rect 23388 19397 23397 19431
rect 23397 19397 23431 19431
rect 23431 19397 23440 19431
rect 23388 19388 23440 19397
rect 23848 19388 23900 19440
rect 27160 19431 27212 19440
rect 27160 19397 27169 19431
rect 27169 19397 27203 19431
rect 27203 19397 27212 19431
rect 27160 19388 27212 19397
rect 27436 19388 27488 19440
rect 30288 19388 30340 19440
rect 19340 19320 19392 19372
rect 21824 19320 21876 19372
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 25780 19363 25832 19372
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 25872 19320 25924 19372
rect 28356 19363 28408 19372
rect 28356 19329 28365 19363
rect 28365 19329 28399 19363
rect 28399 19329 28408 19363
rect 28356 19320 28408 19329
rect 28540 19363 28592 19372
rect 28540 19329 28549 19363
rect 28549 19329 28583 19363
rect 28583 19329 28592 19363
rect 28540 19320 28592 19329
rect 29828 19320 29880 19372
rect 11980 19252 12032 19304
rect 13544 19252 13596 19304
rect 13728 19252 13780 19304
rect 17592 19295 17644 19304
rect 17592 19261 17601 19295
rect 17601 19261 17635 19295
rect 17635 19261 17644 19295
rect 17592 19252 17644 19261
rect 8668 19184 8720 19236
rect 24860 19227 24912 19236
rect 24860 19193 24869 19227
rect 24869 19193 24903 19227
rect 24903 19193 24912 19227
rect 24860 19184 24912 19193
rect 28816 19252 28868 19304
rect 29736 19295 29788 19304
rect 29736 19261 29745 19295
rect 29745 19261 29779 19295
rect 29779 19261 29788 19295
rect 29736 19252 29788 19261
rect 30196 19295 30248 19304
rect 30196 19261 30205 19295
rect 30205 19261 30239 19295
rect 30239 19261 30248 19295
rect 30196 19252 30248 19261
rect 31392 19320 31444 19372
rect 40776 19363 40828 19372
rect 40776 19329 40785 19363
rect 40785 19329 40819 19363
rect 40819 19329 40828 19363
rect 40776 19320 40828 19329
rect 42984 19320 43036 19372
rect 44916 19388 44968 19440
rect 45376 19456 45428 19508
rect 47308 19456 47360 19508
rect 47032 19388 47084 19440
rect 45100 19295 45152 19304
rect 45100 19261 45109 19295
rect 45109 19261 45143 19295
rect 45143 19261 45152 19295
rect 45100 19252 45152 19261
rect 45744 19252 45796 19304
rect 46388 19320 46440 19372
rect 46756 19320 46808 19372
rect 27896 19184 27948 19236
rect 30380 19184 30432 19236
rect 43444 19184 43496 19236
rect 46112 19184 46164 19236
rect 46296 19184 46348 19236
rect 9772 19116 9824 19168
rect 11244 19116 11296 19168
rect 11796 19116 11848 19168
rect 12808 19116 12860 19168
rect 13176 19116 13228 19168
rect 13360 19116 13412 19168
rect 18236 19116 18288 19168
rect 20260 19116 20312 19168
rect 21916 19116 21968 19168
rect 22652 19116 22704 19168
rect 29552 19116 29604 19168
rect 31208 19159 31260 19168
rect 31208 19125 31217 19159
rect 31217 19125 31251 19159
rect 31251 19125 31260 19159
rect 31208 19116 31260 19125
rect 32312 19116 32364 19168
rect 33508 19116 33560 19168
rect 43812 19116 43864 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 2044 18844 2096 18896
rect 16304 18912 16356 18964
rect 16580 18912 16632 18964
rect 30472 18912 30524 18964
rect 32128 18912 32180 18964
rect 43996 18912 44048 18964
rect 45100 18912 45152 18964
rect 18328 18887 18380 18896
rect 11796 18819 11848 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 11796 18785 11805 18819
rect 11805 18785 11839 18819
rect 11839 18785 11848 18819
rect 11796 18776 11848 18785
rect 2136 18708 2188 18717
rect 8116 18708 8168 18760
rect 9036 18708 9088 18760
rect 13176 18708 13228 18760
rect 15200 18776 15252 18828
rect 18328 18853 18337 18887
rect 18337 18853 18371 18887
rect 18371 18853 18380 18887
rect 18328 18844 18380 18853
rect 18420 18844 18472 18896
rect 19156 18844 19208 18896
rect 16488 18776 16540 18828
rect 22652 18844 22704 18896
rect 23020 18844 23072 18896
rect 20076 18776 20128 18828
rect 21916 18819 21968 18828
rect 21916 18785 21925 18819
rect 21925 18785 21959 18819
rect 21959 18785 21968 18819
rect 21916 18776 21968 18785
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 33508 18844 33560 18896
rect 9404 18683 9456 18692
rect 9404 18649 9413 18683
rect 9413 18649 9447 18683
rect 9447 18649 9456 18683
rect 9404 18640 9456 18649
rect 10784 18640 10836 18692
rect 8392 18572 8444 18624
rect 10232 18572 10284 18624
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 27068 18776 27120 18828
rect 29828 18819 29880 18828
rect 29828 18785 29837 18819
rect 29837 18785 29871 18819
rect 29871 18785 29880 18819
rect 29828 18776 29880 18785
rect 15660 18683 15712 18692
rect 15660 18649 15669 18683
rect 15669 18649 15703 18683
rect 15703 18649 15712 18683
rect 15660 18640 15712 18649
rect 13084 18572 13136 18624
rect 14280 18572 14332 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 18972 18640 19024 18692
rect 25780 18708 25832 18760
rect 26240 18708 26292 18760
rect 26976 18708 27028 18760
rect 27160 18751 27212 18760
rect 27160 18717 27169 18751
rect 27169 18717 27203 18751
rect 27203 18717 27212 18751
rect 27160 18708 27212 18717
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 27620 18708 27672 18760
rect 28540 18708 28592 18760
rect 18144 18572 18196 18624
rect 22192 18640 22244 18692
rect 25964 18683 26016 18692
rect 25964 18649 25973 18683
rect 25973 18649 26007 18683
rect 26007 18649 26016 18683
rect 25964 18640 26016 18649
rect 28356 18640 28408 18692
rect 29552 18708 29604 18760
rect 30288 18708 30340 18760
rect 30380 18751 30432 18760
rect 30380 18717 30389 18751
rect 30389 18717 30423 18751
rect 30423 18717 30432 18751
rect 30380 18708 30432 18717
rect 31208 18708 31260 18760
rect 25596 18572 25648 18624
rect 43812 18708 43864 18760
rect 45100 18776 45152 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 45008 18751 45060 18760
rect 45008 18717 45017 18751
rect 45017 18717 45051 18751
rect 45051 18717 45060 18751
rect 45008 18708 45060 18717
rect 45192 18751 45244 18760
rect 45192 18717 45201 18751
rect 45201 18717 45235 18751
rect 45235 18717 45244 18751
rect 45192 18708 45244 18717
rect 46296 18751 46348 18760
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 47676 18640 47728 18692
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 9404 18368 9456 18420
rect 8116 18300 8168 18352
rect 10692 18368 10744 18420
rect 10784 18368 10836 18420
rect 11520 18368 11572 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 12440 18368 12492 18420
rect 16396 18368 16448 18420
rect 17592 18368 17644 18420
rect 18144 18411 18196 18420
rect 18144 18377 18153 18411
rect 18153 18377 18187 18411
rect 18187 18377 18196 18411
rect 18144 18368 18196 18377
rect 25872 18368 25924 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 2412 18232 2464 18284
rect 8576 18232 8628 18284
rect 9128 18232 9180 18284
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 11336 18300 11388 18352
rect 16120 18343 16172 18352
rect 10232 18275 10284 18284
rect 10232 18241 10241 18275
rect 10241 18241 10275 18275
rect 10275 18241 10284 18275
rect 10232 18232 10284 18241
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 10876 18232 10928 18284
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11980 18232 12032 18284
rect 16120 18309 16129 18343
rect 16129 18309 16163 18343
rect 16163 18309 16172 18343
rect 16120 18300 16172 18309
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 18328 18300 18380 18352
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 17776 18232 17828 18284
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 15660 18164 15712 18216
rect 25228 18300 25280 18352
rect 29000 18300 29052 18352
rect 32312 18343 32364 18352
rect 32312 18309 32321 18343
rect 32321 18309 32355 18343
rect 32355 18309 32364 18343
rect 32312 18300 32364 18309
rect 20720 18232 20772 18284
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 25964 18232 26016 18284
rect 27068 18232 27120 18284
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 21272 18164 21324 18216
rect 26240 18164 26292 18216
rect 1952 18028 2004 18080
rect 8576 18028 8628 18080
rect 13268 18028 13320 18080
rect 13360 18028 13412 18080
rect 16764 18028 16816 18080
rect 20812 18071 20864 18080
rect 20812 18037 20821 18071
rect 20821 18037 20855 18071
rect 20855 18037 20864 18071
rect 20812 18028 20864 18037
rect 20904 18028 20956 18080
rect 27804 18164 27856 18216
rect 27896 18207 27948 18216
rect 27896 18173 27905 18207
rect 27905 18173 27939 18207
rect 27939 18173 27948 18207
rect 27896 18164 27948 18173
rect 30196 18164 30248 18216
rect 31484 18207 31536 18216
rect 31484 18173 31493 18207
rect 31493 18173 31527 18207
rect 31527 18173 31536 18207
rect 31484 18164 31536 18173
rect 33968 18207 34020 18216
rect 33968 18173 33977 18207
rect 33977 18173 34011 18207
rect 34011 18173 34020 18207
rect 33968 18164 34020 18173
rect 28172 18096 28224 18148
rect 28264 18028 28316 18080
rect 47676 18411 47728 18420
rect 43812 18232 43864 18284
rect 44916 18300 44968 18352
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 45100 18232 45152 18284
rect 45928 18275 45980 18284
rect 45928 18241 45937 18275
rect 45937 18241 45971 18275
rect 45971 18241 45980 18275
rect 45928 18232 45980 18241
rect 44456 18164 44508 18216
rect 46296 18232 46348 18284
rect 47400 18232 47452 18284
rect 44640 18096 44692 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3056 17824 3108 17876
rect 13728 17824 13780 17876
rect 14464 17824 14516 17876
rect 21272 17824 21324 17876
rect 27620 17824 27672 17876
rect 27804 17867 27856 17876
rect 27804 17833 27813 17867
rect 27813 17833 27847 17867
rect 27847 17833 27856 17867
rect 27804 17824 27856 17833
rect 28264 17824 28316 17876
rect 28448 17824 28500 17876
rect 29000 17824 29052 17876
rect 29736 17824 29788 17876
rect 44456 17867 44508 17876
rect 44456 17833 44465 17867
rect 44465 17833 44499 17867
rect 44499 17833 44508 17867
rect 44456 17824 44508 17833
rect 45100 17824 45152 17876
rect 11704 17756 11756 17808
rect 16396 17756 16448 17808
rect 3700 17688 3752 17740
rect 1768 17620 1820 17672
rect 11152 17620 11204 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11520 17552 11572 17604
rect 13176 17620 13228 17672
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 17776 17620 17828 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 12072 17595 12124 17604
rect 11612 17484 11664 17536
rect 12072 17561 12081 17595
rect 12081 17561 12115 17595
rect 12115 17561 12124 17595
rect 12072 17552 12124 17561
rect 15108 17552 15160 17604
rect 13360 17484 13412 17536
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 16396 17484 16448 17536
rect 16856 17484 16908 17536
rect 20904 17595 20956 17604
rect 20904 17561 20913 17595
rect 20913 17561 20947 17595
rect 20947 17561 20956 17595
rect 20904 17552 20956 17561
rect 21180 17484 21232 17536
rect 21272 17484 21324 17536
rect 24676 17688 24728 17740
rect 25596 17731 25648 17740
rect 25596 17697 25605 17731
rect 25605 17697 25639 17731
rect 25639 17697 25648 17731
rect 25596 17688 25648 17697
rect 26148 17688 26200 17740
rect 26240 17688 26292 17740
rect 30288 17756 30340 17808
rect 22928 17620 22980 17672
rect 23112 17620 23164 17672
rect 25504 17620 25556 17672
rect 22192 17552 22244 17604
rect 23480 17552 23532 17604
rect 27988 17620 28040 17672
rect 29552 17663 29604 17672
rect 29552 17629 29561 17663
rect 29561 17629 29595 17663
rect 29595 17629 29604 17663
rect 29552 17620 29604 17629
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 23940 17484 23992 17536
rect 43536 17620 43588 17672
rect 44272 17663 44324 17672
rect 44272 17629 44281 17663
rect 44281 17629 44315 17663
rect 44315 17629 44324 17663
rect 44272 17620 44324 17629
rect 46296 17663 46348 17672
rect 46296 17629 46305 17663
rect 46305 17629 46339 17663
rect 46339 17629 46348 17663
rect 46296 17620 46348 17629
rect 44456 17552 44508 17604
rect 45008 17595 45060 17604
rect 45008 17561 45017 17595
rect 45017 17561 45051 17595
rect 45051 17561 45060 17595
rect 45008 17552 45060 17561
rect 45192 17595 45244 17604
rect 45192 17561 45201 17595
rect 45201 17561 45235 17595
rect 45235 17561 45244 17595
rect 45192 17552 45244 17561
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 44824 17484 44876 17536
rect 47400 17484 47452 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 12624 17280 12676 17332
rect 13176 17323 13228 17332
rect 13176 17289 13185 17323
rect 13185 17289 13219 17323
rect 13219 17289 13228 17323
rect 13176 17280 13228 17289
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 23112 17323 23164 17332
rect 23112 17289 23137 17323
rect 23137 17289 23164 17323
rect 23112 17280 23164 17289
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 11152 17212 11204 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 11612 17212 11664 17264
rect 11980 17144 12032 17196
rect 12440 17144 12492 17196
rect 18604 17212 18656 17264
rect 20720 17212 20772 17264
rect 23480 17212 23532 17264
rect 23940 17255 23992 17264
rect 12716 17144 12768 17196
rect 12808 17144 12860 17196
rect 13176 17144 13228 17196
rect 14004 17144 14056 17196
rect 14556 17144 14608 17196
rect 14648 17144 14700 17196
rect 15108 17144 15160 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 23848 17144 23900 17196
rect 24676 17280 24728 17332
rect 27252 17280 27304 17332
rect 45008 17280 45060 17332
rect 47676 17323 47728 17332
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 45928 17212 45980 17264
rect 46296 17212 46348 17264
rect 26976 17187 27028 17196
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 2964 17076 3016 17128
rect 15936 17119 15988 17128
rect 15936 17085 15945 17119
rect 15945 17085 15979 17119
rect 15979 17085 15988 17119
rect 15936 17076 15988 17085
rect 18328 17076 18380 17128
rect 18512 17076 18564 17128
rect 19432 17119 19484 17128
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 21088 17076 21140 17128
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 27436 17144 27488 17196
rect 44272 17187 44324 17196
rect 44272 17153 44281 17187
rect 44281 17153 44315 17187
rect 44315 17153 44324 17187
rect 44272 17144 44324 17153
rect 44456 17187 44508 17196
rect 44456 17153 44465 17187
rect 44465 17153 44499 17187
rect 44499 17153 44508 17187
rect 44456 17144 44508 17153
rect 46388 17187 46440 17196
rect 46388 17153 46397 17187
rect 46397 17153 46431 17187
rect 46431 17153 46440 17187
rect 46388 17144 46440 17153
rect 47400 17144 47452 17196
rect 46204 17076 46256 17128
rect 20812 17008 20864 17060
rect 11612 16940 11664 16992
rect 12164 16940 12216 16992
rect 12348 16983 12400 16992
rect 12348 16949 12357 16983
rect 12357 16949 12391 16983
rect 12391 16949 12400 16983
rect 12348 16940 12400 16949
rect 14556 16940 14608 16992
rect 19064 16940 19116 16992
rect 21272 16940 21324 16992
rect 23204 17008 23256 17060
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 23756 16983 23808 16992
rect 23756 16949 23765 16983
rect 23765 16949 23799 16983
rect 23799 16949 23808 16983
rect 23756 16940 23808 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 12072 16736 12124 16788
rect 17776 16736 17828 16788
rect 19432 16736 19484 16788
rect 11980 16668 12032 16720
rect 13544 16668 13596 16720
rect 12348 16600 12400 16652
rect 12624 16600 12676 16652
rect 15936 16668 15988 16720
rect 47032 16736 47084 16788
rect 20628 16668 20680 16720
rect 21088 16668 21140 16720
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 16948 16532 17000 16584
rect 19064 16600 19116 16652
rect 23296 16668 23348 16720
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 19248 16532 19300 16584
rect 20260 16532 20312 16584
rect 20720 16532 20772 16584
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 22192 16532 22244 16584
rect 22652 16532 22704 16584
rect 22836 16575 22888 16584
rect 22836 16541 22837 16575
rect 22837 16541 22871 16575
rect 22871 16541 22888 16575
rect 22836 16532 22888 16541
rect 23756 16600 23808 16652
rect 23940 16600 23992 16652
rect 24676 16600 24728 16652
rect 27528 16643 27580 16652
rect 27528 16609 27537 16643
rect 27537 16609 27571 16643
rect 27571 16609 27580 16643
rect 27528 16600 27580 16609
rect 28632 16600 28684 16652
rect 24308 16532 24360 16584
rect 47768 16600 47820 16652
rect 29552 16575 29604 16584
rect 29552 16541 29561 16575
rect 29561 16541 29595 16575
rect 29595 16541 29604 16575
rect 29552 16532 29604 16541
rect 38660 16532 38712 16584
rect 26056 16507 26108 16516
rect 17592 16439 17644 16448
rect 17592 16405 17601 16439
rect 17601 16405 17635 16439
rect 17635 16405 17644 16439
rect 17592 16396 17644 16405
rect 22836 16396 22888 16448
rect 22928 16439 22980 16448
rect 22928 16405 22937 16439
rect 22937 16405 22971 16439
rect 22971 16405 22980 16439
rect 23572 16439 23624 16448
rect 22928 16396 22980 16405
rect 23572 16405 23581 16439
rect 23581 16405 23615 16439
rect 23615 16405 23624 16439
rect 23572 16396 23624 16405
rect 24492 16439 24544 16448
rect 24492 16405 24501 16439
rect 24501 16405 24535 16439
rect 24535 16405 24544 16439
rect 24492 16396 24544 16405
rect 26056 16473 26065 16507
rect 26065 16473 26099 16507
rect 26099 16473 26108 16507
rect 26056 16464 26108 16473
rect 45560 16464 45612 16516
rect 46848 16464 46900 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 13176 16056 13228 16108
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 16948 16192 17000 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 18420 16192 18472 16244
rect 24492 16124 24544 16176
rect 25320 16192 25372 16244
rect 46848 16235 46900 16244
rect 16580 16056 16632 16108
rect 16948 16056 17000 16108
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 19248 16056 19300 16108
rect 21180 16056 21232 16108
rect 22836 16099 22888 16108
rect 22836 16065 22845 16099
rect 22845 16065 22879 16099
rect 22879 16065 22888 16099
rect 22836 16056 22888 16065
rect 25228 16099 25280 16108
rect 25228 16065 25237 16099
rect 25237 16065 25271 16099
rect 25271 16065 25280 16099
rect 38200 16124 38252 16176
rect 25964 16099 26016 16108
rect 25228 16056 25280 16065
rect 25964 16065 25973 16099
rect 25973 16065 26007 16099
rect 26007 16065 26016 16099
rect 25964 16056 26016 16065
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 28172 16099 28224 16108
rect 26056 16056 26108 16065
rect 28172 16065 28181 16099
rect 28181 16065 28215 16099
rect 28215 16065 28224 16099
rect 28172 16056 28224 16065
rect 30472 16056 30524 16108
rect 46848 16201 46857 16235
rect 46857 16201 46891 16235
rect 46891 16201 46900 16235
rect 46848 16192 46900 16201
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 17132 15988 17184 16040
rect 23572 15988 23624 16040
rect 24676 15988 24728 16040
rect 28448 15988 28500 16040
rect 16764 15920 16816 15972
rect 19248 15920 19300 15972
rect 11060 15852 11112 15904
rect 12348 15895 12400 15904
rect 12348 15861 12357 15895
rect 12357 15861 12391 15895
rect 12391 15861 12400 15895
rect 12348 15852 12400 15861
rect 14004 15852 14056 15904
rect 16396 15852 16448 15904
rect 18420 15852 18472 15904
rect 19340 15852 19392 15904
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 25320 15895 25372 15904
rect 25320 15861 25329 15895
rect 25329 15861 25363 15895
rect 25363 15861 25372 15895
rect 25320 15852 25372 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 12716 15648 12768 15700
rect 17592 15648 17644 15700
rect 22652 15648 22704 15700
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 29552 15580 29604 15632
rect 11796 15512 11848 15564
rect 12072 15512 12124 15564
rect 16948 15512 17000 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 22376 15512 22428 15564
rect 1768 15444 1820 15496
rect 12348 15444 12400 15496
rect 15200 15444 15252 15496
rect 15752 15444 15804 15496
rect 16764 15376 16816 15428
rect 17040 15376 17092 15428
rect 17776 15444 17828 15496
rect 22928 15512 22980 15564
rect 25320 15555 25372 15564
rect 25320 15521 25329 15555
rect 25329 15521 25363 15555
rect 25363 15521 25372 15555
rect 25320 15512 25372 15521
rect 26700 15555 26752 15564
rect 26700 15521 26709 15555
rect 26709 15521 26743 15555
rect 26743 15521 26752 15555
rect 26700 15512 26752 15521
rect 12072 15308 12124 15360
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 17960 15308 18012 15360
rect 18052 15308 18104 15360
rect 19984 15308 20036 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 15292 15036 15344 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 12256 14968 12308 15020
rect 12900 14968 12952 15020
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 18512 15104 18564 15156
rect 19984 15104 20036 15156
rect 16948 15036 17000 15088
rect 17960 15036 18012 15088
rect 19340 15036 19392 15088
rect 15200 14968 15252 14977
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 17132 14943 17184 14952
rect 11428 14764 11480 14816
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 14924 14832 14976 14884
rect 16580 14832 16632 14884
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17132 14900 17184 14909
rect 15108 14764 15160 14816
rect 16028 14764 16080 14816
rect 17224 14764 17276 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 14924 14492 14976 14544
rect 17132 14560 17184 14612
rect 16120 14492 16172 14544
rect 17040 14492 17092 14544
rect 17224 14535 17276 14544
rect 17224 14501 17233 14535
rect 17233 14501 17267 14535
rect 17267 14501 17276 14535
rect 17224 14492 17276 14501
rect 27712 14424 27764 14476
rect 2136 14356 2188 14365
rect 16028 14356 16080 14408
rect 16856 14356 16908 14408
rect 11704 14331 11756 14340
rect 11704 14297 11713 14331
rect 11713 14297 11747 14331
rect 11747 14297 11756 14331
rect 11704 14288 11756 14297
rect 13268 14288 13320 14340
rect 14280 14288 14332 14340
rect 14924 14331 14976 14340
rect 14924 14297 14933 14331
rect 14933 14297 14967 14331
rect 14967 14297 14976 14331
rect 14924 14288 14976 14297
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 15844 14288 15896 14340
rect 16120 14331 16172 14340
rect 16120 14297 16129 14331
rect 16129 14297 16163 14331
rect 16163 14297 16172 14331
rect 16120 14288 16172 14297
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 15108 14220 15160 14272
rect 15384 14220 15436 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 20628 14356 20680 14408
rect 16488 14220 16540 14229
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 18420 14220 18472 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 11704 14016 11756 14068
rect 15200 14016 15252 14068
rect 17132 14016 17184 14068
rect 12716 13948 12768 14000
rect 12440 13880 12492 13932
rect 11704 13812 11756 13864
rect 13176 13880 13228 13932
rect 14556 13948 14608 14000
rect 17868 13948 17920 14000
rect 18604 13948 18656 14000
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 3424 13744 3476 13796
rect 15476 13744 15528 13796
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14556 13472 14608 13524
rect 15752 13472 15804 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 17316 13472 17368 13524
rect 18604 13472 18656 13524
rect 12440 13404 12492 13456
rect 17776 13268 17828 13320
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 13912 13200 13964 13252
rect 15476 13243 15528 13252
rect 15476 13209 15485 13243
rect 15485 13209 15519 13243
rect 15519 13209 15528 13243
rect 15476 13200 15528 13209
rect 16120 13200 16172 13252
rect 12624 13175 12676 13184
rect 12624 13141 12659 13175
rect 12659 13141 12676 13175
rect 12624 13132 12676 13141
rect 15384 13132 15436 13184
rect 16672 13175 16724 13184
rect 16672 13141 16681 13175
rect 16681 13141 16715 13175
rect 16715 13141 16724 13175
rect 16672 13132 16724 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 27620 12928 27672 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 14188 12792 14240 12844
rect 15292 12792 15344 12844
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 12624 12724 12676 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 15016 12588 15068 12640
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 47768 12631 47820 12640
rect 47768 12597 47777 12631
rect 47777 12597 47811 12631
rect 47811 12597 47820 12631
rect 47768 12588 47820 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12808 12384 12860 12436
rect 14188 12427 14240 12436
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 12256 12180 12308 12232
rect 15844 12248 15896 12300
rect 16488 12248 16540 12300
rect 16672 12248 16724 12300
rect 47768 12248 47820 12300
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15384 12180 15436 12232
rect 15752 12180 15804 12232
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 18052 12112 18104 12164
rect 47676 12112 47728 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 18052 11840 18104 11892
rect 47676 11883 47728 11892
rect 47676 11849 47685 11883
rect 47685 11849 47719 11883
rect 47719 11849 47728 11883
rect 47676 11840 47728 11849
rect 15476 11772 15528 11824
rect 16580 11772 16632 11824
rect 12256 11747 12308 11756
rect 12256 11713 12265 11747
rect 12265 11713 12299 11747
rect 12299 11713 12308 11747
rect 12256 11704 12308 11713
rect 12624 11704 12676 11756
rect 14096 11704 14148 11756
rect 15016 11636 15068 11688
rect 15384 11704 15436 11756
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 18420 11704 18472 11756
rect 25596 11704 25648 11756
rect 25964 11704 26016 11756
rect 28632 11636 28684 11688
rect 15292 11568 15344 11620
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 46480 11500 46532 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12900 11160 12952 11212
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 16580 11160 16632 11212
rect 46480 11203 46532 11212
rect 46480 11169 46489 11203
rect 46489 11169 46523 11203
rect 46523 11169 46532 11203
rect 46480 11160 46532 11169
rect 13912 11092 13964 11144
rect 16764 11092 16816 11144
rect 47768 11024 47820 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 3516 10956 3568 11008
rect 4804 10956 4856 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 12440 10684 12492 10736
rect 13820 10684 13872 10736
rect 14648 10684 14700 10736
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 15108 10523 15160 10532
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 46388 10548 46440 10600
rect 46756 10591 46808 10600
rect 46756 10557 46765 10591
rect 46765 10557 46799 10591
rect 46799 10557 46808 10591
rect 46756 10548 46808 10557
rect 45652 10480 45704 10532
rect 13912 10412 13964 10464
rect 14096 10412 14148 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 47032 10072 47084 10124
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 13820 10004 13872 10056
rect 14924 10004 14976 10056
rect 16764 9936 16816 9988
rect 25872 9936 25924 9988
rect 47676 9936 47728 9988
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 11796 9528 11848 9580
rect 14004 9596 14056 9648
rect 13820 9528 13872 9580
rect 14464 9639 14516 9648
rect 14464 9605 14473 9639
rect 14473 9605 14507 9639
rect 14507 9605 14516 9639
rect 14464 9596 14516 9605
rect 15384 9664 15436 9716
rect 15108 9596 15160 9648
rect 16764 9639 16816 9648
rect 16764 9605 16773 9639
rect 16773 9605 16807 9639
rect 16807 9605 16816 9639
rect 16764 9596 16816 9605
rect 47676 9639 47728 9648
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 47032 9571 47084 9580
rect 47032 9537 47041 9571
rect 47041 9537 47075 9571
rect 47075 9537 47084 9571
rect 47032 9528 47084 9537
rect 47492 9528 47544 9580
rect 13636 9392 13688 9444
rect 11888 9324 11940 9376
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 12072 9052 12124 9104
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 13544 8891 13596 8900
rect 13544 8857 13553 8891
rect 13553 8857 13587 8891
rect 13587 8857 13596 8891
rect 13544 8848 13596 8857
rect 3792 8780 3844 8832
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 17960 9027 18012 9036
rect 17960 8993 17969 9027
rect 17969 8993 18003 9027
rect 18003 8993 18012 9027
rect 17960 8984 18012 8993
rect 46848 8984 46900 9036
rect 46388 8916 46440 8968
rect 14464 8891 14516 8900
rect 14464 8857 14473 8891
rect 14473 8857 14507 8891
rect 14507 8857 14516 8891
rect 14464 8848 14516 8857
rect 16764 8891 16816 8900
rect 16764 8857 16773 8891
rect 16773 8857 16807 8891
rect 16807 8857 16816 8891
rect 16764 8848 16816 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 13728 8508 13780 8560
rect 47768 8551 47820 8560
rect 47768 8517 47777 8551
rect 47777 8517 47811 8551
rect 47811 8517 47820 8551
rect 47768 8508 47820 8517
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 14832 8415 14884 8424
rect 4068 8236 4120 8288
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 42708 8372 42760 8424
rect 46940 8372 46992 8424
rect 24768 8304 24820 8356
rect 13544 8236 13596 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11888 8032 11940 8084
rect 14464 8032 14516 8084
rect 16764 8032 16816 8084
rect 46572 7896 46624 7948
rect 46664 7896 46716 7948
rect 10416 7828 10468 7880
rect 11796 7828 11848 7880
rect 13820 7828 13872 7880
rect 47492 7760 47544 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1676 7420 1728 7472
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 45192 7327 45244 7336
rect 45192 7293 45201 7327
rect 45201 7293 45235 7327
rect 45235 7293 45244 7327
rect 45192 7284 45244 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6808 4120 6860
rect 17960 6808 18012 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47492 6808 47544 6860
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 48136 6307 48188 6316
rect 48136 6273 48145 6307
rect 48145 6273 48179 6307
rect 48179 6273 48188 6307
rect 48136 6264 48188 6273
rect 14372 6128 14424 6180
rect 32220 6128 32272 6180
rect 47952 6103 48004 6112
rect 47952 6069 47961 6103
rect 47961 6069 47995 6103
rect 47995 6069 48004 6103
rect 47952 6060 48004 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 46848 5720 46900 5772
rect 46204 5652 46256 5704
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 47952 5244 48004 5296
rect 18144 5176 18196 5228
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 21364 5176 21416 5228
rect 47860 5219 47912 5228
rect 47860 5185 47869 5219
rect 47869 5185 47903 5219
rect 47903 5185 47912 5219
rect 47860 5176 47912 5185
rect 45652 5108 45704 5160
rect 45192 5040 45244 5092
rect 17592 4972 17644 5024
rect 20720 4972 20772 5024
rect 21916 4972 21968 5024
rect 32772 4972 32824 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20076 4768 20128 4820
rect 21364 4811 21416 4820
rect 21364 4777 21373 4811
rect 21373 4777 21407 4811
rect 21407 4777 21416 4811
rect 21364 4768 21416 4777
rect 31484 4768 31536 4820
rect 45100 4768 45152 4820
rect 45836 4768 45888 4820
rect 6920 4632 6972 4684
rect 9404 4564 9456 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 19892 4564 19944 4616
rect 20904 4632 20956 4684
rect 45652 4632 45704 4684
rect 46296 4675 46348 4684
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 20720 4564 20772 4616
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 42892 4607 42944 4616
rect 42892 4573 42901 4607
rect 42901 4573 42935 4607
rect 42935 4573 42944 4607
rect 42892 4564 42944 4573
rect 45192 4564 45244 4616
rect 15568 4496 15620 4548
rect 43996 4496 44048 4548
rect 46020 4539 46072 4548
rect 46020 4505 46029 4539
rect 46029 4505 46063 4539
rect 46063 4505 46072 4539
rect 46020 4496 46072 4505
rect 17040 4428 17092 4480
rect 20720 4428 20772 4480
rect 23020 4428 23072 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 11520 4224 11572 4276
rect 18236 4224 18288 4276
rect 41328 4224 41380 4276
rect 10416 4131 10468 4140
rect 3148 4020 3200 4072
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 7104 4063 7156 4072
rect 3240 4020 3292 4029
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8208 4020 8260 4072
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 16672 4156 16724 4208
rect 16856 4088 16908 4140
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17776 4088 17828 4140
rect 18512 4088 18564 4140
rect 19340 4088 19392 4140
rect 20812 4131 20864 4140
rect 3884 3952 3936 4004
rect 7196 3952 7248 4004
rect 15660 4020 15712 4072
rect 19248 4020 19300 4072
rect 20812 4097 20821 4131
rect 20821 4097 20855 4131
rect 20855 4097 20864 4131
rect 20812 4088 20864 4097
rect 23112 4088 23164 4140
rect 25596 4088 25648 4140
rect 25780 4088 25832 4140
rect 30932 4088 30984 4140
rect 39764 4131 39816 4140
rect 39764 4097 39773 4131
rect 39773 4097 39807 4131
rect 39807 4097 39816 4131
rect 39764 4088 39816 4097
rect 42708 4156 42760 4208
rect 45652 4156 45704 4208
rect 46112 4131 46164 4140
rect 46112 4097 46121 4131
rect 46121 4097 46155 4131
rect 46155 4097 46164 4131
rect 46112 4088 46164 4097
rect 46664 4088 46716 4140
rect 46848 4088 46900 4140
rect 3976 3884 4028 3936
rect 10048 3952 10100 4004
rect 17224 3952 17276 4004
rect 30012 4020 30064 4072
rect 31392 4063 31444 4072
rect 31392 4029 31401 4063
rect 31401 4029 31435 4063
rect 31435 4029 31444 4063
rect 31392 4020 31444 4029
rect 36176 4020 36228 4072
rect 22744 3952 22796 4004
rect 36544 3952 36596 4004
rect 37832 3952 37884 4004
rect 43904 4020 43956 4072
rect 43996 4020 44048 4072
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9588 3884 9640 3936
rect 11704 3884 11756 3936
rect 14004 3884 14056 3936
rect 16948 3884 17000 3936
rect 17684 3884 17736 3936
rect 18328 3884 18380 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 19064 3927 19116 3936
rect 18420 3884 18472 3893
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 19432 3884 19484 3936
rect 20260 3884 20312 3936
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 23664 3884 23716 3936
rect 25320 3884 25372 3936
rect 25872 3884 25924 3936
rect 30840 3884 30892 3936
rect 33232 3927 33284 3936
rect 33232 3893 33241 3927
rect 33241 3893 33275 3927
rect 33275 3893 33284 3927
rect 33232 3884 33284 3893
rect 39856 3927 39908 3936
rect 39856 3893 39865 3927
rect 39865 3893 39899 3927
rect 39899 3893 39908 3927
rect 39856 3884 39908 3893
rect 42800 3884 42852 3936
rect 43536 3884 43588 3936
rect 46480 3884 46532 3936
rect 48044 3927 48096 3936
rect 48044 3893 48053 3927
rect 48053 3893 48087 3927
rect 48087 3893 48096 3927
rect 48044 3884 48096 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 3884 3680 3936 3732
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 1768 3476 1820 3528
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 9036 3612 9088 3664
rect 10048 3680 10100 3732
rect 17224 3680 17276 3732
rect 17776 3723 17828 3732
rect 17776 3689 17785 3723
rect 17785 3689 17819 3723
rect 17819 3689 17828 3723
rect 17776 3680 17828 3689
rect 18512 3680 18564 3732
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 20168 3680 20220 3732
rect 33968 3680 34020 3732
rect 36544 3680 36596 3732
rect 41236 3680 41288 3732
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 15108 3612 15160 3664
rect 42616 3680 42668 3732
rect 5816 3519 5868 3528
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 11520 3476 11572 3528
rect 13820 3476 13872 3528
rect 1952 3340 2004 3392
rect 4068 3340 4120 3392
rect 13636 3408 13688 3460
rect 7288 3340 7340 3392
rect 15384 3587 15436 3596
rect 15384 3553 15393 3587
rect 15393 3553 15427 3587
rect 15427 3553 15436 3587
rect 15384 3544 15436 3553
rect 16764 3476 16816 3528
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 18420 3476 18472 3528
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 20352 3544 20404 3596
rect 20812 3544 20864 3596
rect 25320 3587 25372 3596
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 22100 3476 22152 3528
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23664 3519 23716 3528
rect 23112 3476 23164 3485
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 21088 3408 21140 3460
rect 21180 3408 21232 3460
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 25412 3544 25464 3596
rect 27528 3544 27580 3596
rect 42524 3544 42576 3596
rect 42892 3612 42944 3664
rect 45652 3612 45704 3664
rect 47400 3612 47452 3664
rect 42800 3587 42852 3596
rect 42800 3553 42809 3587
rect 42809 3553 42843 3587
rect 42843 3553 42852 3587
rect 42800 3544 42852 3553
rect 43168 3587 43220 3596
rect 43168 3553 43177 3587
rect 43177 3553 43211 3587
rect 43211 3553 43220 3587
rect 43168 3544 43220 3553
rect 46480 3587 46532 3596
rect 33048 3476 33100 3528
rect 35992 3519 36044 3528
rect 35992 3485 36001 3519
rect 36001 3485 36035 3519
rect 36035 3485 36044 3519
rect 35992 3476 36044 3485
rect 37832 3519 37884 3528
rect 37832 3485 37841 3519
rect 37841 3485 37875 3519
rect 37875 3485 37884 3519
rect 37832 3476 37884 3485
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39948 3476 40000 3528
rect 40316 3519 40368 3528
rect 40316 3485 40325 3519
rect 40325 3485 40359 3519
rect 40359 3485 40368 3519
rect 40316 3476 40368 3485
rect 40408 3476 40460 3528
rect 41328 3519 41380 3528
rect 41328 3485 41337 3519
rect 41337 3485 41371 3519
rect 41371 3485 41380 3519
rect 41328 3476 41380 3485
rect 41512 3519 41564 3528
rect 41512 3485 41521 3519
rect 41521 3485 41555 3519
rect 41555 3485 41564 3519
rect 41512 3476 41564 3485
rect 45652 3519 45704 3528
rect 45652 3485 45661 3519
rect 45661 3485 45695 3519
rect 45695 3485 45704 3519
rect 45652 3476 45704 3485
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 16672 3340 16724 3392
rect 17316 3340 17368 3392
rect 19340 3340 19392 3392
rect 21272 3340 21324 3392
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 28632 3408 28684 3460
rect 36176 3451 36228 3460
rect 36176 3417 36185 3451
rect 36185 3417 36219 3451
rect 36219 3417 36228 3451
rect 36176 3408 36228 3417
rect 36452 3408 36504 3460
rect 30932 3340 30984 3392
rect 31392 3340 31444 3392
rect 36544 3340 36596 3392
rect 37740 3340 37792 3392
rect 48044 3408 48096 3460
rect 48964 3408 49016 3460
rect 42432 3340 42484 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3884 3136 3936 3188
rect 7288 3136 7340 3188
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 16856 3136 16908 3188
rect 19248 3136 19300 3188
rect 20904 3136 20956 3188
rect 21088 3136 21140 3188
rect 30196 3136 30248 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 9496 3068 9548 3120
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 16396 3068 16448 3120
rect 21180 3068 21232 3120
rect 22284 3111 22336 3120
rect 22284 3077 22293 3111
rect 22293 3077 22327 3111
rect 22327 3077 22336 3111
rect 22284 3068 22336 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 5816 3000 5868 3052
rect 7104 3000 7156 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 20076 3000 20128 3052
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 664 2932 716 2984
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 7748 2864 7800 2916
rect 10968 2932 11020 2984
rect 14188 2932 14240 2984
rect 17408 2932 17460 2984
rect 20168 2932 20220 2984
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 15108 2864 15160 2916
rect 26516 3068 26568 3120
rect 28908 3068 28960 3120
rect 24400 2975 24452 2984
rect 24400 2941 24409 2975
rect 24409 2941 24443 2975
rect 24443 2941 24452 2975
rect 24400 2932 24452 2941
rect 26148 2975 26200 2984
rect 26148 2941 26157 2975
rect 26157 2941 26191 2975
rect 26191 2941 26200 2975
rect 26148 2932 26200 2941
rect 36452 3136 36504 3188
rect 36544 3136 36596 3188
rect 46296 3136 46348 3188
rect 33232 3111 33284 3120
rect 33232 3077 33241 3111
rect 33241 3077 33275 3111
rect 33275 3077 33284 3111
rect 33232 3068 33284 3077
rect 39764 3068 39816 3120
rect 41604 3068 41656 3120
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 47768 3111 47820 3120
rect 47768 3077 47777 3111
rect 47777 3077 47811 3111
rect 47811 3077 47820 3111
rect 47768 3068 47820 3077
rect 33048 3043 33100 3052
rect 33048 3009 33057 3043
rect 33057 3009 33091 3043
rect 33091 3009 33100 3043
rect 33048 3000 33100 3009
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 41236 3000 41288 3052
rect 42432 3043 42484 3052
rect 30380 2975 30432 2984
rect 30380 2941 30389 2975
rect 30389 2941 30423 2975
rect 30423 2941 30432 2975
rect 33508 2975 33560 2984
rect 30380 2932 30432 2941
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 35992 2932 36044 2984
rect 35716 2864 35768 2916
rect 40316 2932 40368 2984
rect 41328 2975 41380 2984
rect 41328 2941 41337 2975
rect 41337 2941 41371 2975
rect 41371 2941 41380 2975
rect 41328 2932 41380 2941
rect 40408 2864 40460 2916
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 44272 2975 44324 2984
rect 44272 2941 44281 2975
rect 44281 2941 44315 2975
rect 44315 2941 44324 2975
rect 44272 2932 44324 2941
rect 46572 2932 46624 2984
rect 47676 2932 47728 2984
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18236 2796 18288 2848
rect 28264 2796 28316 2848
rect 30380 2796 30432 2848
rect 40592 2796 40644 2848
rect 42892 2796 42944 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 17316 2592 17368 2644
rect 17960 2592 18012 2644
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19984 2592 20036 2644
rect 20444 2635 20496 2644
rect 20444 2601 20453 2635
rect 20453 2601 20487 2635
rect 20487 2601 20496 2635
rect 20444 2592 20496 2601
rect 21824 2592 21876 2644
rect 24400 2592 24452 2644
rect 24492 2592 24544 2644
rect 8024 2524 8076 2576
rect 24584 2524 24636 2576
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 30656 2592 30708 2644
rect 35716 2635 35768 2644
rect 35716 2601 35725 2635
rect 35725 2601 35759 2635
rect 35759 2601 35768 2635
rect 35716 2592 35768 2601
rect 28356 2524 28408 2576
rect 28448 2524 28500 2576
rect 36176 2592 36228 2644
rect 39120 2592 39172 2644
rect 39304 2592 39356 2644
rect 42984 2635 43036 2644
rect 42984 2601 42993 2635
rect 42993 2601 43027 2635
rect 43027 2601 43036 2635
rect 42984 2592 43036 2601
rect 5172 2388 5224 2440
rect 15476 2388 15528 2440
rect 16120 2388 16172 2440
rect 16948 2388 17000 2440
rect 18052 2431 18104 2440
rect 18052 2397 18061 2431
rect 18061 2397 18095 2431
rect 18095 2397 18104 2431
rect 18052 2388 18104 2397
rect 19432 2388 19484 2440
rect 1308 2320 1360 2372
rect 2596 2320 2648 2372
rect 8392 2320 8444 2372
rect 29000 2456 29052 2508
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 32404 2456 32456 2508
rect 41512 2456 41564 2508
rect 43904 2499 43956 2508
rect 43904 2465 43913 2499
rect 43913 2465 43947 2499
rect 43947 2465 43956 2499
rect 43904 2456 43956 2465
rect 47032 2456 47084 2508
rect 23756 2388 23808 2440
rect 20628 2320 20680 2372
rect 23204 2320 23256 2372
rect 29644 2388 29696 2440
rect 36084 2388 36136 2440
rect 39856 2388 39908 2440
rect 41236 2388 41288 2440
rect 42892 2431 42944 2440
rect 42892 2397 42901 2431
rect 42901 2397 42935 2431
rect 42935 2397 42944 2431
rect 42892 2388 42944 2397
rect 43812 2388 43864 2440
rect 46020 2388 46072 2440
rect 24492 2320 24544 2372
rect 26424 2320 26476 2372
rect 27068 2320 27120 2372
rect 28356 2320 28408 2372
rect 35440 2320 35492 2372
rect 38016 2320 38068 2372
rect 39304 2320 39356 2372
rect 46388 2320 46440 2372
rect 48320 2320 48372 2372
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 15384 2252 15436 2304
rect 19156 2252 19208 2304
rect 21824 2252 21876 2304
rect 21916 2252 21968 2304
rect 25044 2252 25096 2304
rect 45468 2295 45520 2304
rect 45468 2261 45477 2295
rect 45477 2261 45511 2295
rect 45511 2261 45520 2295
rect 45468 2252 45520 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 17316 2048 17368 2100
rect 25504 2048 25556 2100
rect 3056 1980 3108 2032
rect 28080 1980 28132 2032
rect 20996 1912 21048 1964
rect 45468 1912 45520 1964
rect 21824 1844 21876 1896
rect 35992 1844 36044 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 19174 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 2608 47138 2636 49200
rect 2608 47110 2820 47138
rect 2792 47054 2820 47110
rect 3056 47116 3108 47122
rect 3056 47058 3108 47064
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2780 47048 2832 47054
rect 3068 47025 3096 47058
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 2780 46990 2832 46996
rect 3054 47016 3110 47025
rect 2320 46980 2372 46986
rect 3240 46990 3292 46996
rect 3054 46951 3110 46960
rect 2320 46922 2372 46928
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 1952 46368 2004 46374
rect 1952 46310 2004 46316
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 35698 1440 36110
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1504 35578 1532 43182
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1688 35894 1716 46310
rect 1964 45490 1992 46310
rect 1952 45484 2004 45490
rect 1952 45426 2004 45432
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 2044 40452 2096 40458
rect 2044 40394 2096 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 2056 36378 2084 40394
rect 2044 36372 2096 36378
rect 2044 36314 2096 36320
rect 2228 36100 2280 36106
rect 2228 36042 2280 36048
rect 1688 35866 1900 35894
rect 1504 35550 1808 35578
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1596 35086 1624 35391
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 34886
rect 1676 33448 1728 33454
rect 1676 33390 1728 33396
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1400 32836 1452 32842
rect 1400 32778 1452 32784
rect 1412 32026 1440 32778
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 1596 31822 1624 32671
rect 1688 32502 1716 33390
rect 1676 32496 1728 32502
rect 1676 32438 1728 32444
rect 1780 32314 1808 35550
rect 1688 32286 1808 32314
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1688 26234 1716 32286
rect 1768 31952 1820 31958
rect 1768 31894 1820 31900
rect 1596 26206 1716 26234
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23225 1440 23666
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1596 21350 1624 26206
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 20 19168 72 19174
rect 20 19110 72 19116
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 7478 1716 25162
rect 1780 23866 1808 31894
rect 1872 28762 1900 35866
rect 2240 35290 2268 36042
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2044 35216 2096 35222
rect 2044 35158 2096 35164
rect 1952 32360 2004 32366
rect 1952 32302 2004 32308
rect 1860 28756 1912 28762
rect 1860 28698 1912 28704
rect 1964 26234 1992 32302
rect 2056 31958 2084 35158
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2044 31952 2096 31958
rect 2044 31894 2096 31900
rect 2044 31816 2096 31822
rect 2044 31758 2096 31764
rect 2056 31346 2084 31758
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1964 26206 2084 26234
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18902 2084 26206
rect 2044 18896 2096 18902
rect 2044 18838 2096 18844
rect 2148 18766 2176 35022
rect 2332 23254 2360 46922
rect 3148 46912 3200 46918
rect 3148 46854 3200 46860
rect 3160 46646 3188 46854
rect 3148 46640 3200 46646
rect 3148 46582 3200 46588
rect 3896 46594 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 5828 47054 5856 49200
rect 7116 47054 7144 49200
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 3896 46566 4016 46594
rect 3988 46510 4016 46566
rect 3884 46504 3936 46510
rect 3884 46446 3936 46452
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2792 45422 2820 46271
rect 3896 46170 3924 46446
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 2872 45824 2924 45830
rect 2872 45766 2924 45772
rect 2884 45558 2912 45766
rect 2872 45552 2924 45558
rect 2872 45494 2924 45500
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 3330 44976 3386 44985
rect 3330 44911 3386 44920
rect 2412 41132 2464 41138
rect 2412 41074 2464 41080
rect 2320 23248 2372 23254
rect 2320 23190 2372 23196
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2424 18290 2452 41074
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36242 2820 36751
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 3344 35894 3372 44911
rect 3422 43616 3478 43625
rect 3422 43551 3478 43560
rect 3436 38842 3464 43551
rect 3514 39536 3570 39545
rect 3514 39471 3570 39480
rect 3528 39030 3556 39471
rect 3516 39024 3568 39030
rect 3516 38966 3568 38972
rect 3436 38814 3556 38842
rect 3344 35866 3464 35894
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2792 31278 2820 31991
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17202 1808 17614
rect 1964 17270 1992 18022
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 2976 17134 3004 31758
rect 3056 31680 3108 31686
rect 3056 31622 3108 31628
rect 3068 31414 3096 31622
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 3146 28656 3202 28665
rect 3146 28591 3202 28600
rect 3160 28490 3188 28591
rect 3148 28484 3200 28490
rect 3148 28426 3200 28432
rect 3436 23610 3464 35866
rect 3528 25770 3556 38814
rect 3792 32836 3844 32842
rect 3792 32778 3844 32784
rect 3804 32366 3832 32778
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 3698 31376 3754 31385
rect 3698 31311 3754 31320
rect 3516 25764 3568 25770
rect 3516 25706 3568 25712
rect 3436 23582 3556 23610
rect 3528 20602 3556 23582
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3436 19825 3464 20470
rect 3422 19816 3478 19825
rect 3422 19751 3478 19760
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 3068 18465 3096 19178
rect 3054 18456 3110 18465
rect 3054 18391 3110 18400
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2964 17128 3016 17134
rect 3068 17105 3096 17818
rect 3712 17746 3740 31311
rect 3804 19990 3832 32302
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 2964 17070 3016 17076
rect 3054 17096 3110 17105
rect 2792 16425 2820 17070
rect 3054 17031 3110 17040
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 2778 15056 2834 15065
rect 1768 15020 1820 15026
rect 2778 14991 2834 15000
rect 1768 14962 1820 14968
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 2148 3534 2176 14350
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13705 3464 13738
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 4080 12434 4108 46922
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3988 12406 4108 12434
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10305 3556 10950
rect 3514 10296 3570 10305
rect 3514 10231 3570 10240
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3160 3738 3188 4014
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1780 3058 1808 3470
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 1320 800 1348 2314
rect 2608 800 2636 2314
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 2038 3096 2246
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 3252 921 3280 4014
rect 3804 1465 3832 8774
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3896 3738 3924 3946
rect 3988 3942 4016 12406
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4816 11014 4844 20198
rect 5000 19961 5028 46922
rect 6920 46912 6972 46918
rect 6920 46854 6972 46860
rect 4986 19952 5042 19961
rect 4986 19887 5042 19896
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7585 4108 8230
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4066 6896 4122 6905
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6932 4690 6960 46854
rect 7564 39024 7616 39030
rect 7564 38966 7616 38972
rect 7576 27334 7604 38966
rect 7852 28422 7880 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9312 46912 9364 46918
rect 9312 46854 9364 46860
rect 8312 45526 8432 45554
rect 8312 29034 8340 45526
rect 9324 31890 9352 46854
rect 10980 46374 11008 49200
rect 11624 47054 11652 49200
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 11980 47048 12032 47054
rect 11980 46990 12032 46996
rect 11704 46504 11756 46510
rect 11704 46446 11756 46452
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 11716 46170 11744 46446
rect 11704 46164 11756 46170
rect 11704 46106 11756 46112
rect 11992 37194 12020 46990
rect 12268 46918 12296 49200
rect 12912 47054 12940 49200
rect 12900 47048 12952 47054
rect 13740 47036 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 13820 47048 13872 47054
rect 13740 47008 13820 47036
rect 12900 46990 12952 46996
rect 13820 46990 13872 46996
rect 12256 46912 12308 46918
rect 12256 46854 12308 46860
rect 14200 46510 14228 49200
rect 14648 46980 14700 46986
rect 14648 46922 14700 46928
rect 15384 46980 15436 46986
rect 15384 46922 15436 46928
rect 13820 46504 13872 46510
rect 13820 46446 13872 46452
rect 14004 46504 14056 46510
rect 14004 46446 14056 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 13832 46170 13860 46446
rect 13820 46164 13872 46170
rect 13820 46106 13872 46112
rect 14016 45626 14044 46446
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 45626 14136 45902
rect 14004 45620 14056 45626
rect 14004 45562 14056 45568
rect 14096 45620 14148 45626
rect 14096 45562 14148 45568
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 11980 37188 12032 37194
rect 11980 37130 12032 37136
rect 9312 31884 9364 31890
rect 9312 31826 9364 31832
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 12256 28008 12308 28014
rect 12256 27950 12308 27956
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12268 27674 12296 27950
rect 12544 27674 12572 27950
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8220 26926 8248 27270
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 8128 26586 8156 26862
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 7472 26240 7524 26246
rect 8036 26217 8064 26318
rect 7472 26182 7524 26188
rect 8022 26208 8078 26217
rect 7484 25974 7512 26182
rect 8022 26143 8078 26152
rect 7472 25968 7524 25974
rect 7472 25910 7524 25916
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8312 23322 8340 25774
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24818 8524 25230
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8496 23730 8524 24754
rect 9324 24614 9352 26794
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26450 9720 26726
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9416 25498 9444 26318
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 23798 9352 24550
rect 9876 24206 9904 25842
rect 10336 25294 10364 26794
rect 11164 26450 11192 26930
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10428 26042 10456 26250
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 11440 25294 11468 27406
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12360 26450 12388 27338
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12164 26376 12216 26382
rect 12360 26353 12388 26386
rect 12164 26318 12216 26324
rect 12346 26344 12402 26353
rect 11612 25832 11664 25838
rect 11612 25774 11664 25780
rect 11624 25498 11652 25774
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9876 23730 9904 24142
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8312 22710 8340 22918
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8404 22574 8432 23462
rect 9140 23118 9168 23598
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9600 22982 9628 23258
rect 9692 23186 9720 23666
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9600 22778 9628 22918
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8128 21010 8156 22034
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21418 9720 21830
rect 9784 21622 9812 23054
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9876 21554 9904 23666
rect 10060 23594 10088 25230
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10152 24750 10180 25094
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10244 24410 10272 24754
rect 10336 24682 10364 25230
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10048 23588 10100 23594
rect 10048 23530 10100 23536
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10152 22710 10180 23462
rect 10428 23322 10456 23462
rect 11900 23322 11928 25230
rect 12176 24682 12204 26318
rect 12346 26279 12402 26288
rect 12452 25838 12480 26726
rect 12544 26586 12572 26930
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12636 26217 12664 26726
rect 12622 26208 12678 26217
rect 12622 26143 12678 26152
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12072 23792 12124 23798
rect 12072 23734 12124 23740
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 10244 23066 10272 23258
rect 10600 23112 10652 23118
rect 10244 23038 10364 23066
rect 10600 23054 10652 23060
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10244 22438 10272 22918
rect 10336 22710 10364 23038
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10060 21894 10088 22374
rect 10336 21894 10364 22646
rect 10612 22506 10640 23054
rect 10968 23044 11020 23050
rect 10968 22986 11020 22992
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 10980 22778 11008 22986
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 11256 22098 11284 22986
rect 11808 22114 11836 22986
rect 12084 22438 12112 23734
rect 12452 22642 12480 24142
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12544 23662 12572 24006
rect 12820 23866 12848 24754
rect 12912 24206 12940 26998
rect 13280 26518 13308 27406
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13280 26382 13308 26454
rect 13372 26382 13400 27338
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 13268 26376 13320 26382
rect 13174 26344 13230 26353
rect 13268 26318 13320 26324
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13174 26279 13176 26288
rect 13228 26279 13230 26288
rect 13176 26250 13228 26256
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 13096 25498 13124 25842
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13268 24880 13320 24886
rect 13268 24822 13320 24828
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 13280 23730 13308 24822
rect 13372 24818 13400 26318
rect 13464 26246 13492 26386
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13464 25702 13492 26182
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13360 24132 13412 24138
rect 13360 24074 13412 24080
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 13280 23594 13308 23666
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13372 23050 13400 24074
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 12636 22642 12664 22986
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 11808 22098 11928 22114
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11808 22092 11940 22098
rect 11808 22086 11888 22092
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 7576 20466 7604 20878
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7944 20058 7972 20334
rect 8956 20058 8984 20878
rect 9876 20466 9904 21490
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 21146 9996 21286
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20534 9996 20810
rect 10060 20806 10088 21830
rect 10612 21078 10640 21966
rect 10876 21956 10928 21962
rect 10876 21898 10928 21904
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 10704 20466 10732 21286
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10888 20330 10916 21898
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8312 18970 8340 19382
rect 9140 19310 9168 19790
rect 8392 19304 8444 19310
rect 9128 19304 9180 19310
rect 8392 19246 8444 19252
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8128 18358 8156 18702
rect 8404 18630 8432 19246
rect 8496 19242 8708 19258
rect 9128 19246 9180 19252
rect 8484 19236 8720 19242
rect 8536 19230 8668 19236
rect 8484 19178 8536 19184
rect 8668 19178 8720 19184
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 9048 18426 9076 18702
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5816 3528 5868 3534
rect 4066 3496 4122 3505
rect 5816 3470 5868 3476
rect 4066 3431 4122 3440
rect 4080 3398 4108 3431
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3790 1456 3846 1465
rect 3790 1391 3846 1400
rect 3238 912 3294 921
rect 3238 847 3294 856
rect 3896 800 3924 3130
rect 5828 3058 5856 3470
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5184 800 5212 2382
rect 6472 800 6500 3538
rect 7116 3058 7144 4014
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2122 7236 3946
rect 8128 3534 8156 18294
rect 9140 18290 9168 19246
rect 11256 19174 11284 22034
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 21690 11376 21898
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11808 20466 11836 22086
rect 11888 22034 11940 22040
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11992 20262 12020 20878
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11992 19310 12020 20198
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 18426 9444 18634
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9784 18290 9812 19110
rect 11808 18834 11836 19110
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10244 18290 10272 18566
rect 10690 18456 10746 18465
rect 10796 18426 10824 18634
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10690 18391 10692 18400
rect 10744 18391 10746 18400
rect 10784 18420 10836 18426
rect 10692 18362 10744 18368
rect 10784 18362 10836 18368
rect 10782 18320 10838 18329
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 10232 18284 10284 18290
rect 10888 18290 10916 18566
rect 12084 18426 12112 22374
rect 12636 22094 12664 22578
rect 12452 22066 12664 22094
rect 12452 21554 12480 22066
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12452 19378 12480 21490
rect 12636 20466 12664 21830
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 20058 12848 20334
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 19174 12848 19314
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12438 18456 12494 18465
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 12072 18420 12124 18426
rect 12438 18391 12440 18400
rect 12072 18362 12124 18368
rect 12492 18391 12494 18400
rect 12440 18362 12492 18368
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 10782 18255 10784 18264
rect 10232 18226 10284 18232
rect 10836 18255 10838 18264
rect 10876 18284 10928 18290
rect 10784 18226 10836 18232
rect 10876 18226 10928 18232
rect 8588 18086 8616 18226
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 11348 17678 11376 18294
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11164 17270 11192 17614
rect 11532 17610 11560 18362
rect 12820 18329 12848 19110
rect 12806 18320 12862 18329
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11980 18284 12032 18290
rect 12806 18255 12862 18264
rect 11980 18226 12032 18232
rect 11716 17814 11744 18226
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11532 17082 11560 17546
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17270 11652 17478
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11992 17202 12020 18226
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11532 17054 11652 17082
rect 11624 16998 11652 17054
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11624 16574 11652 16934
rect 11992 16726 12020 17138
rect 12084 16794 12112 17546
rect 12636 17338 12664 18158
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12440 17196 12492 17202
rect 12176 17156 12440 17184
rect 12176 16998 12204 17156
rect 12440 17138 12492 17144
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 12360 16658 12388 16934
rect 12636 16658 12664 17274
rect 12820 17202 12848 18255
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 11624 16546 11836 16574
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15570 11100 15846
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11716 15026 11744 16050
rect 11808 15570 11836 16546
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 15366 12112 15506
rect 12360 15502 12388 15846
rect 12728 15706 12756 17138
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14482 11468 14758
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11716 14074 11744 14282
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11716 8498 11744 13806
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11808 7886 11836 9522
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9042 11928 9318
rect 12084 9110 12112 15302
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 12238 12296 14962
rect 12728 14822 12756 15642
rect 12912 15026 12940 22714
rect 13464 19378 13492 25638
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 23730 13584 25094
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 22778 13584 23666
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13648 22710 13676 22918
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13740 19922 13768 45426
rect 14660 34202 14688 46922
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 15396 29510 15424 46922
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 17420 47410 17448 49200
rect 16592 47382 17448 47410
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 15488 45526 16528 45554
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14200 27606 14228 28086
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 26382 13860 26930
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 13924 24954 13952 25774
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 14016 24834 14044 25230
rect 14108 25226 14136 27406
rect 14292 26518 14320 29038
rect 14476 28762 14504 29038
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 14660 28150 14688 28494
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14280 26512 14332 26518
rect 14280 26454 14332 26460
rect 14292 26042 14320 26454
rect 14464 26376 14516 26382
rect 14568 26353 14596 27950
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14660 26382 14688 27406
rect 15016 27396 15068 27402
rect 15016 27338 15068 27344
rect 15028 27130 15056 27338
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15028 26790 15056 26930
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 14648 26376 14700 26382
rect 14464 26318 14516 26324
rect 14554 26344 14610 26353
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 14200 25498 14228 25774
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 14292 25430 14320 25978
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14096 25220 14148 25226
rect 14096 25162 14148 25168
rect 13924 24806 14044 24834
rect 14384 24818 14412 26250
rect 14476 25498 14504 26318
rect 14648 26318 14700 26324
rect 14554 26279 14610 26288
rect 14568 26246 14596 26279
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14372 24812 14424 24818
rect 13924 24614 13952 24806
rect 14372 24754 14424 24760
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13832 23118 13860 23598
rect 13924 23186 13952 24550
rect 14384 23866 14412 24754
rect 14476 24614 14504 24754
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 14476 23118 14504 24550
rect 14844 23118 14872 25162
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 13832 21010 13860 23054
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22574 14320 22918
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 14476 22234 14504 23054
rect 14844 22438 14872 23054
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 14936 22710 14964 22918
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14844 21690 14872 22374
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14292 21010 14320 21286
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 15028 20534 15056 26726
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15304 25498 15332 25842
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15396 25294 15424 28494
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15580 28218 15608 28426
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 16500 27538 16528 45526
rect 16592 27946 16620 47382
rect 18708 47054 18736 49200
rect 19996 48226 20024 49200
rect 19996 48198 20116 48226
rect 19984 47252 20036 47258
rect 19984 47194 20036 47200
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 16960 32502 16988 46990
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19432 46504 19484 46510
rect 19432 46446 19484 46452
rect 19444 45490 19472 46446
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19432 45484 19484 45490
rect 19432 45426 19484 45432
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19168 33658 19196 35566
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 19904 35290 19932 35430
rect 19892 35284 19944 35290
rect 19892 35226 19944 35232
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19260 34406 19288 35022
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34610 20024 47194
rect 20088 47122 20116 48198
rect 20260 47184 20312 47190
rect 20260 47126 20312 47132
rect 20076 47116 20128 47122
rect 20076 47058 20128 47064
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 20180 46170 20208 46446
rect 20168 46164 20220 46170
rect 20168 46106 20220 46112
rect 20076 45960 20128 45966
rect 20076 45902 20128 45908
rect 20088 45422 20116 45902
rect 20076 45416 20128 45422
rect 20076 45358 20128 45364
rect 20088 35816 20116 45358
rect 20272 35873 20300 47126
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 20258 35864 20314 35873
rect 20088 35788 20208 35816
rect 20258 35799 20314 35808
rect 20074 35728 20130 35737
rect 20074 35663 20130 35672
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19248 34400 19300 34406
rect 19248 34342 19300 34348
rect 19260 33998 19288 34342
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19260 33538 19288 33934
rect 19432 33856 19484 33862
rect 19432 33798 19484 33804
rect 19444 33590 19472 33798
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 19168 33510 19288 33538
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 18524 32978 18552 33458
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 17224 32836 17276 32842
rect 17224 32778 17276 32784
rect 17236 32570 17264 32778
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 16948 32496 17000 32502
rect 16948 32438 17000 32444
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17788 31958 17816 32370
rect 17776 31952 17828 31958
rect 17776 31894 17828 31900
rect 17972 31482 18000 32914
rect 19168 32910 19196 33510
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32366 18092 32710
rect 18144 32496 18196 32502
rect 18144 32438 18196 32444
rect 18156 32366 18184 32438
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18144 32360 18196 32366
rect 18144 32302 18196 32308
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17868 30184 17920 30190
rect 17920 30132 18000 30138
rect 17868 30126 18000 30132
rect 17880 30110 18000 30126
rect 17972 29306 18000 30110
rect 18340 29714 18368 32370
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18616 30938 18644 31350
rect 19168 31346 19196 32846
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19340 32292 19392 32298
rect 19340 32234 19392 32240
rect 19156 31340 19208 31346
rect 19156 31282 19208 31288
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 19076 30802 19104 31078
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 19168 30734 19196 31282
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 19260 30938 19288 31214
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19352 30870 19380 32234
rect 19996 31822 20024 34546
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 19156 30728 19208 30734
rect 19156 30670 19208 30676
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 18340 29594 18368 29650
rect 18248 29566 18368 29594
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17328 28762 17356 29038
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 18248 28558 18276 29566
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 18328 29232 18380 29238
rect 18328 29174 18380 29180
rect 17684 28552 17736 28558
rect 17684 28494 17736 28500
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 17696 28014 17724 28494
rect 17880 28370 17908 28494
rect 18144 28484 18196 28490
rect 18144 28426 18196 28432
rect 18156 28370 18184 28426
rect 17880 28342 18184 28370
rect 18144 28144 18196 28150
rect 18144 28086 18196 28092
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 16580 27940 16632 27946
rect 16580 27882 16632 27888
rect 16868 27674 16896 27950
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16488 27532 16540 27538
rect 16488 27474 16540 27480
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16132 25498 16160 25842
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 15396 24818 15424 25230
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 15856 24954 15884 25094
rect 16316 24954 16344 25094
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15304 23798 15332 24346
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15120 22778 15148 23598
rect 15212 23594 15240 23666
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15304 23118 15332 23734
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15488 23050 15516 23666
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15212 22098 15240 22374
rect 15200 22092 15252 22098
rect 15488 22094 15516 22986
rect 15568 22094 15620 22098
rect 15200 22034 15252 22040
rect 15396 22092 15620 22094
rect 15396 22066 15568 22092
rect 15396 21622 15424 22066
rect 15568 22034 15620 22040
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15488 21486 15516 21898
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13188 18766 13216 19110
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18222 13124 18566
rect 13372 18408 13400 19110
rect 13280 18380 13400 18408
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13280 18086 13308 18380
rect 13556 18290 13584 19246
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13188 17338 13216 17614
rect 13372 17542 13400 18022
rect 13740 17882 13768 19246
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18290 14320 18566
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 16114 13216 17138
rect 13556 16726 13584 17478
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13188 15026 13216 16050
rect 14016 15910 14044 17138
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12728 14006 12756 14758
rect 13280 14346 13308 14758
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 13188 13938 13216 14214
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 12452 13462 12480 13874
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 13924 13258 13952 13670
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 12782 12664 13126
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11762 12296 12174
rect 12636 11762 12664 12718
rect 12820 12442 12848 12718
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 12268 10674 12296 11494
rect 12912 11218 12940 11494
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10742 12480 10950
rect 13832 10742 13860 11494
rect 13924 11150 13952 13194
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 13924 10470 13952 11086
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13832 9586 13860 9998
rect 14016 9654 14044 15846
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14200 12442 14228 12786
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11762 14136 12174
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 8090 11928 8366
rect 13556 8294 13584 8842
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3738 8248 4014
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7300 3194 7328 3334
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7116 2094 7236 2122
rect 7116 800 7144 2094
rect 7760 800 7788 2858
rect 8036 2582 8064 2926
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 3606
rect 9416 3602 9444 4558
rect 10428 4146 10456 7822
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11532 4146 11560 4218
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9508 3126 9536 3878
rect 9600 3602 9628 3878
rect 10060 3738 10088 3946
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 11532 3058 11560 3470
rect 11716 3126 11744 3878
rect 13648 3466 13676 9386
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 8566 13768 9318
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13832 7886 13860 9522
rect 14108 8498 14136 10406
rect 14292 9042 14320 14282
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 14384 6186 14412 20334
rect 15028 19854 15056 20470
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15212 18834 15240 19450
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17882 14504 18158
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 17202 14596 17614
rect 14660 17202 14688 18566
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15120 17202 15148 17546
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14568 16658 14596 16934
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14660 16114 14688 17138
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14568 13530 14596 13942
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14568 12646 14596 13466
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14660 10742 14688 16050
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 12238 14872 15302
rect 15212 15178 15240 15438
rect 15120 15150 15240 15178
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14936 14550 14964 14826
rect 15120 14822 15148 15150
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14936 14346 14964 14486
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 15120 14278 15148 14758
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15212 14074 15240 14962
rect 15304 14346 15332 15030
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15396 13190 15424 14214
rect 15488 13802 15516 20946
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15672 18222 15700 18634
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 12850 15424 13126
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11218 14964 12038
rect 15028 11694 15056 12582
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 15028 10130 15056 11630
rect 15212 11218 15240 12582
rect 15304 11626 15332 12786
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11762 15424 12174
rect 15488 11830 15516 13194
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14924 10056 14976 10062
rect 15120 10010 15148 10474
rect 14976 10004 15148 10010
rect 14924 9998 15148 10004
rect 14936 9982 15148 9998
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9654 14504 9862
rect 15120 9654 15148 9982
rect 15396 9722 15424 11698
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8090 14504 8842
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 13832 3058 13860 3470
rect 14016 3126 14044 3878
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 10980 800 11008 2926
rect 14200 800 14228 2926
rect 14844 800 14872 8366
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15120 2922 15148 3606
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15396 2310 15424 3538
rect 15580 2514 15608 4490
rect 15672 4078 15700 18158
rect 15764 15502 15792 23530
rect 15856 23322 15884 24142
rect 16316 24070 16344 24890
rect 16408 24750 16436 25230
rect 16868 24954 16896 25230
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16408 24206 16436 24686
rect 16684 24614 16712 24754
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23866 16344 24006
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16684 23730 16712 24550
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16776 23866 16804 24142
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15948 23118 15976 23462
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 21418 15976 23054
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 16132 18358 16160 22986
rect 16684 22642 16712 23666
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16500 21010 16528 22034
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16776 21690 16804 21898
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16316 18873 16344 18906
rect 16302 18864 16358 18873
rect 16302 18799 16358 18808
rect 16408 18426 16436 19858
rect 16592 19122 16620 20334
rect 16960 20262 16988 27406
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17972 25906 18000 26726
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 17144 25362 17172 25638
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 17972 23254 18000 25842
rect 18156 25362 18184 28086
rect 18340 27606 18368 29174
rect 18984 29034 19012 29242
rect 18972 29028 19024 29034
rect 18972 28970 19024 28976
rect 18788 28960 18840 28966
rect 18788 28902 18840 28908
rect 18800 28626 18828 28902
rect 18788 28620 18840 28626
rect 18788 28562 18840 28568
rect 18984 28082 19012 28970
rect 19352 28490 19380 30806
rect 19444 30326 19472 31078
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19982 30152 20038 30161
rect 19982 30087 20038 30096
rect 19996 29714 20024 30087
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19904 28558 19932 29106
rect 19984 28688 20036 28694
rect 19982 28656 19984 28665
rect 20036 28656 20038 28665
rect 19982 28591 20038 28600
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 19352 27606 19380 28086
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 26586 19472 27406
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 26580 19484 26586
rect 19432 26522 19484 26528
rect 19444 25922 19472 26522
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19444 25894 19564 25922
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19156 25424 19208 25430
rect 19156 25366 19208 25372
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 17960 23248 18012 23254
rect 17960 23190 18012 23196
rect 17972 22098 18000 23190
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17972 21554 18000 21830
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18156 21486 18184 25298
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18432 24818 18460 25162
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18248 23730 18276 24754
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18524 24410 18552 24686
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18340 23866 18368 24074
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21010 17080 21286
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17040 20392 17092 20398
rect 17038 20360 17040 20369
rect 17092 20360 17094 20369
rect 17038 20295 17094 20304
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16684 19378 16712 20198
rect 17420 19854 17448 20402
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19718 17448 19790
rect 18156 19718 18184 21422
rect 18248 20466 18276 21830
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18248 19786 18276 19926
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16500 19094 16712 19122
rect 16500 18834 16528 19094
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16592 18766 16620 18906
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16408 17814 16436 18362
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 16726 15976 17070
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 16408 15910 16436 17478
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14414 16068 14758
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16132 14346 16160 14486
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 15856 13530 15884 14282
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15764 12238 15792 13466
rect 16132 13258 16160 14282
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15856 11762 15884 12242
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 16408 3126 16436 15846
rect 16592 14890 16620 16050
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16684 14770 16712 19094
rect 17420 18290 17448 19654
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17604 18426 17632 19246
rect 18248 19174 18276 19722
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18340 18902 18368 21490
rect 18524 21418 18552 22578
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18708 22030 18736 22374
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18328 18896 18380 18902
rect 18420 18896 18472 18902
rect 18328 18838 18380 18844
rect 18418 18864 18420 18873
rect 18472 18864 18474 18873
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18426 18184 18566
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18340 18358 18368 18838
rect 18418 18799 18474 18808
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 16590 16804 18022
rect 17788 17678 17816 18226
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 17202 16896 17478
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 17788 16794 17816 17614
rect 18524 17134 18552 19382
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16776 15978 16804 16526
rect 16960 16250 16988 16526
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16960 16114 16988 16186
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16776 15434 16804 15914
rect 16960 15570 16988 16050
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15570 17172 15982
rect 17604 15706 17632 16390
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16960 15094 16988 15506
rect 17788 15502 17816 16730
rect 18340 16250 18368 17070
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18432 15910 18460 16186
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16592 14742 16712 14770
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 12306 16528 14214
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16592 11914 16620 14742
rect 16960 14498 16988 15030
rect 17052 15026 17080 15370
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 14550 17080 14962
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17144 14618 17172 14894
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16868 14470 16988 14498
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16868 14414 16896 14470
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 17144 14074 17172 14554
rect 17236 14550 17264 14758
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17328 13530 17356 13806
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17788 13326 17816 15438
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17972 15094 18000 15302
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 18064 15026 18092 15302
rect 18524 15162 18552 17070
rect 18616 16590 18644 17206
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 17880 14006 17908 14214
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 18432 13326 18460 14214
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18616 13530 18644 13942
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12306 16712 13126
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 16592 11886 16712 11914
rect 18064 11898 18092 12106
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16592 11218 16620 11766
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16592 9042 16620 11154
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16684 4214 16712 11886
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18432 11762 18460 13262
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 11150 16804 11494
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16776 9654 16804 9930
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16776 8090 16804 8842
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 17972 6866 18000 8978
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4622 17632 4966
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 17052 4146 17080 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16396 3120 16448 3126
rect 16396 3062 16448 3068
rect 16684 3058 16712 3334
rect 16776 3194 16804 3470
rect 16868 3194 16896 4082
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 16960 2446 16988 3878
rect 17236 3738 17264 3946
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17696 3534 17724 3878
rect 17788 3738 17816 4082
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3058 17356 3334
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15488 800 15516 2382
rect 16132 800 16160 2382
rect 17328 2106 17356 2586
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 17420 800 17448 2926
rect 17972 2650 18000 2994
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18064 2446 18092 2790
rect 18156 2650 18184 5170
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18248 2854 18276 4218
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18340 3534 18368 3878
rect 18432 3534 18460 3878
rect 18524 3738 18552 4082
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18708 800 18736 20810
rect 18984 18698 19012 23462
rect 19168 19446 19196 25366
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 24750 19380 25094
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19444 24274 19472 25774
rect 19536 25294 19564 25894
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23730 20024 25230
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19444 23322 19472 23598
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19260 22982 19288 23054
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19260 19394 19288 22918
rect 19444 22642 19472 23258
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19996 21962 20024 22374
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19616 21480 19668 21486
rect 19444 21428 19616 21434
rect 19444 21422 19668 21428
rect 19444 21406 19656 21422
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20534 19380 20742
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19444 19990 19472 21406
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20466 20024 20878
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19720 19922 19748 20198
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19446 19472 19654
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 19440 19484 19446
rect 19260 19378 19380 19394
rect 19432 19382 19484 19388
rect 19260 19372 19392 19378
rect 19260 19366 19340 19372
rect 19340 19314 19392 19320
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 19076 16658 19104 16934
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19076 16114 19104 16594
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 19076 3058 19104 3878
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19168 2310 19196 18838
rect 20088 18834 20116 35663
rect 20180 21486 20208 35788
rect 20260 35760 20312 35766
rect 20260 35702 20312 35708
rect 20272 35290 20300 35702
rect 20260 35284 20312 35290
rect 20260 35226 20312 35232
rect 20364 34134 20392 46990
rect 20640 46510 20668 49200
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 20732 46034 20760 46310
rect 21284 46034 21312 49200
rect 24584 47048 24636 47054
rect 24584 46990 24636 46996
rect 22192 46980 22244 46986
rect 22192 46922 22244 46928
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20824 35630 20852 35974
rect 20812 35624 20864 35630
rect 20812 35566 20864 35572
rect 21364 35624 21416 35630
rect 21364 35566 21416 35572
rect 20352 34128 20404 34134
rect 20352 34070 20404 34076
rect 21088 34128 21140 34134
rect 21088 34070 21140 34076
rect 21100 33998 21128 34070
rect 20720 33992 20772 33998
rect 20904 33992 20956 33998
rect 20720 33934 20772 33940
rect 20902 33960 20904 33969
rect 21088 33992 21140 33998
rect 20956 33960 20958 33969
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20548 32910 20576 33254
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20364 32473 20392 32710
rect 20548 32570 20576 32846
rect 20732 32774 20760 33934
rect 21088 33934 21140 33940
rect 20902 33895 20958 33904
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 20916 33114 20944 33798
rect 21284 33454 21312 33798
rect 21272 33448 21324 33454
rect 21272 33390 21324 33396
rect 21376 33318 21404 35566
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 22006 33960 22062 33969
rect 21732 33584 21784 33590
rect 21928 33572 21956 33934
rect 22006 33895 22008 33904
rect 22060 33895 22062 33904
rect 22008 33866 22060 33872
rect 21784 33544 21956 33572
rect 21732 33526 21784 33532
rect 21180 33312 21232 33318
rect 21180 33254 21232 33260
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 20996 32836 21048 32842
rect 20996 32778 21048 32784
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20350 32464 20406 32473
rect 20350 32399 20406 32408
rect 20260 31816 20312 31822
rect 20260 31758 20312 31764
rect 20272 26382 20300 31758
rect 20548 30938 20576 32506
rect 20536 30932 20588 30938
rect 20536 30874 20588 30880
rect 20628 30864 20680 30870
rect 20628 30806 20680 30812
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20272 25498 20300 25910
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20180 21010 20208 21286
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20272 20806 20300 21490
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20272 19990 20300 20742
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19444 16794 19472 17070
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 20272 16590 20300 19110
rect 19248 16584 19300 16590
rect 20260 16584 20312 16590
rect 19248 16526 19300 16532
rect 20258 16552 20260 16561
rect 20312 16552 20314 16561
rect 19260 16114 19288 16526
rect 20258 16487 20314 16496
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15978 19288 16050
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 15094 19380 15846
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19996 15162 20024 15302
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20364 12434 20392 30670
rect 20640 30666 20668 30806
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20444 30592 20496 30598
rect 20444 30534 20496 30540
rect 20456 29306 20484 30534
rect 20640 30258 20668 30602
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20548 29782 20576 30194
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 20640 29646 20668 29990
rect 20732 29850 20760 32710
rect 20904 31476 20956 31482
rect 20904 31418 20956 31424
rect 20916 31346 20944 31418
rect 21008 31414 21036 32778
rect 20996 31408 21048 31414
rect 20996 31350 21048 31356
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 20904 30864 20956 30870
rect 20904 30806 20956 30812
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20548 29170 20576 29446
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20456 28626 20484 28698
rect 20548 28642 20576 28902
rect 20444 28620 20496 28626
rect 20444 28562 20496 28568
rect 20548 28614 20760 28642
rect 20548 27402 20576 28614
rect 20732 28558 20760 28614
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20640 28014 20668 28494
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20640 27538 20668 27950
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 24682 20484 26930
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20548 24138 20576 26318
rect 20640 24410 20668 26454
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21010 20484 21286
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20640 16726 20668 24346
rect 20824 23050 20852 30330
rect 20916 29102 20944 30806
rect 21100 30734 21128 31282
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 20996 30184 21048 30190
rect 21100 30161 21128 30194
rect 20996 30126 21048 30132
rect 21086 30152 21142 30161
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20916 27878 20944 28358
rect 20904 27872 20956 27878
rect 20904 27814 20956 27820
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20916 22642 20944 23054
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20916 21554 20944 22578
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20732 17678 20760 18226
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20640 14414 20668 16662
rect 20732 16590 20760 17206
rect 20824 17066 20852 18022
rect 20916 17610 20944 18022
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20364 12406 20484 12434
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20088 4826 20116 5170
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19892 4616 19944 4622
rect 19944 4564 20024 4570
rect 19892 4558 20024 4564
rect 19904 4542 20024 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19260 3194 19288 4014
rect 19352 3738 19380 4082
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19352 800 19380 3334
rect 19444 2446 19472 3878
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 2650 20024 4542
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 3058 20116 3470
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20180 2990 20208 3674
rect 20272 3602 20300 3878
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 20364 1714 20392 3538
rect 20456 2650 20484 12406
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4622 20760 4966
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 3058 20760 4422
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20824 3602 20852 4082
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20916 3194 20944 4626
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 19996 1686 20392 1714
rect 19996 800 20024 1686
rect 20640 800 20668 2314
rect 21008 1970 21036 30126
rect 21086 30087 21142 30096
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 21100 29102 21128 29582
rect 21088 29096 21140 29102
rect 21088 29038 21140 29044
rect 21100 28762 21128 29038
rect 21088 28756 21140 28762
rect 21088 28698 21140 28704
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21100 26994 21128 27406
rect 21192 27334 21220 33254
rect 21364 33040 21416 33046
rect 21548 33040 21600 33046
rect 21416 33000 21548 33028
rect 21364 32982 21416 32988
rect 21548 32982 21600 32988
rect 21548 32836 21600 32842
rect 21548 32778 21600 32784
rect 21560 32570 21588 32778
rect 21548 32564 21600 32570
rect 21548 32506 21600 32512
rect 21928 32026 21956 33544
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 21456 31952 21508 31958
rect 21454 31920 21456 31929
rect 21508 31920 21510 31929
rect 21454 31855 21510 31864
rect 22204 31754 22232 46922
rect 24596 46578 24624 46990
rect 24584 46572 24636 46578
rect 24584 46514 24636 46520
rect 25148 46510 25176 49200
rect 25412 47048 25464 47054
rect 25412 46990 25464 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25424 46034 25452 46990
rect 25792 46034 25820 49200
rect 26608 47116 26660 47122
rect 26608 47058 26660 47064
rect 25412 46028 25464 46034
rect 25412 45970 25464 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 24676 45960 24728 45966
rect 24676 45902 24728 45908
rect 24688 45558 24716 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25320 45824 25372 45830
rect 25320 45766 25372 45772
rect 24676 45552 24728 45558
rect 24676 45494 24728 45500
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22664 37466 22692 38286
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22848 37942 22876 38150
rect 22836 37936 22888 37942
rect 22836 37878 22888 37884
rect 23848 37936 23900 37942
rect 23848 37878 23900 37884
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23388 37392 23440 37398
rect 23388 37334 23440 37340
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22572 36242 22600 36858
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 23204 36236 23256 36242
rect 23204 36178 23256 36184
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22480 35630 22508 35974
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 22376 34196 22428 34202
rect 22376 34138 22428 34144
rect 22284 33652 22336 33658
rect 22284 33594 22336 33600
rect 22296 32570 22324 33594
rect 22388 33590 22416 34138
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22468 33312 22520 33318
rect 22468 33254 22520 33260
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 22282 32056 22338 32065
rect 22282 31991 22338 32000
rect 22296 31890 22324 31991
rect 22388 31958 22416 32506
rect 22376 31952 22428 31958
rect 22376 31894 22428 31900
rect 22284 31884 22336 31890
rect 22284 31826 22336 31832
rect 22100 31748 22152 31754
rect 22204 31726 22416 31754
rect 22100 31690 22152 31696
rect 22112 31634 22140 31690
rect 22112 31606 22324 31634
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21836 30802 21864 31078
rect 21824 30796 21876 30802
rect 21824 30738 21876 30744
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21376 30326 21404 30670
rect 21640 30592 21692 30598
rect 21640 30534 21692 30540
rect 21364 30320 21416 30326
rect 21364 30262 21416 30268
rect 21652 29238 21680 30534
rect 22204 30258 22232 31350
rect 22296 31346 22324 31606
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22284 30796 22336 30802
rect 22284 30738 22336 30744
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21652 27606 21680 29174
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 22020 28558 22048 28902
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 28218 21864 28358
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21916 27600 21968 27606
rect 21916 27542 21968 27548
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 21192 27062 21220 27270
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21836 26450 21864 26930
rect 21928 26790 21956 27542
rect 22296 27538 22324 30738
rect 22284 27532 22336 27538
rect 22284 27474 22336 27480
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 22020 26926 22048 27338
rect 22204 26976 22232 27406
rect 22296 27130 22324 27474
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22284 26988 22336 26994
rect 22204 26948 22284 26976
rect 22284 26930 22336 26936
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 22020 26586 22048 26862
rect 22008 26580 22060 26586
rect 22008 26522 22060 26528
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 21548 26308 21600 26314
rect 21548 26250 21600 26256
rect 21560 25702 21588 26250
rect 22020 26246 22048 26318
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 21548 25696 21600 25702
rect 21548 25638 21600 25644
rect 21560 25158 21588 25638
rect 22020 25362 22048 26182
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 21088 25152 21140 25158
rect 21088 25094 21140 25100
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21100 24138 21128 25094
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 21376 24070 21404 25094
rect 22020 24410 22048 25298
rect 22296 25294 22324 26386
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24954 22140 25162
rect 22100 24948 22152 24954
rect 22100 24890 22152 24896
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 24410 22324 24686
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 21088 23248 21140 23254
rect 21088 23190 21140 23196
rect 21100 22642 21128 23190
rect 22112 23066 22140 23258
rect 22284 23112 22336 23118
rect 22112 23060 22284 23066
rect 22112 23054 22336 23060
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22112 23038 22324 23054
rect 22020 22778 22048 22986
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22030 21312 22578
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21284 21486 21312 21966
rect 22020 21962 22048 22714
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 21690 21956 21830
rect 22020 21690 22048 21898
rect 22112 21876 22140 23038
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22204 22234 22232 22918
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22388 22094 22416 31726
rect 22480 27614 22508 33254
rect 22664 33114 22692 33798
rect 22744 33584 22796 33590
rect 22744 33526 22796 33532
rect 22652 33108 22704 33114
rect 22652 33050 22704 33056
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22664 32434 22692 32846
rect 22652 32428 22704 32434
rect 22652 32370 22704 32376
rect 22756 31482 22784 33526
rect 22836 33040 22888 33046
rect 22836 32982 22888 32988
rect 22848 31686 22876 32982
rect 23032 32910 23060 34342
rect 23124 33386 23152 35634
rect 23112 33380 23164 33386
rect 23112 33322 23164 33328
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23032 32774 23060 32846
rect 23020 32768 23072 32774
rect 23020 32710 23072 32716
rect 23032 31958 23060 32710
rect 23020 31952 23072 31958
rect 23020 31894 23072 31900
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 22836 31680 22888 31686
rect 22836 31622 22888 31628
rect 22560 31476 22612 31482
rect 22560 31418 22612 31424
rect 22744 31476 22796 31482
rect 22744 31418 22796 31424
rect 22572 30734 22600 31418
rect 23032 31414 23060 31758
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 23216 31260 23244 36178
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23308 35086 23336 35566
rect 23296 35080 23348 35086
rect 23296 35022 23348 35028
rect 23308 34678 23336 35022
rect 23296 34672 23348 34678
rect 23296 34614 23348 34620
rect 23400 34406 23428 37334
rect 23492 37194 23520 37402
rect 23860 37262 23888 37878
rect 24216 37664 24268 37670
rect 24216 37606 24268 37612
rect 24308 37664 24360 37670
rect 24308 37606 24360 37612
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23480 37188 23532 37194
rect 23480 37130 23532 37136
rect 24228 36718 24256 37606
rect 24320 37262 24348 37606
rect 24492 37324 24544 37330
rect 24492 37266 24544 37272
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 24216 36712 24268 36718
rect 24216 36654 24268 36660
rect 23940 35080 23992 35086
rect 23940 35022 23992 35028
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23388 34400 23440 34406
rect 23388 34342 23440 34348
rect 23296 34196 23348 34202
rect 23296 34138 23348 34144
rect 23308 33318 23336 34138
rect 23388 33992 23440 33998
rect 23492 33980 23520 34886
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23584 34134 23612 34342
rect 23572 34128 23624 34134
rect 23572 34070 23624 34076
rect 23440 33952 23520 33980
rect 23388 33934 23440 33940
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23584 32910 23612 33254
rect 23676 32978 23704 34614
rect 23848 34400 23900 34406
rect 23848 34342 23900 34348
rect 23860 33862 23888 34342
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23664 32972 23716 32978
rect 23664 32914 23716 32920
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23584 32434 23612 32846
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23846 32464 23902 32473
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23480 32360 23532 32366
rect 23480 32302 23532 32308
rect 23296 32292 23348 32298
rect 23296 32234 23348 32240
rect 23308 31906 23336 32234
rect 23388 32224 23440 32230
rect 23388 32166 23440 32172
rect 23400 32026 23428 32166
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23308 31878 23428 31906
rect 22848 31232 23244 31260
rect 22560 30728 22612 30734
rect 22560 30670 22612 30676
rect 22572 29170 22600 30670
rect 22848 30054 22876 31232
rect 23400 30802 23428 31878
rect 23492 31822 23520 32302
rect 23572 31952 23624 31958
rect 23570 31920 23572 31929
rect 23624 31920 23626 31929
rect 23570 31855 23626 31864
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23664 31748 23716 31754
rect 23664 31690 23716 31696
rect 23676 31482 23704 31690
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22664 29306 22692 29990
rect 22652 29300 22704 29306
rect 22652 29242 22704 29248
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22480 27586 22600 27614
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22480 26994 22508 27066
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22572 26450 22600 27586
rect 22664 27470 22692 28018
rect 22848 27962 22876 29990
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 22940 28150 22968 29106
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 22744 27940 22796 27946
rect 22848 27934 22968 27962
rect 22744 27882 22796 27888
rect 22756 27606 22784 27882
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 22744 27600 22796 27606
rect 22744 27542 22796 27548
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22572 24818 22600 26250
rect 22664 25498 22692 26318
rect 22744 26308 22796 26314
rect 22848 26296 22876 27814
rect 22796 26268 22876 26296
rect 22744 26250 22796 26256
rect 22652 25492 22704 25498
rect 22652 25434 22704 25440
rect 22756 25226 22784 26250
rect 22744 25220 22796 25226
rect 22744 25162 22796 25168
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22940 24750 22968 27934
rect 23032 26994 23060 30194
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29050 23244 30126
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23584 29170 23612 29650
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23216 29034 23336 29050
rect 23216 29028 23348 29034
rect 23216 29022 23296 29028
rect 23296 28970 23348 28976
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23308 27470 23336 28970
rect 23492 28626 23520 28970
rect 23570 28656 23626 28665
rect 23480 28620 23532 28626
rect 23570 28591 23626 28600
rect 23480 28562 23532 28568
rect 23584 28558 23612 28591
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23124 26586 23152 26862
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23112 26444 23164 26450
rect 23112 26386 23164 26392
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25906 23060 26182
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 23124 25770 23152 26386
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 23216 25430 23244 26522
rect 23204 25424 23256 25430
rect 23204 25366 23256 25372
rect 23308 24750 23336 27406
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25362 23428 25842
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 23492 24834 23520 28358
rect 23584 27062 23612 28358
rect 23676 27946 23704 31418
rect 23768 30598 23796 32438
rect 23846 32399 23848 32408
rect 23900 32399 23902 32408
rect 23848 32370 23900 32376
rect 23952 31482 23980 35022
rect 24228 34542 24256 36654
rect 24504 36378 24532 37266
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 24596 36378 24624 37198
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24584 36372 24636 36378
rect 24584 36314 24636 36320
rect 24216 34536 24268 34542
rect 24216 34478 24268 34484
rect 24032 34060 24084 34066
rect 24032 34002 24084 34008
rect 24044 33969 24072 34002
rect 24030 33960 24086 33969
rect 24030 33895 24086 33904
rect 24228 33658 24256 34478
rect 24492 33992 24544 33998
rect 24492 33934 24544 33940
rect 24308 33924 24360 33930
rect 24308 33866 24360 33872
rect 24216 33652 24268 33658
rect 24216 33594 24268 33600
rect 24320 33538 24348 33866
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24228 33510 24348 33538
rect 24136 32570 24164 33458
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 24124 32360 24176 32366
rect 24122 32328 24124 32337
rect 24176 32328 24178 32337
rect 24122 32263 24178 32272
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 24136 31226 24164 31962
rect 23952 31198 24164 31226
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23848 30592 23900 30598
rect 23848 30534 23900 30540
rect 23768 29238 23796 30534
rect 23860 30190 23888 30534
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23952 30138 23980 31198
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 24044 30326 24072 31078
rect 24032 30320 24084 30326
rect 24032 30262 24084 30268
rect 23952 30110 24072 30138
rect 23848 29776 23900 29782
rect 23848 29718 23900 29724
rect 23756 29232 23808 29238
rect 23756 29174 23808 29180
rect 23860 29034 23888 29718
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 23848 29028 23900 29034
rect 23848 28970 23900 28976
rect 23952 28082 23980 29106
rect 24044 28150 24072 30110
rect 24228 28422 24256 33510
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 24320 32842 24348 33390
rect 24400 32972 24452 32978
rect 24400 32914 24452 32920
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 24308 30864 24360 30870
rect 24308 30806 24360 30812
rect 24320 28626 24348 30806
rect 24412 29646 24440 32914
rect 24400 29640 24452 29646
rect 24400 29582 24452 29588
rect 24308 28620 24360 28626
rect 24308 28562 24360 28568
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24032 28144 24084 28150
rect 24032 28086 24084 28092
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23584 26042 23612 26998
rect 23768 26382 23796 28018
rect 23952 27130 23980 28018
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 23492 24806 23612 24834
rect 23584 24750 23612 24806
rect 22928 24744 22980 24750
rect 22928 24686 22980 24692
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22296 22066 22416 22094
rect 22560 22092 22612 22098
rect 22192 21888 22244 21894
rect 22112 21848 22192 21876
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21928 21570 21956 21626
rect 21928 21542 22048 21570
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 20874 21220 21286
rect 22020 21010 22048 21542
rect 22112 21486 22140 21848
rect 22192 21830 22244 21836
rect 22100 21480 22152 21486
rect 22100 21422 22152 21428
rect 22192 21412 22244 21418
rect 22192 21354 22244 21360
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 22020 19854 22048 20946
rect 22204 20874 22232 21354
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21284 17882 21312 18158
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21192 17338 21220 17478
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21100 16726 21128 17070
rect 21284 16998 21312 17478
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21192 16114 21220 16526
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15570 21128 15846
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21376 12434 21404 19722
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21836 18290 21864 19314
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21928 18834 21956 19110
rect 22296 18834 22324 22066
rect 22560 22034 22612 22040
rect 22572 21690 22600 22034
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22664 21894 22692 21966
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22560 21072 22612 21078
rect 22560 21014 22612 21020
rect 22572 20466 22600 21014
rect 22664 20942 22692 21830
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19990 22508 20198
rect 22468 19984 22520 19990
rect 22468 19926 22520 19932
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 19825 22692 19858
rect 22650 19816 22706 19825
rect 22650 19751 22706 19760
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22664 18902 22692 19110
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 22204 17610 22232 18634
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22204 16590 22232 17546
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22388 15570 22416 16594
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 15706 22692 16526
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 21284 12406 21404 12434
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21100 3194 21128 3402
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21192 3126 21220 3402
rect 21284 3398 21312 12406
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21376 4826 21404 5170
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21928 4622 21956 4966
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22756 4010 22784 24550
rect 23308 24274 23336 24686
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22710 22968 22918
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 22234 22876 22510
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 20466 22876 21286
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 23216 20466 23244 20742
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 22848 19938 22876 20402
rect 22848 19922 23060 19938
rect 22848 19916 23072 19922
rect 22848 19910 23020 19916
rect 22940 17678 22968 19910
rect 23020 19858 23072 19864
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23032 18902 23060 19450
rect 23124 19378 23152 19654
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17338 23152 17614
rect 23308 17542 23336 19722
rect 23400 19446 23428 19858
rect 23676 19854 23704 20878
rect 23664 19848 23716 19854
rect 24308 19848 24360 19854
rect 23664 19790 23716 19796
rect 23938 19816 23994 19825
rect 24308 19790 24360 19796
rect 23938 19751 23994 19760
rect 23952 19718 23980 19751
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23860 19446 23888 19654
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23848 19440 23900 19446
rect 23848 19382 23900 19388
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23308 17082 23336 17478
rect 23492 17270 23520 17546
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17270 23980 17478
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23216 17066 23336 17082
rect 23204 17060 23336 17066
rect 23256 17054 23336 17060
rect 23860 17082 23888 17138
rect 23860 17054 23980 17082
rect 23204 17002 23256 17008
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23308 16726 23336 16934
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23768 16658 23796 16934
rect 23952 16658 23980 17054
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 24320 16590 24348 19790
rect 22836 16584 22888 16590
rect 22834 16552 22836 16561
rect 24308 16584 24360 16590
rect 22888 16552 22890 16561
rect 22834 16487 22890 16496
rect 24306 16552 24308 16561
rect 24360 16552 24362 16561
rect 24306 16487 24362 16496
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 22848 16114 22876 16390
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22940 15570 22968 16390
rect 23584 16046 23612 16390
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 24412 6914 24440 25842
rect 24504 20890 24532 33934
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24596 32502 24624 33594
rect 24584 32496 24636 32502
rect 24584 32438 24636 32444
rect 24596 32230 24624 32438
rect 24584 32224 24636 32230
rect 24584 32166 24636 32172
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24596 30734 24624 31078
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24596 29102 24624 29582
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24596 28082 24624 29038
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24688 26908 24716 45494
rect 25332 45490 25360 45766
rect 25424 45626 25452 45834
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 25320 45484 25372 45490
rect 25320 45426 25372 45432
rect 25228 37324 25280 37330
rect 25228 37266 25280 37272
rect 25044 36100 25096 36106
rect 25044 36042 25096 36048
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24872 35154 24900 35634
rect 25056 35494 25084 36042
rect 25240 35834 25268 37266
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 25044 35488 25096 35494
rect 25044 35430 25096 35436
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24780 32570 24808 34886
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 24860 33924 24912 33930
rect 24860 33866 24912 33872
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24780 32026 24808 32506
rect 24872 32230 24900 33866
rect 24860 32224 24912 32230
rect 24964 32212 24992 34002
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 25056 32910 25084 33254
rect 25228 33040 25280 33046
rect 25228 32982 25280 32988
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25148 32366 25176 32914
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 24964 32184 25176 32212
rect 24860 32166 24912 32172
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24780 28558 24808 29650
rect 24872 29170 24900 32166
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24964 30190 24992 31282
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24780 26994 24808 28018
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24596 26880 24716 26908
rect 24596 21486 24624 26880
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24688 23866 24716 24754
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24504 20862 24624 20890
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24504 20534 24532 20742
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24504 16182 24532 16390
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24412 6886 24532 6914
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21180 3120 21232 3126
rect 21180 3062 21232 3068
rect 22112 3058 22140 3470
rect 22296 3126 22324 3878
rect 23032 3534 23060 4422
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23124 3534 23152 4082
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23676 3534 23704 3878
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21836 2310 21864 2586
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 20996 1964 21048 1970
rect 20996 1906 21048 1912
rect 21836 1902 21864 2246
rect 21824 1896 21876 1902
rect 21824 1838 21876 1844
rect 21928 800 21956 2246
rect 22572 800 22600 2926
rect 23768 2446 23796 3334
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24412 2650 24440 2926
rect 24504 2650 24532 6886
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 24596 2582 24624 20862
rect 24688 17746 24716 23666
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17338 24716 17682
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24688 16046 24716 16594
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24780 8362 24808 26930
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24964 24274 24992 25094
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 24964 22098 24992 22510
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 19786 24900 20878
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24872 19242 24900 19722
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 23216 800 23244 2314
rect 24504 800 24532 2314
rect 25056 2310 25084 30194
rect 25148 29782 25176 32184
rect 25240 31958 25268 32982
rect 25228 31952 25280 31958
rect 25228 31894 25280 31900
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25240 31346 25268 31758
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25136 29776 25188 29782
rect 25136 29718 25188 29724
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25148 21554 25176 21966
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25148 20262 25176 21490
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25240 20330 25268 20538
rect 25228 20324 25280 20330
rect 25228 20266 25280 20272
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 19990 25176 20198
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25240 16114 25268 18294
rect 25332 16250 25360 45426
rect 26620 38554 26648 47058
rect 26700 46980 26752 46986
rect 26700 46922 26752 46928
rect 26608 38548 26660 38554
rect 26608 38490 26660 38496
rect 26148 38208 26200 38214
rect 26148 38150 26200 38156
rect 26160 37942 26188 38150
rect 26148 37936 26200 37942
rect 26148 37878 26200 37884
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25516 36854 25544 37062
rect 25504 36848 25556 36854
rect 25504 36790 25556 36796
rect 25504 36576 25556 36582
rect 25504 36518 25556 36524
rect 25516 36174 25544 36518
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25412 35488 25464 35494
rect 25412 35430 25464 35436
rect 25424 29646 25452 35430
rect 25700 35222 25728 35634
rect 25780 35488 25832 35494
rect 25780 35430 25832 35436
rect 25688 35216 25740 35222
rect 25688 35158 25740 35164
rect 25792 35086 25820 35430
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25780 34672 25832 34678
rect 25780 34614 25832 34620
rect 25792 34202 25820 34614
rect 25884 34610 25912 37198
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 26160 36378 26188 36654
rect 26332 36576 26384 36582
rect 26332 36518 26384 36524
rect 26148 36372 26200 36378
rect 26148 36314 26200 36320
rect 26056 36304 26108 36310
rect 26344 36258 26372 36518
rect 26056 36246 26108 36252
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 25976 35737 26004 36110
rect 25962 35728 26018 35737
rect 25962 35663 26018 35672
rect 25964 35624 26016 35630
rect 25964 35566 26016 35572
rect 25976 35494 26004 35566
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25976 34746 26004 35430
rect 26068 35086 26096 36246
rect 26160 36242 26372 36258
rect 26148 36236 26372 36242
rect 26200 36230 26372 36236
rect 26148 36178 26200 36184
rect 26344 36174 26372 36230
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26056 35080 26108 35086
rect 26056 35022 26108 35028
rect 26160 34898 26188 35974
rect 26252 35834 26280 36042
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 26344 35086 26372 36110
rect 26608 36032 26660 36038
rect 26608 35974 26660 35980
rect 26620 35698 26648 35974
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26068 34870 26188 34898
rect 25964 34740 26016 34746
rect 25964 34682 26016 34688
rect 25872 34604 25924 34610
rect 25872 34546 25924 34552
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25596 33108 25648 33114
rect 25596 33050 25648 33056
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25516 32366 25544 32778
rect 25504 32360 25556 32366
rect 25504 32302 25556 32308
rect 25504 31272 25556 31278
rect 25504 31214 25556 31220
rect 25516 30122 25544 31214
rect 25504 30116 25556 30122
rect 25504 30058 25556 30064
rect 25412 29640 25464 29646
rect 25412 29582 25464 29588
rect 25424 29306 25452 29582
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 25424 28626 25452 29242
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25516 28762 25544 29106
rect 25608 29034 25636 33050
rect 25884 33046 25912 34546
rect 26068 33522 26096 34870
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 26160 33590 26188 34682
rect 26240 33992 26292 33998
rect 26240 33934 26292 33940
rect 26148 33584 26200 33590
rect 26148 33526 26200 33532
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 26068 33114 26096 33458
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 25872 33040 25924 33046
rect 25872 32982 25924 32988
rect 25884 32774 25912 32982
rect 26160 32978 26188 33526
rect 26148 32972 26200 32978
rect 26148 32914 26200 32920
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 25872 32768 25924 32774
rect 25872 32710 25924 32716
rect 26068 32434 26096 32846
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26160 32434 26188 32710
rect 26252 32570 26280 33934
rect 26332 33380 26384 33386
rect 26332 33322 26384 33328
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 25872 31952 25924 31958
rect 25872 31894 25924 31900
rect 25884 30326 25912 31894
rect 25964 30660 26016 30666
rect 25964 30602 26016 30608
rect 25872 30320 25924 30326
rect 25872 30262 25924 30268
rect 25688 29300 25740 29306
rect 25688 29242 25740 29248
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25700 28558 25728 29242
rect 25688 28552 25740 28558
rect 25688 28494 25740 28500
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 25792 25294 25820 25638
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25976 24682 26004 30602
rect 26068 26994 26096 32370
rect 26344 32337 26372 33322
rect 26330 32328 26386 32337
rect 26330 32263 26332 32272
rect 26384 32263 26386 32272
rect 26332 32234 26384 32240
rect 26344 32203 26372 32234
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 26252 30802 26280 31214
rect 26240 30796 26292 30802
rect 26240 30738 26292 30744
rect 26252 29850 26280 30738
rect 26344 30258 26372 31758
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26240 29844 26292 29850
rect 26240 29786 26292 29792
rect 26344 29646 26372 30194
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26344 29306 26372 29582
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 26608 28960 26660 28966
rect 26608 28902 26660 28908
rect 26240 28688 26292 28694
rect 26240 28630 26292 28636
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26252 25294 26280 28630
rect 26620 28558 26648 28902
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 26344 27402 26372 27814
rect 26436 27674 26464 28358
rect 26516 28076 26568 28082
rect 26516 28018 26568 28024
rect 26424 27668 26476 27674
rect 26424 27610 26476 27616
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26528 27334 26556 28018
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26528 27130 26556 27270
rect 26516 27124 26568 27130
rect 26516 27066 26568 27072
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26528 25974 26556 26454
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26252 24750 26280 25230
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25700 23866 25728 24074
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25504 22024 25556 22030
rect 25504 21966 25556 21972
rect 25516 20874 25544 21966
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 26252 21690 26280 21898
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 21010 25820 21286
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25424 20369 25452 20538
rect 25516 20398 25544 20810
rect 25504 20392 25556 20398
rect 25410 20360 25466 20369
rect 25504 20334 25556 20340
rect 25410 20295 25466 20304
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25792 19378 25820 19790
rect 26160 19514 26188 20198
rect 26516 19984 26568 19990
rect 26516 19926 26568 19932
rect 26528 19786 26556 19926
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25792 18766 25820 19314
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 17746 25636 18566
rect 25884 18426 25912 19314
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25332 15570 25360 15846
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25332 3602 25360 3878
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 25424 1850 25452 3538
rect 25516 2106 25544 17614
rect 25884 12434 25912 18362
rect 25976 18290 26004 18634
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25976 16114 26004 18226
rect 26252 18222 26280 18702
rect 26240 18216 26292 18222
rect 26240 18158 26292 18164
rect 26252 17746 26280 18158
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 16114 26096 16458
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 25792 12406 25912 12434
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25608 4146 25636 11698
rect 25792 4146 25820 12406
rect 25976 11762 26004 16050
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25884 3942 25912 9930
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 26160 2990 26188 17682
rect 26528 3126 26556 19722
rect 26712 15570 26740 46922
rect 26792 34944 26844 34950
rect 26792 34886 26844 34892
rect 26804 34542 26832 34886
rect 26792 34536 26844 34542
rect 26792 34478 26844 34484
rect 26804 33998 26832 34478
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26804 30734 26832 31078
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 26804 28694 26832 30670
rect 26792 28688 26844 28694
rect 26792 28630 26844 28636
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 26896 28014 26924 28494
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26884 28008 26936 28014
rect 26884 27950 26936 27956
rect 26896 27674 26924 27950
rect 26884 27668 26936 27674
rect 26884 27610 26936 27616
rect 26988 27062 27016 28018
rect 26976 27056 27028 27062
rect 26976 26998 27028 27004
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26804 25906 26832 26182
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26804 25226 26832 25842
rect 26988 25770 27016 26998
rect 26976 25764 27028 25770
rect 26976 25706 27028 25712
rect 26792 25220 26844 25226
rect 26792 25162 26844 25168
rect 26804 24410 26832 25162
rect 26792 24404 26844 24410
rect 26792 24346 26844 24352
rect 27080 22778 27108 49200
rect 28368 47054 28396 49200
rect 29368 47184 29420 47190
rect 29368 47126 29420 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28264 46912 28316 46918
rect 28264 46854 28316 46860
rect 28276 46578 28304 46854
rect 28264 46572 28316 46578
rect 28264 46514 28316 46520
rect 27528 38412 27580 38418
rect 27528 38354 27580 38360
rect 27436 38208 27488 38214
rect 27436 38150 27488 38156
rect 27252 37800 27304 37806
rect 27252 37742 27304 37748
rect 27264 37262 27292 37742
rect 27448 37466 27476 38150
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 27540 37398 27568 38354
rect 27988 37936 28040 37942
rect 27988 37878 28040 37884
rect 27528 37392 27580 37398
rect 27528 37334 27580 37340
rect 28000 37262 28028 37878
rect 28540 37664 28592 37670
rect 28540 37606 28592 37612
rect 27252 37256 27304 37262
rect 27252 37198 27304 37204
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 27264 35766 27292 37198
rect 27816 36106 27844 37198
rect 28552 36786 28580 37606
rect 28540 36780 28592 36786
rect 28540 36722 28592 36728
rect 28264 36644 28316 36650
rect 28264 36586 28316 36592
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 27804 36100 27856 36106
rect 27804 36042 27856 36048
rect 27712 35828 27764 35834
rect 27712 35770 27764 35776
rect 27160 35760 27212 35766
rect 27160 35702 27212 35708
rect 27252 35760 27304 35766
rect 27252 35702 27304 35708
rect 27172 35086 27200 35702
rect 27344 35624 27396 35630
rect 27344 35566 27396 35572
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 27264 34678 27292 35430
rect 27356 35086 27384 35566
rect 27724 35494 27752 35770
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 27620 35216 27672 35222
rect 27620 35158 27672 35164
rect 27344 35080 27396 35086
rect 27344 35022 27396 35028
rect 27252 34672 27304 34678
rect 27252 34614 27304 34620
rect 27632 34134 27660 35158
rect 27712 35012 27764 35018
rect 27712 34954 27764 34960
rect 27724 34610 27752 34954
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27620 34128 27672 34134
rect 27620 34070 27672 34076
rect 27632 33522 27660 34070
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27724 33454 27752 34546
rect 27816 34066 27844 36042
rect 28080 36032 28132 36038
rect 28080 35974 28132 35980
rect 27894 35728 27950 35737
rect 28092 35698 28120 35974
rect 27894 35663 27950 35672
rect 28080 35692 28132 35698
rect 27804 34060 27856 34066
rect 27804 34002 27856 34008
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27252 33040 27304 33046
rect 27252 32982 27304 32988
rect 27264 31346 27292 32982
rect 27724 31686 27752 33390
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27816 31482 27844 31690
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 27252 31340 27304 31346
rect 27528 31340 27580 31346
rect 27252 31282 27304 31288
rect 27448 31300 27528 31328
rect 27448 29170 27476 31300
rect 27528 31282 27580 31288
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27632 29646 27660 31282
rect 27908 30938 27936 35663
rect 28080 35634 28132 35640
rect 28184 34950 28212 36110
rect 28276 35698 28304 36586
rect 28264 35692 28316 35698
rect 28264 35634 28316 35640
rect 28172 34944 28224 34950
rect 28172 34886 28224 34892
rect 27988 33312 28040 33318
rect 27988 33254 28040 33260
rect 28000 32910 28028 33254
rect 28080 32972 28132 32978
rect 28080 32914 28132 32920
rect 27988 32904 28040 32910
rect 27988 32846 28040 32852
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 28000 31754 28028 32166
rect 27988 31748 28040 31754
rect 27988 31690 28040 31696
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27448 28626 27476 29106
rect 27436 28620 27488 28626
rect 27436 28562 27488 28568
rect 27160 28484 27212 28490
rect 27160 28426 27212 28432
rect 27172 25974 27200 28426
rect 27540 27946 27568 29106
rect 27632 29102 27660 29582
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27724 28082 27752 28494
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27632 27606 27660 28018
rect 27620 27600 27672 27606
rect 27620 27542 27672 27548
rect 27724 27554 27752 28018
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 27724 27526 27844 27554
rect 27816 27470 27844 27526
rect 27804 27464 27856 27470
rect 27804 27406 27856 27412
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27264 25362 27292 26318
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 27264 25226 27292 25298
rect 27252 25220 27304 25226
rect 27252 25162 27304 25168
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 27172 22574 27200 23054
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 27356 21622 27384 25842
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27632 24818 27660 25434
rect 27724 25158 27752 26386
rect 27816 25498 27844 27406
rect 27908 27402 27936 27814
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27804 25492 27856 25498
rect 27804 25434 27856 25440
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27632 24426 27660 24754
rect 27724 24750 27752 25094
rect 27712 24744 27764 24750
rect 27712 24686 27764 24692
rect 27632 24398 27844 24426
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 20466 26832 20810
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 26804 20262 26832 20402
rect 27264 20262 27292 20402
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27264 20074 27292 20198
rect 27080 20046 27292 20074
rect 27080 18834 27108 20046
rect 27158 19952 27214 19961
rect 27158 19887 27214 19896
rect 27172 19446 27200 19887
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 27172 18766 27200 19382
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 26988 17202 27016 18702
rect 27068 18284 27120 18290
rect 27264 18272 27292 19790
rect 27448 19446 27476 21626
rect 27540 21554 27568 21898
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27540 20874 27568 21490
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27448 18766 27476 19382
rect 27632 18850 27660 24210
rect 27816 24206 27844 24398
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27816 23882 27844 24142
rect 28000 24138 28028 24346
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 27816 23866 27936 23882
rect 27816 23860 27948 23866
rect 27816 23854 27896 23860
rect 27896 23802 27948 23808
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 28000 21894 28028 22034
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27724 19718 27752 20334
rect 28000 19922 28028 21830
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27540 18822 27660 18850
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27120 18244 27292 18272
rect 27068 18226 27120 18232
rect 27264 17338 27292 18244
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27448 17202 27476 18702
rect 27540 17762 27568 18822
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27632 17882 27660 18702
rect 27816 18306 27844 19722
rect 27896 19236 27948 19242
rect 27896 19178 27948 19184
rect 27724 18278 27844 18306
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27540 17734 27660 17762
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 27540 3602 27568 16594
rect 27632 12986 27660 17734
rect 27724 14482 27752 18278
rect 27908 18222 27936 19178
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27896 18216 27948 18222
rect 27896 18158 27948 18164
rect 27816 17882 27844 18158
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 28000 17678 28028 19858
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 26516 3120 26568 3126
rect 26516 3062 26568 3068
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 25504 2100 25556 2106
rect 25504 2042 25556 2048
rect 25148 1822 25452 1850
rect 25148 800 25176 1822
rect 26436 800 26464 2314
rect 27080 800 27108 2314
rect 28092 2038 28120 32914
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28184 32502 28212 32846
rect 28276 32570 28304 35634
rect 28356 35284 28408 35290
rect 28356 35226 28408 35232
rect 28368 34542 28396 35226
rect 28552 35154 28580 36722
rect 28816 36712 28868 36718
rect 28816 36654 28868 36660
rect 28724 36372 28776 36378
rect 28724 36314 28776 36320
rect 28630 35728 28686 35737
rect 28630 35663 28632 35672
rect 28684 35663 28686 35672
rect 28632 35634 28684 35640
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 28540 35148 28592 35154
rect 28540 35090 28592 35096
rect 28540 34944 28592 34950
rect 28540 34886 28592 34892
rect 28552 34678 28580 34886
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28356 34536 28408 34542
rect 28356 34478 28408 34484
rect 28368 33998 28396 34478
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 28368 33590 28396 33934
rect 28356 33584 28408 33590
rect 28356 33526 28408 33532
rect 28368 33318 28396 33526
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28460 33114 28488 34546
rect 28644 33658 28672 35430
rect 28632 33652 28684 33658
rect 28632 33594 28684 33600
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28644 32994 28672 33594
rect 28552 32966 28672 32994
rect 28552 32774 28580 32966
rect 28736 32858 28764 36314
rect 28828 35834 28856 36654
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 29288 35834 29316 36110
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 29276 35828 29328 35834
rect 29276 35770 29328 35776
rect 28816 33312 28868 33318
rect 28816 33254 28868 33260
rect 28828 32910 28856 33254
rect 28644 32830 28764 32858
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 28540 32768 28592 32774
rect 28540 32710 28592 32716
rect 28264 32564 28316 32570
rect 28264 32506 28316 32512
rect 28172 32496 28224 32502
rect 28644 32450 28672 32830
rect 29012 32502 29040 32846
rect 28172 32438 28224 32444
rect 28184 31414 28212 32438
rect 28460 32434 28672 32450
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 29000 32496 29052 32502
rect 29000 32438 29052 32444
rect 28448 32428 28672 32434
rect 28500 32422 28672 32428
rect 28448 32370 28500 32376
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28276 32230 28304 32302
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 28644 32026 28672 32422
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28632 32020 28684 32026
rect 28632 31962 28684 31968
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28172 31408 28224 31414
rect 28172 31350 28224 31356
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28172 29572 28224 29578
rect 28172 29514 28224 29520
rect 28184 29170 28212 29514
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28172 28484 28224 28490
rect 28172 28426 28224 28432
rect 28184 28218 28212 28426
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28172 18148 28224 18154
rect 28172 18090 28224 18096
rect 28184 16114 28212 18090
rect 28276 18086 28304 31282
rect 28460 31278 28488 31622
rect 28448 31272 28500 31278
rect 28448 31214 28500 31220
rect 28448 30932 28500 30938
rect 28448 30874 28500 30880
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28368 29850 28396 30194
rect 28356 29844 28408 29850
rect 28356 29786 28408 29792
rect 28460 28422 28488 30874
rect 28736 30734 28764 32370
rect 28828 31822 28856 32438
rect 28906 32056 28962 32065
rect 28906 31991 28962 32000
rect 28920 31958 28948 31991
rect 28908 31952 28960 31958
rect 28908 31894 28960 31900
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28540 30320 28592 30326
rect 28540 30262 28592 30268
rect 28552 30054 28580 30262
rect 28736 30258 28764 30670
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28448 28416 28500 28422
rect 28448 28358 28500 28364
rect 28460 25838 28488 28358
rect 28552 28082 28580 29106
rect 28724 29096 28776 29102
rect 28724 29038 28776 29044
rect 28736 28558 28764 29038
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28632 28144 28684 28150
rect 28632 28086 28684 28092
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 28552 27878 28580 28018
rect 28540 27872 28592 27878
rect 28540 27814 28592 27820
rect 28644 27470 28672 28086
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28828 26858 28856 31758
rect 29276 31408 29328 31414
rect 29276 31350 29328 31356
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 29196 30666 29224 31282
rect 29184 30660 29236 30666
rect 29184 30602 29236 30608
rect 29288 30598 29316 31350
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 28906 30152 28962 30161
rect 28906 30087 28962 30096
rect 28920 30054 28948 30087
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29104 28218 29132 28902
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 28920 27878 28948 27950
rect 28908 27872 28960 27878
rect 28908 27814 28960 27820
rect 28920 27402 28948 27814
rect 28908 27396 28960 27402
rect 28908 27338 28960 27344
rect 29000 27328 29052 27334
rect 29000 27270 29052 27276
rect 29012 27130 29040 27270
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 29184 26988 29236 26994
rect 29012 26946 29184 26974
rect 28816 26852 28868 26858
rect 28816 26794 28868 26800
rect 28908 25900 28960 25906
rect 28908 25842 28960 25848
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28632 25696 28684 25702
rect 28632 25638 28684 25644
rect 28644 25294 28672 25638
rect 28920 25498 28948 25842
rect 29012 25838 29040 26946
rect 29184 26930 29236 26936
rect 29092 26852 29144 26858
rect 29092 26794 29144 26800
rect 29184 26852 29236 26858
rect 29184 26794 29236 26800
rect 29000 25832 29052 25838
rect 29000 25774 29052 25780
rect 28908 25492 28960 25498
rect 28908 25434 28960 25440
rect 28448 25288 28500 25294
rect 28448 25230 28500 25236
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28460 24206 28488 25230
rect 28736 24410 28764 25230
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28920 24410 28948 24686
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29012 24449 29040 24550
rect 28998 24440 29054 24449
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28908 24404 28960 24410
rect 28998 24375 29054 24384
rect 28908 24346 28960 24352
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28920 23866 28948 24210
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 28368 18698 28396 19314
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28276 2854 28304 17818
rect 28264 2848 28316 2854
rect 28264 2790 28316 2796
rect 28368 2582 28396 18634
rect 28460 17882 28488 21422
rect 28736 21010 28764 23666
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 28724 21004 28776 21010
rect 28724 20946 28776 20952
rect 28632 20868 28684 20874
rect 28632 20810 28684 20816
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28552 19378 28580 19994
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28552 18766 28580 19314
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28448 17876 28500 17882
rect 28448 17818 28500 17824
rect 28644 16658 28672 20810
rect 28828 20534 28856 21830
rect 28920 21690 28948 21830
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28816 20528 28868 20534
rect 28816 20470 28868 20476
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 19310 28856 19790
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28816 19304 28868 19310
rect 28816 19246 28868 19252
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28448 16040 28500 16046
rect 28448 15982 28500 15988
rect 28460 2582 28488 15982
rect 28644 11694 28672 16594
rect 28632 11688 28684 11694
rect 28632 11630 28684 11636
rect 28644 3466 28672 11630
rect 28632 3460 28684 3466
rect 28632 3402 28684 3408
rect 28920 3126 28948 19654
rect 29000 18352 29052 18358
rect 29000 18294 29052 18300
rect 29012 17882 29040 18294
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29104 6914 29132 26794
rect 29196 24750 29224 26794
rect 29288 25362 29316 30534
rect 29276 25356 29328 25362
rect 29276 25298 29328 25304
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29196 23526 29224 24686
rect 29288 24070 29316 25298
rect 29276 24064 29328 24070
rect 29276 24006 29328 24012
rect 29184 23520 29236 23526
rect 29184 23462 29236 23468
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29288 21690 29316 22510
rect 29380 22098 29408 47126
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49314 40030 50000
rect 39500 49286 40030 49314
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 31024 47048 31076 47054
rect 31024 46990 31076 46996
rect 29828 36848 29880 36854
rect 29828 36790 29880 36796
rect 29840 36378 29868 36790
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 29828 36372 29880 36378
rect 29828 36314 29880 36320
rect 30300 35698 30328 36518
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 29920 35012 29972 35018
rect 29920 34954 29972 34960
rect 30932 35012 30984 35018
rect 30932 34954 30984 34960
rect 29932 34746 29960 34954
rect 30944 34746 30972 34954
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 30932 34740 30984 34746
rect 30932 34682 30984 34688
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 30472 34536 30524 34542
rect 30472 34478 30524 34484
rect 29840 33318 29868 34478
rect 29920 34400 29972 34406
rect 29920 34342 29972 34348
rect 29932 34134 29960 34342
rect 29920 34128 29972 34134
rect 29920 34070 29972 34076
rect 29828 33312 29880 33318
rect 29828 33254 29880 33260
rect 29840 33046 29868 33254
rect 29828 33040 29880 33046
rect 29828 32982 29880 32988
rect 30012 33040 30064 33046
rect 30012 32982 30064 32988
rect 30024 32910 30052 32982
rect 30484 32910 30512 34478
rect 30564 33108 30616 33114
rect 30564 33050 30616 33056
rect 30576 32910 30604 33050
rect 30656 32972 30708 32978
rect 30656 32914 30708 32920
rect 30012 32904 30064 32910
rect 30012 32846 30064 32852
rect 30472 32904 30524 32910
rect 30472 32846 30524 32852
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 29552 32836 29604 32842
rect 29552 32778 29604 32784
rect 29564 30326 29592 32778
rect 30380 32768 30432 32774
rect 30380 32710 30432 32716
rect 30392 32502 30420 32710
rect 30380 32496 30432 32502
rect 30380 32438 30432 32444
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 29840 31890 29868 32302
rect 30378 32192 30434 32201
rect 30378 32127 30434 32136
rect 30392 32026 30420 32127
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30286 31920 30342 31929
rect 29828 31884 29880 31890
rect 30286 31855 30342 31864
rect 29828 31826 29880 31832
rect 30300 31822 30328 31855
rect 30288 31816 30340 31822
rect 30288 31758 30340 31764
rect 30380 31748 30432 31754
rect 30380 31690 30432 31696
rect 30392 31210 30420 31690
rect 30380 31204 30432 31210
rect 30380 31146 30432 31152
rect 30484 30734 30512 32846
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 29552 30320 29604 30326
rect 29552 30262 29604 30268
rect 30288 30320 30340 30326
rect 30288 30262 30340 30268
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29645 29640 29697 29646
rect 29645 29582 29697 29588
rect 29656 29306 29684 29582
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29736 27872 29788 27878
rect 29736 27814 29788 27820
rect 29748 27538 29776 27814
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29460 27396 29512 27402
rect 29460 27338 29512 27344
rect 29472 26790 29500 27338
rect 29840 26926 29868 29106
rect 29932 27946 29960 30194
rect 30104 30184 30156 30190
rect 30104 30126 30156 30132
rect 30012 29776 30064 29782
rect 30012 29718 30064 29724
rect 30024 29238 30052 29718
rect 30012 29232 30064 29238
rect 30012 29174 30064 29180
rect 29920 27940 29972 27946
rect 29920 27882 29972 27888
rect 29932 27674 29960 27882
rect 29920 27668 29972 27674
rect 29920 27610 29972 27616
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 29460 25152 29512 25158
rect 29460 25094 29512 25100
rect 29472 24750 29500 25094
rect 29840 24954 29868 25230
rect 29828 24948 29880 24954
rect 29828 24890 29880 24896
rect 29460 24744 29512 24750
rect 29460 24686 29512 24692
rect 29918 24440 29974 24449
rect 29918 24375 29920 24384
rect 29972 24375 29974 24384
rect 29920 24346 29972 24352
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29564 23662 29592 24006
rect 30024 23730 30052 27066
rect 30116 25294 30144 30126
rect 30196 29504 30248 29510
rect 30196 29446 30248 29452
rect 30208 29238 30236 29446
rect 30196 29232 30248 29238
rect 30196 29174 30248 29180
rect 30300 28150 30328 30262
rect 30288 28144 30340 28150
rect 30288 28086 30340 28092
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 30208 26926 30236 27406
rect 30196 26920 30248 26926
rect 30196 26862 30248 26868
rect 30300 25430 30328 28086
rect 30564 28076 30616 28082
rect 30564 28018 30616 28024
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30392 27334 30420 27950
rect 30576 27402 30604 28018
rect 30564 27396 30616 27402
rect 30564 27338 30616 27344
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30288 25424 30340 25430
rect 30288 25366 30340 25372
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30116 24206 30144 25230
rect 30300 24274 30328 25366
rect 30576 25294 30604 26318
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30576 24818 30604 25094
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30288 24268 30340 24274
rect 30288 24210 30340 24216
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 29552 23656 29604 23662
rect 29552 23598 29604 23604
rect 30380 23044 30432 23050
rect 30380 22986 30432 22992
rect 29368 22092 29420 22098
rect 29368 22034 29420 22040
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29276 21684 29328 21690
rect 29276 21626 29328 21632
rect 29564 19174 29592 21966
rect 30196 21004 30248 21010
rect 30392 20992 30420 22986
rect 30472 21004 30524 21010
rect 30392 20964 30472 20992
rect 30196 20946 30248 20952
rect 30472 20946 30524 20952
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29736 19304 29788 19310
rect 29736 19246 29788 19252
rect 29552 19168 29604 19174
rect 29552 19110 29604 19116
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29564 17678 29592 18702
rect 29748 17882 29776 19246
rect 29840 18834 29868 19314
rect 30208 19310 30236 20946
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 30208 18222 30236 19246
rect 30300 18766 30328 19382
rect 30380 19236 30432 19242
rect 30380 19178 30432 19184
rect 30392 18766 30420 19178
rect 30484 18970 30512 20946
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 30380 18760 30432 18766
rect 30380 18702 30432 18708
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30392 18034 30420 18702
rect 30300 18006 30420 18034
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 30300 17814 30328 18006
rect 30288 17808 30340 17814
rect 30288 17750 30340 17756
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29564 15638 29592 16526
rect 30484 16114 30512 18906
rect 30472 16108 30524 16114
rect 30472 16050 30524 16056
rect 29552 15632 29604 15638
rect 29552 15574 29604 15580
rect 30484 12434 30512 16050
rect 29012 6886 29132 6914
rect 30392 12406 30512 12434
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28448 2576 28500 2582
rect 28448 2518 28500 2524
rect 29012 2514 29040 6886
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 30024 2514 30052 4014
rect 30392 3210 30420 12406
rect 30208 3194 30420 3210
rect 30196 3188 30420 3194
rect 30248 3182 30420 3188
rect 30196 3130 30248 3136
rect 30392 2990 30420 3182
rect 30380 2984 30432 2990
rect 30380 2926 30432 2932
rect 30392 2854 30420 2926
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30668 2650 30696 32914
rect 30748 31204 30800 31210
rect 30748 31146 30800 31152
rect 30760 29646 30788 31146
rect 30748 29640 30800 29646
rect 30748 29582 30800 29588
rect 31036 29578 31064 46990
rect 32232 46442 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 45626 32352 46446
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 33324 45824 33376 45830
rect 33324 45766 33376 45772
rect 32312 45620 32364 45626
rect 32312 45562 32364 45568
rect 32220 45484 32272 45490
rect 32220 45426 32272 45432
rect 32232 37874 32260 45426
rect 32220 37868 32272 37874
rect 32220 37810 32272 37816
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31208 35624 31260 35630
rect 31208 35566 31260 35572
rect 31220 35086 31248 35566
rect 31208 35080 31260 35086
rect 31208 35022 31260 35028
rect 31404 34678 31432 35634
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 31944 35488 31996 35494
rect 31944 35430 31996 35436
rect 31956 35154 31984 35430
rect 32140 35222 32168 35566
rect 32128 35216 32180 35222
rect 32128 35158 32180 35164
rect 31944 35148 31996 35154
rect 31944 35090 31996 35096
rect 32232 35034 32260 37810
rect 32864 35624 32916 35630
rect 32864 35566 32916 35572
rect 32876 35290 32904 35566
rect 33140 35488 33192 35494
rect 33140 35430 33192 35436
rect 32864 35284 32916 35290
rect 32864 35226 32916 35232
rect 32956 35216 33008 35222
rect 32956 35158 33008 35164
rect 32772 35148 32824 35154
rect 32772 35090 32824 35096
rect 32140 35006 32260 35034
rect 31392 34672 31444 34678
rect 31392 34614 31444 34620
rect 31760 33312 31812 33318
rect 31760 33254 31812 33260
rect 31576 33108 31628 33114
rect 31576 33050 31628 33056
rect 31392 32768 31444 32774
rect 31392 32710 31444 32716
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31220 31482 31248 32370
rect 31404 32366 31432 32710
rect 31588 32366 31616 33050
rect 31772 32978 31800 33254
rect 31760 32972 31812 32978
rect 31760 32914 31812 32920
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 31392 32360 31444 32366
rect 31392 32302 31444 32308
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 31588 31822 31616 32302
rect 31680 32026 31708 32846
rect 31852 32564 31904 32570
rect 31852 32506 31904 32512
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31576 31816 31628 31822
rect 31576 31758 31628 31764
rect 31208 31476 31260 31482
rect 31208 31418 31260 31424
rect 31864 31346 31892 32506
rect 32036 32292 32088 32298
rect 32036 32234 32088 32240
rect 32048 31822 32076 32234
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 31852 31340 31904 31346
rect 31852 31282 31904 31288
rect 31392 30660 31444 30666
rect 31392 30602 31444 30608
rect 31024 29572 31076 29578
rect 31024 29514 31076 29520
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31220 28762 31248 29106
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 30932 28552 30984 28558
rect 30932 28494 30984 28500
rect 30944 27606 30972 28494
rect 31404 28014 31432 30602
rect 32140 28506 32168 35006
rect 32784 33318 32812 35090
rect 32864 35080 32916 35086
rect 32864 35022 32916 35028
rect 32876 34746 32904 35022
rect 32864 34740 32916 34746
rect 32864 34682 32916 34688
rect 32968 34542 32996 35158
rect 33152 35018 33180 35430
rect 33140 35012 33192 35018
rect 33140 34954 33192 34960
rect 33152 34610 33180 34954
rect 33048 34604 33100 34610
rect 33048 34546 33100 34552
rect 33140 34604 33192 34610
rect 33140 34546 33192 34552
rect 32956 34536 33008 34542
rect 32956 34478 33008 34484
rect 32772 33312 32824 33318
rect 32772 33254 32824 33260
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32232 32366 32260 32846
rect 32588 32768 32640 32774
rect 32588 32710 32640 32716
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32220 32360 32272 32366
rect 32220 32302 32272 32308
rect 32416 32026 32444 32370
rect 32496 32224 32548 32230
rect 32494 32192 32496 32201
rect 32548 32192 32550 32201
rect 32494 32127 32550 32136
rect 32220 32020 32272 32026
rect 32220 31962 32272 31968
rect 32404 32020 32456 32026
rect 32404 31962 32456 31968
rect 32232 31906 32260 31962
rect 32402 31920 32458 31929
rect 32232 31878 32352 31906
rect 32324 30734 32352 31878
rect 32402 31855 32458 31864
rect 32416 31822 32444 31855
rect 32404 31816 32456 31822
rect 32404 31758 32456 31764
rect 32508 30802 32536 32127
rect 32600 31754 32628 32710
rect 32968 32586 32996 34478
rect 33060 33114 33088 34546
rect 33336 34474 33364 45766
rect 38028 45554 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38384 46640 38436 46646
rect 38384 46582 38436 46588
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38396 45966 38424 46582
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 38384 45960 38436 45966
rect 38384 45902 38436 45908
rect 37292 45526 38056 45554
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34532 35222 34560 35974
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 35348 35148 35400 35154
rect 35348 35090 35400 35096
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 34532 34678 34560 34886
rect 34520 34672 34572 34678
rect 34520 34614 34572 34620
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 33324 34468 33376 34474
rect 33324 34410 33376 34416
rect 33048 33108 33100 33114
rect 33048 33050 33100 33056
rect 33428 33046 33456 34546
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35360 34202 35388 35090
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 35808 35080 35860 35086
rect 35808 35022 35860 35028
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 34796 34060 34848 34066
rect 34796 34002 34848 34008
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34532 33522 34560 33934
rect 34520 33516 34572 33522
rect 34520 33458 34572 33464
rect 33416 33040 33468 33046
rect 33416 32982 33468 32988
rect 32692 32570 32996 32586
rect 32680 32564 32996 32570
rect 32732 32558 32996 32564
rect 32680 32506 32732 32512
rect 32968 32502 32996 32558
rect 32956 32496 33008 32502
rect 32956 32438 33008 32444
rect 33416 32360 33468 32366
rect 33416 32302 33468 32308
rect 33428 31958 33456 32302
rect 34336 32020 34388 32026
rect 34336 31962 34388 31968
rect 33416 31952 33468 31958
rect 32678 31920 32734 31929
rect 33416 31894 33468 31900
rect 33600 31952 33652 31958
rect 33600 31894 33652 31900
rect 32678 31855 32734 31864
rect 32588 31748 32640 31754
rect 32588 31690 32640 31696
rect 32496 30796 32548 30802
rect 32496 30738 32548 30744
rect 32600 30734 32628 31690
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32496 30660 32548 30666
rect 32496 30602 32548 30608
rect 32404 30592 32456 30598
rect 32404 30534 32456 30540
rect 32416 29170 32444 30534
rect 32508 29850 32536 30602
rect 32692 30410 32720 31855
rect 33612 31822 33640 31894
rect 34348 31822 34376 31962
rect 32864 31816 32916 31822
rect 32600 30382 32720 30410
rect 32784 31764 32864 31770
rect 32784 31758 32916 31764
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 34336 31816 34388 31822
rect 34336 31758 34388 31764
rect 34428 31816 34480 31822
rect 34428 31758 34480 31764
rect 32784 31742 32904 31758
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32404 29164 32456 29170
rect 32404 29106 32456 29112
rect 32508 29102 32536 29786
rect 32600 29170 32628 30382
rect 32784 30122 32812 31742
rect 32956 31680 33008 31686
rect 32956 31622 33008 31628
rect 32968 31414 32996 31622
rect 34348 31482 34376 31758
rect 34336 31476 34388 31482
rect 34336 31418 34388 31424
rect 32956 31408 33008 31414
rect 32956 31350 33008 31356
rect 33508 31408 33560 31414
rect 33508 31350 33560 31356
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33428 30734 33456 31214
rect 33520 30938 33548 31350
rect 33508 30932 33560 30938
rect 33508 30874 33560 30880
rect 33416 30728 33468 30734
rect 33416 30670 33468 30676
rect 33428 30258 33456 30670
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 32772 30116 32824 30122
rect 32772 30058 32824 30064
rect 32680 29572 32732 29578
rect 32680 29514 32732 29520
rect 32692 29238 32720 29514
rect 32680 29232 32732 29238
rect 32680 29174 32732 29180
rect 32784 29186 32812 30058
rect 33692 30048 33744 30054
rect 33692 29990 33744 29996
rect 33704 29578 33732 29990
rect 34440 29850 34468 31758
rect 34532 31754 34560 33458
rect 34612 33448 34664 33454
rect 34612 33390 34664 33396
rect 34624 31958 34652 33390
rect 34808 33386 34836 34002
rect 34796 33380 34848 33386
rect 34796 33322 34848 33328
rect 35348 33380 35400 33386
rect 35348 33322 35400 33328
rect 34808 32910 34836 33322
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34796 32904 34848 32910
rect 34796 32846 34848 32852
rect 35072 32768 35124 32774
rect 35072 32710 35124 32716
rect 35084 32502 35112 32710
rect 35072 32496 35124 32502
rect 35072 32438 35124 32444
rect 34704 32360 34756 32366
rect 34704 32302 34756 32308
rect 34612 31952 34664 31958
rect 34612 31894 34664 31900
rect 34716 31890 34744 32302
rect 34796 32292 34848 32298
rect 34796 32234 34848 32240
rect 34808 32026 34836 32234
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34796 32020 34848 32026
rect 34796 31962 34848 31968
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 34888 31884 34940 31890
rect 34888 31826 34940 31832
rect 34520 31748 34572 31754
rect 34520 31690 34572 31696
rect 34716 31482 34744 31826
rect 34796 31748 34848 31754
rect 34796 31690 34848 31696
rect 34704 31476 34756 31482
rect 34704 31418 34756 31424
rect 34808 31142 34836 31690
rect 34900 31346 34928 31826
rect 35360 31414 35388 33322
rect 35452 32910 35480 35022
rect 35532 35012 35584 35018
rect 35532 34954 35584 34960
rect 35544 34202 35572 34954
rect 35716 34944 35768 34950
rect 35716 34886 35768 34892
rect 35728 34678 35756 34886
rect 35716 34672 35768 34678
rect 35716 34614 35768 34620
rect 35716 34400 35768 34406
rect 35716 34342 35768 34348
rect 35532 34196 35584 34202
rect 35532 34138 35584 34144
rect 35728 34066 35756 34342
rect 35716 34060 35768 34066
rect 35716 34002 35768 34008
rect 35532 33312 35584 33318
rect 35532 33254 35584 33260
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 35544 31346 35572 33254
rect 35716 32972 35768 32978
rect 35716 32914 35768 32920
rect 35624 32836 35676 32842
rect 35624 32778 35676 32784
rect 35636 32026 35664 32778
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 35728 31482 35756 32914
rect 35820 32910 35848 35022
rect 36268 34740 36320 34746
rect 36268 34682 36320 34688
rect 36176 34060 36228 34066
rect 36176 34002 36228 34008
rect 35900 33992 35952 33998
rect 35900 33934 35952 33940
rect 35912 33114 35940 33934
rect 35900 33108 35952 33114
rect 35900 33050 35952 33056
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35808 32224 35860 32230
rect 35808 32166 35860 32172
rect 35820 31890 35848 32166
rect 35808 31884 35860 31890
rect 35808 31826 35860 31832
rect 35912 31686 35940 33050
rect 36084 32768 36136 32774
rect 36084 32710 36136 32716
rect 36096 32502 36124 32710
rect 36084 32496 36136 32502
rect 36084 32438 36136 32444
rect 35900 31680 35952 31686
rect 35900 31622 35952 31628
rect 35716 31476 35768 31482
rect 35716 31418 35768 31424
rect 34888 31340 34940 31346
rect 34888 31282 34940 31288
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 34796 31136 34848 31142
rect 34796 31078 34848 31084
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34428 29844 34480 29850
rect 34428 29786 34480 29792
rect 33692 29572 33744 29578
rect 33692 29514 33744 29520
rect 32784 29170 32904 29186
rect 32588 29164 32640 29170
rect 32784 29164 32916 29170
rect 32784 29158 32864 29164
rect 32588 29106 32640 29112
rect 32864 29106 32916 29112
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32772 29096 32824 29102
rect 32772 29038 32824 29044
rect 32140 28478 32628 28506
rect 32496 28416 32548 28422
rect 32496 28358 32548 28364
rect 32508 28082 32536 28358
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 31392 28008 31444 28014
rect 31392 27950 31444 27956
rect 32220 28008 32272 28014
rect 32220 27950 32272 27956
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 31036 27674 31064 27814
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 31392 27532 31444 27538
rect 31392 27474 31444 27480
rect 31116 27056 31168 27062
rect 31116 26998 31168 27004
rect 31128 26586 31156 26998
rect 31404 26994 31432 27474
rect 32232 27334 32260 27950
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32312 27396 32364 27402
rect 32312 27338 32364 27344
rect 32220 27328 32272 27334
rect 32220 27270 32272 27276
rect 32324 27062 32352 27338
rect 32312 27056 32364 27062
rect 32312 26998 32364 27004
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 31404 26382 31432 26930
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31404 19378 31432 21490
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 31208 19168 31260 19174
rect 31208 19110 31260 19116
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 31220 18766 31248 19110
rect 32128 18964 32180 18970
rect 32128 18906 32180 18912
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 32140 18290 32168 18906
rect 32324 18358 32352 19110
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 31484 18216 31536 18222
rect 31484 18158 31536 18164
rect 31496 4826 31524 18158
rect 32220 6180 32272 6186
rect 32220 6122 32272 6128
rect 31484 4820 31536 4826
rect 31484 4762 31536 4768
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30656 2644 30708 2650
rect 30656 2586 30708 2592
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28080 2032 28132 2038
rect 28080 1974 28132 1980
rect 28368 800 28396 2314
rect 29656 800 29684 2382
rect 30852 1986 30880 3878
rect 30944 3398 30972 4082
rect 31392 4072 31444 4078
rect 31392 4014 31444 4020
rect 31404 3398 31432 4014
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 30852 1958 30972 1986
rect 30944 800 30972 1958
rect 32232 800 32260 6122
rect 32416 2514 32444 27814
rect 32600 20806 32628 28478
rect 32588 20800 32640 20806
rect 32588 20742 32640 20748
rect 32784 5030 32812 29038
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 33784 20596 33836 20602
rect 33784 20538 33836 20544
rect 33796 20398 33824 20538
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 33508 19168 33560 19174
rect 33508 19110 33560 19116
rect 33520 18902 33548 19110
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 33508 18896 33560 18902
rect 33508 18838 33560 18844
rect 33968 18216 34020 18222
rect 33968 18158 34020 18164
rect 32772 5024 32824 5030
rect 32772 4966 32824 4972
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33060 3058 33088 3470
rect 33244 3126 33272 3878
rect 33980 3738 34008 18158
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 36188 4078 36216 34002
rect 36280 33998 36308 34682
rect 36268 33992 36320 33998
rect 36268 33934 36320 33940
rect 36280 31822 36308 33934
rect 36268 31816 36320 31822
rect 36268 31758 36320 31764
rect 37292 22030 37320 45526
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 38212 16182 38240 45902
rect 39500 45554 39528 49286
rect 39918 49200 40030 49286
rect 40562 49200 40674 50000
rect 41206 49314 41318 50000
rect 40788 49286 41318 49314
rect 40788 47410 40816 49286
rect 41206 49200 41318 49286
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 41892 47546 41920 49200
rect 41892 47518 42012 47546
rect 38672 45526 39528 45554
rect 40052 47382 40816 47410
rect 38568 21888 38620 21894
rect 38568 21830 38620 21836
rect 38580 21418 38608 21830
rect 38568 21412 38620 21418
rect 38568 21354 38620 21360
rect 38672 16590 38700 45526
rect 40052 22574 40080 47382
rect 41880 47048 41932 47054
rect 41880 46990 41932 46996
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40420 25362 40448 46922
rect 41892 46578 41920 46990
rect 41880 46572 41932 46578
rect 41880 46514 41932 46520
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41340 46034 41368 46310
rect 41984 46034 42012 47518
rect 42536 46442 42564 49200
rect 42616 47048 42668 47054
rect 42616 46990 42668 46996
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41972 46028 42024 46034
rect 41972 45970 42024 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45626 41552 45834
rect 41512 45620 41564 45626
rect 41512 45562 41564 45568
rect 40684 45552 40736 45558
rect 40684 45494 40736 45500
rect 40696 45014 40724 45494
rect 42628 45082 42656 46990
rect 42800 46980 42852 46986
rect 42800 46922 42852 46928
rect 42812 45558 42840 46922
rect 43180 46918 43208 49200
rect 43168 46912 43220 46918
rect 43168 46854 43220 46860
rect 43536 46368 43588 46374
rect 43536 46310 43588 46316
rect 42800 45552 42852 45558
rect 42800 45494 42852 45500
rect 42616 45076 42668 45082
rect 42616 45018 42668 45024
rect 40684 45008 40736 45014
rect 40684 44950 40736 44956
rect 43444 40928 43496 40934
rect 43444 40870 43496 40876
rect 40408 25356 40460 25362
rect 40408 25298 40460 25304
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 40040 22568 40092 22574
rect 40040 22510 40092 22516
rect 39580 21956 39632 21962
rect 39580 21898 39632 21904
rect 39592 21486 39620 21898
rect 42812 21622 42840 22918
rect 43456 22030 43484 40870
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 42800 21616 42852 21622
rect 42800 21558 42852 21564
rect 39304 21480 39356 21486
rect 39304 21422 39356 21428
rect 39580 21480 39632 21486
rect 39580 21422 39632 21428
rect 38660 16584 38712 16590
rect 38660 16526 38712 16532
rect 38200 16176 38252 16182
rect 38200 16118 38252 16124
rect 36176 4072 36228 4078
rect 36176 4014 36228 4020
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 37832 4004 37884 4010
rect 37832 3946 37884 3952
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 36556 3738 36584 3946
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 37844 3534 37872 3946
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37832 3528 37884 3534
rect 37832 3470 37884 3476
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 33232 3120 33284 3126
rect 33232 3062 33284 3068
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 36004 2990 36032 3470
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 36452 3460 36504 3466
rect 36452 3402 36504 3408
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 32404 2508 32456 2514
rect 32404 2450 32456 2456
rect 33520 800 33548 2926
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35728 2650 35756 2858
rect 35716 2644 35768 2650
rect 35716 2586 35768 2592
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 35452 800 35480 2314
rect 36004 1902 36032 2926
rect 36188 2650 36216 3402
rect 36464 3194 36492 3402
rect 36544 3392 36596 3398
rect 36544 3334 36596 3340
rect 37740 3392 37792 3398
rect 37740 3334 37792 3340
rect 36556 3194 36584 3334
rect 36452 3188 36504 3194
rect 36452 3130 36504 3136
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 37752 3058 37780 3334
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 39132 2650 39160 3470
rect 39316 2650 39344 21422
rect 40776 20324 40828 20330
rect 40776 20266 40828 20272
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40696 19786 40724 20198
rect 40684 19780 40736 19786
rect 40684 19722 40736 19728
rect 40788 19378 40816 20266
rect 40960 19780 41012 19786
rect 40960 19722 41012 19728
rect 42616 19780 42668 19786
rect 42616 19722 42668 19728
rect 40972 19514 41000 19722
rect 40960 19508 41012 19514
rect 40960 19450 41012 19456
rect 40776 19372 40828 19378
rect 40776 19314 40828 19320
rect 41328 4276 41380 4282
rect 41328 4218 41380 4224
rect 39764 4140 39816 4146
rect 39764 4082 39816 4088
rect 39776 3126 39804 4082
rect 39856 3936 39908 3942
rect 39856 3878 39908 3884
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 39304 2644 39356 2650
rect 39304 2586 39356 2592
rect 39868 2446 39896 3878
rect 41236 3732 41288 3738
rect 41236 3674 41288 3680
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 35992 1896 36044 1902
rect 35992 1838 36044 1844
rect 36096 800 36124 2382
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 38028 800 38056 2314
rect 39316 800 39344 2314
rect 39960 800 39988 3470
rect 40328 2990 40356 3470
rect 40316 2984 40368 2990
rect 40316 2926 40368 2932
rect 40420 2922 40448 3470
rect 41248 3058 41276 3674
rect 41340 3534 41368 4218
rect 42628 3738 42656 19722
rect 43444 19712 43496 19718
rect 43444 19654 43496 19660
rect 42984 19372 43036 19378
rect 42984 19314 43036 19320
rect 42708 8424 42760 8430
rect 42708 8366 42760 8372
rect 42720 4214 42748 8366
rect 42892 4616 42944 4622
rect 42892 4558 42944 4564
rect 42708 4208 42760 4214
rect 42708 4150 42760 4156
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42616 3732 42668 3738
rect 42616 3674 42668 3680
rect 42812 3602 42840 3878
rect 42904 3670 42932 4558
rect 42892 3664 42944 3670
rect 42892 3606 42944 3612
rect 42524 3596 42576 3602
rect 42524 3538 42576 3544
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 41524 3074 41552 3470
rect 42432 3392 42484 3398
rect 42432 3334 42484 3340
rect 41604 3120 41656 3126
rect 41524 3068 41604 3074
rect 41524 3062 41656 3068
rect 41236 3052 41288 3058
rect 41236 2994 41288 3000
rect 41524 3046 41644 3062
rect 42444 3058 42472 3334
rect 42432 3052 42484 3058
rect 41328 2984 41380 2990
rect 41326 2952 41328 2961
rect 41380 2952 41382 2961
rect 40408 2916 40460 2922
rect 41326 2887 41382 2896
rect 40408 2858 40460 2864
rect 40592 2848 40644 2854
rect 40592 2790 40644 2796
rect 40604 800 40632 2790
rect 41524 2514 41552 3046
rect 42432 2994 42484 3000
rect 41512 2508 41564 2514
rect 41512 2450 41564 2456
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 41248 800 41276 2382
rect 42536 800 42564 3538
rect 42892 2848 42944 2854
rect 42892 2790 42944 2796
rect 42904 2446 42932 2790
rect 42996 2650 43024 19314
rect 43456 19242 43484 19654
rect 43444 19236 43496 19242
rect 43444 19178 43496 19184
rect 43548 17678 43576 46310
rect 43824 45966 43852 49200
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 44468 45554 44496 49200
rect 45112 45626 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 44192 45526 44496 45554
rect 44192 45490 44220 45526
rect 44180 45484 44232 45490
rect 44180 45426 44232 45432
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 43996 45280 44048 45286
rect 43996 45222 44048 45228
rect 44008 29306 44036 45222
rect 44468 45082 44496 45358
rect 45112 45082 45140 45358
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 44916 44872 44968 44878
rect 44916 44814 44968 44820
rect 43996 29300 44048 29306
rect 43996 29242 44048 29248
rect 44928 26234 44956 44814
rect 45204 44402 45232 46990
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45388 45558 45416 46922
rect 45756 45966 45784 49200
rect 46296 46504 46348 46510
rect 46296 46446 46348 46452
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 45560 45824 45612 45830
rect 45560 45766 45612 45772
rect 45376 45552 45428 45558
rect 45376 45494 45428 45500
rect 45468 45280 45520 45286
rect 45468 45222 45520 45228
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 45376 29708 45428 29714
rect 45376 29650 45428 29656
rect 44836 26206 44956 26234
rect 44640 22636 44692 22642
rect 44640 22578 44692 22584
rect 43628 22024 43680 22030
rect 43628 21966 43680 21972
rect 43536 17672 43588 17678
rect 43536 17614 43588 17620
rect 43548 3942 43576 17614
rect 43640 12434 43668 21966
rect 44456 21956 44508 21962
rect 44456 21898 44508 21904
rect 44468 21690 44496 21898
rect 44652 21690 44680 22578
rect 44456 21684 44508 21690
rect 44456 21626 44508 21632
rect 44640 21684 44692 21690
rect 44640 21626 44692 21632
rect 44456 21548 44508 21554
rect 44456 21490 44508 21496
rect 44468 20602 44496 21490
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 44192 20466 44404 20482
rect 43812 20460 43864 20466
rect 43812 20402 43864 20408
rect 44180 20460 44404 20466
rect 44232 20454 44404 20460
rect 44180 20402 44232 20408
rect 43824 19768 43852 20402
rect 44376 20330 44404 20454
rect 44456 20392 44508 20398
rect 44454 20360 44456 20369
rect 44640 20392 44692 20398
rect 44508 20360 44510 20369
rect 44272 20324 44324 20330
rect 44272 20266 44324 20272
rect 44364 20324 44416 20330
rect 44640 20334 44692 20340
rect 44454 20295 44510 20304
rect 44364 20266 44416 20272
rect 44284 20058 44312 20266
rect 44272 20052 44324 20058
rect 44272 19994 44324 20000
rect 44652 19990 44680 20334
rect 44640 19984 44692 19990
rect 44640 19926 44692 19932
rect 43996 19848 44048 19854
rect 43996 19790 44048 19796
rect 43904 19780 43956 19786
rect 43824 19740 43904 19768
rect 43824 19514 43852 19740
rect 43904 19722 43956 19728
rect 43812 19508 43864 19514
rect 43812 19450 43864 19456
rect 43812 19168 43864 19174
rect 43812 19110 43864 19116
rect 43824 18766 43852 19110
rect 44008 18970 44036 19790
rect 43996 18964 44048 18970
rect 43996 18906 44048 18912
rect 43812 18760 43864 18766
rect 43812 18702 43864 18708
rect 43824 18290 43852 18702
rect 43812 18284 43864 18290
rect 43812 18226 43864 18232
rect 44456 18216 44508 18222
rect 44456 18158 44508 18164
rect 44468 17882 44496 18158
rect 44652 18154 44680 19926
rect 44640 18148 44692 18154
rect 44640 18090 44692 18096
rect 44456 17876 44508 17882
rect 44456 17818 44508 17824
rect 44272 17672 44324 17678
rect 44272 17614 44324 17620
rect 44284 17202 44312 17614
rect 44456 17604 44508 17610
rect 44456 17546 44508 17552
rect 44468 17202 44496 17546
rect 44836 17542 44864 26206
rect 45388 23798 45416 29650
rect 45376 23792 45428 23798
rect 45376 23734 45428 23740
rect 45480 23118 45508 45222
rect 45572 36922 45600 45766
rect 45652 45620 45704 45626
rect 45652 45562 45704 45568
rect 45664 45422 45692 45562
rect 45848 45554 45876 45902
rect 45756 45526 45876 45554
rect 45652 45416 45704 45422
rect 45652 45358 45704 45364
rect 45652 44872 45704 44878
rect 45652 44814 45704 44820
rect 45664 44334 45692 44814
rect 45756 44402 45784 45526
rect 46308 44538 46336 46446
rect 46400 45626 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46756 47116 46808 47122
rect 46756 47058 46808 47064
rect 46768 47025 46796 47058
rect 46754 47016 46810 47025
rect 46754 46951 46810 46960
rect 46756 46640 46808 46646
rect 46756 46582 46808 46588
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46388 45620 46440 45626
rect 46388 45562 46440 45568
rect 46492 45082 46520 45834
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 46296 44532 46348 44538
rect 46296 44474 46348 44480
rect 46020 44464 46072 44470
rect 46020 44406 46072 44412
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45652 44328 45704 44334
rect 45652 44270 45704 44276
rect 45560 36916 45612 36922
rect 45560 36858 45612 36864
rect 45664 26234 45692 44270
rect 45928 28076 45980 28082
rect 45928 28018 45980 28024
rect 45572 26206 45692 26234
rect 45468 23112 45520 23118
rect 45468 23054 45520 23060
rect 45192 22976 45244 22982
rect 45192 22918 45244 22924
rect 44916 22636 44968 22642
rect 44916 22578 44968 22584
rect 44928 22166 44956 22578
rect 44916 22160 44968 22166
rect 44916 22102 44968 22108
rect 45204 21962 45232 22918
rect 45376 22568 45428 22574
rect 45376 22510 45428 22516
rect 45284 22024 45336 22030
rect 45284 21966 45336 21972
rect 45192 21956 45244 21962
rect 45192 21898 45244 21904
rect 45296 21622 45324 21966
rect 45284 21616 45336 21622
rect 45284 21558 45336 21564
rect 45296 21146 45324 21558
rect 45284 21140 45336 21146
rect 45284 21082 45336 21088
rect 45388 20534 45416 22510
rect 45480 20942 45508 23054
rect 45468 20936 45520 20942
rect 45468 20878 45520 20884
rect 45376 20528 45428 20534
rect 45376 20470 45428 20476
rect 45100 20460 45152 20466
rect 45100 20402 45152 20408
rect 45112 19718 45140 20402
rect 45376 20324 45428 20330
rect 45376 20266 45428 20272
rect 45388 19990 45416 20266
rect 45376 19984 45428 19990
rect 45376 19926 45428 19932
rect 45100 19712 45152 19718
rect 45100 19654 45152 19660
rect 45388 19514 45416 19926
rect 45572 19718 45600 26206
rect 45744 23656 45796 23662
rect 45744 23598 45796 23604
rect 45756 23186 45784 23598
rect 45744 23180 45796 23186
rect 45744 23122 45796 23128
rect 45652 21956 45704 21962
rect 45652 21898 45704 21904
rect 45664 21554 45692 21898
rect 45652 21548 45704 21554
rect 45652 21490 45704 21496
rect 45560 19712 45612 19718
rect 45560 19654 45612 19660
rect 45376 19508 45428 19514
rect 45376 19450 45428 19456
rect 44916 19440 44968 19446
rect 44916 19382 44968 19388
rect 44928 18358 44956 19382
rect 45756 19310 45784 23122
rect 45836 23112 45888 23118
rect 45836 23054 45888 23060
rect 45848 20874 45876 23054
rect 45940 21894 45968 28018
rect 45928 21888 45980 21894
rect 45928 21830 45980 21836
rect 45836 20868 45888 20874
rect 45836 20810 45888 20816
rect 45100 19304 45152 19310
rect 45100 19246 45152 19252
rect 45744 19304 45796 19310
rect 45744 19246 45796 19252
rect 45112 18970 45140 19246
rect 45100 18964 45152 18970
rect 45100 18906 45152 18912
rect 45100 18828 45152 18834
rect 45100 18770 45152 18776
rect 45008 18760 45060 18766
rect 45008 18702 45060 18708
rect 44916 18352 44968 18358
rect 44916 18294 44968 18300
rect 45020 17610 45048 18702
rect 45112 18290 45140 18770
rect 45192 18760 45244 18766
rect 45192 18702 45244 18708
rect 45100 18284 45152 18290
rect 45100 18226 45152 18232
rect 45112 17882 45140 18226
rect 45100 17876 45152 17882
rect 45100 17818 45152 17824
rect 45204 17610 45232 18702
rect 45008 17604 45060 17610
rect 45008 17546 45060 17552
rect 45192 17604 45244 17610
rect 45192 17546 45244 17552
rect 44824 17536 44876 17542
rect 44824 17478 44876 17484
rect 45020 17338 45048 17546
rect 45008 17332 45060 17338
rect 45008 17274 45060 17280
rect 44272 17196 44324 17202
rect 44272 17138 44324 17144
rect 44456 17196 44508 17202
rect 44456 17138 44508 17144
rect 43640 12406 44036 12434
rect 44008 4554 44036 12406
rect 45204 7342 45232 17546
rect 45560 16516 45612 16522
rect 45560 16458 45612 16464
rect 45572 15745 45600 16458
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45652 10532 45704 10538
rect 45652 10474 45704 10480
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 45192 7336 45244 7342
rect 45192 7278 45244 7284
rect 45204 5098 45232 7278
rect 45664 5166 45692 10474
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45192 5092 45244 5098
rect 45192 5034 45244 5040
rect 45100 4820 45152 4826
rect 45100 4762 45152 4768
rect 43996 4548 44048 4554
rect 43996 4490 44048 4496
rect 44008 4078 44036 4490
rect 43904 4072 43956 4078
rect 43904 4014 43956 4020
rect 43996 4072 44048 4078
rect 43996 4014 44048 4020
rect 43536 3936 43588 3942
rect 43536 3878 43588 3884
rect 43168 3596 43220 3602
rect 43168 3538 43220 3544
rect 42984 2644 43036 2650
rect 42984 2586 43036 2592
rect 42892 2440 42944 2446
rect 42892 2382 42944 2388
rect 43180 800 43208 3538
rect 43916 2514 43944 4014
rect 44272 2984 44324 2990
rect 44270 2952 44272 2961
rect 44324 2952 44326 2961
rect 44270 2887 44326 2896
rect 43904 2508 43956 2514
rect 43904 2450 43956 2456
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 4762
rect 45664 4690 45692 5102
rect 45848 4826 45876 20810
rect 46032 20262 46060 44406
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46768 41138 46796 46582
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47768 46436 47820 46442
rect 47768 46378 47820 46384
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 47584 45484 47636 45490
rect 47584 45426 47636 45432
rect 47400 45416 47452 45422
rect 47400 45358 47452 45364
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 46940 44804 46992 44810
rect 46940 44746 46992 44752
rect 46952 44538 46980 44746
rect 46940 44532 46992 44538
rect 46940 44474 46992 44480
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 47412 42226 47440 45358
rect 47596 45014 47624 45426
rect 47584 45008 47636 45014
rect 47584 44950 47636 44956
rect 47400 42220 47452 42226
rect 47400 42162 47452 42168
rect 46756 41132 46808 41138
rect 46756 41074 46808 41080
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46662 39536 46718 39545
rect 46296 39500 46348 39506
rect 46662 39471 46718 39480
rect 46296 39442 46348 39448
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46308 37466 46336 38286
rect 46296 37460 46348 37466
rect 46296 37402 46348 37408
rect 46204 33856 46256 33862
rect 46204 33798 46256 33804
rect 46216 23338 46244 33798
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 32026 46336 32846
rect 46296 32020 46348 32026
rect 46296 31962 46348 31968
rect 46386 30016 46442 30025
rect 46386 29951 46442 29960
rect 46296 25696 46348 25702
rect 46296 25638 46348 25644
rect 46308 25362 46336 25638
rect 46296 25356 46348 25362
rect 46296 25298 46348 25304
rect 46400 24410 46428 29951
rect 46480 27872 46532 27878
rect 46480 27814 46532 27820
rect 46492 27538 46520 27814
rect 46480 27532 46532 27538
rect 46480 27474 46532 27480
rect 46572 24812 46624 24818
rect 46572 24754 46624 24760
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46388 24404 46440 24410
rect 46388 24346 46440 24352
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46584 24154 46612 24754
rect 46492 24126 46612 24154
rect 46216 23310 46428 23338
rect 46202 23216 46258 23225
rect 46202 23151 46258 23160
rect 46112 23044 46164 23050
rect 46112 22986 46164 22992
rect 46124 22545 46152 22986
rect 46216 22574 46244 23151
rect 46204 22568 46256 22574
rect 46110 22536 46166 22545
rect 46204 22510 46256 22516
rect 46110 22471 46166 22480
rect 46296 20936 46348 20942
rect 46296 20878 46348 20884
rect 46020 20256 46072 20262
rect 46020 20198 46072 20204
rect 46308 19242 46336 20878
rect 46400 19378 46428 23310
rect 46388 19372 46440 19378
rect 46388 19314 46440 19320
rect 46112 19236 46164 19242
rect 46112 19178 46164 19184
rect 46296 19236 46348 19242
rect 46296 19178 46348 19184
rect 46124 18850 46152 19178
rect 46492 18850 46520 24126
rect 46676 22098 46704 39471
rect 46940 39364 46992 39370
rect 46940 39306 46992 39312
rect 46952 39098 46980 39306
rect 46940 39092 46992 39098
rect 46940 39034 46992 39040
rect 46756 38956 46808 38962
rect 46756 38898 46808 38904
rect 46768 24886 46796 38898
rect 47308 35080 47360 35086
rect 47308 35022 47360 35028
rect 47320 34105 47348 35022
rect 47306 34096 47362 34105
rect 47306 34031 47362 34040
rect 46848 32428 46900 32434
rect 46848 32370 46900 32376
rect 46860 32337 46888 32370
rect 46846 32328 46902 32337
rect 46846 32263 46902 32272
rect 46848 32224 46900 32230
rect 46848 32166 46900 32172
rect 46860 31890 46888 32166
rect 46848 31884 46900 31890
rect 46848 31826 46900 31832
rect 46846 31376 46902 31385
rect 46846 31311 46902 31320
rect 46860 30394 46888 31311
rect 46848 30388 46900 30394
rect 46848 30330 46900 30336
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 46846 28656 46902 28665
rect 46846 28591 46902 28600
rect 46860 27130 46888 28591
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47044 27606 47072 27814
rect 47032 27600 47084 27606
rect 47032 27542 47084 27548
rect 46848 27124 46900 27130
rect 46848 27066 46900 27072
rect 46846 26616 46902 26625
rect 46846 26551 46902 26560
rect 46860 26450 46888 26551
rect 46848 26444 46900 26450
rect 46848 26386 46900 26392
rect 46846 25936 46902 25945
rect 46846 25871 46902 25880
rect 46756 24880 46808 24886
rect 46756 24822 46808 24828
rect 46756 24744 46808 24750
rect 46756 24686 46808 24692
rect 46768 23905 46796 24686
rect 46754 23896 46810 23905
rect 46754 23831 46810 23840
rect 46756 23656 46808 23662
rect 46756 23598 46808 23604
rect 46572 22092 46624 22098
rect 46572 22034 46624 22040
rect 46664 22092 46716 22098
rect 46664 22034 46716 22040
rect 46584 21350 46612 22034
rect 46572 21344 46624 21350
rect 46572 21286 46624 21292
rect 46124 18822 46520 18850
rect 45928 18284 45980 18290
rect 45928 18226 45980 18232
rect 45940 17270 45968 18226
rect 45928 17264 45980 17270
rect 45928 17206 45980 17212
rect 45836 4820 45888 4826
rect 45836 4762 45888 4768
rect 45652 4684 45704 4690
rect 45652 4626 45704 4632
rect 45192 4616 45244 4622
rect 45192 4558 45244 4564
rect 45204 3058 45232 4558
rect 45664 4214 45692 4626
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45652 4208 45704 4214
rect 45652 4150 45704 4156
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 45664 3534 45692 3606
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 46032 2446 46060 4490
rect 46124 4146 46152 18822
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46308 18290 46336 18702
rect 46386 18456 46442 18465
rect 46386 18391 46442 18400
rect 46296 18284 46348 18290
rect 46296 18226 46348 18232
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 17270 46336 17614
rect 46296 17264 46348 17270
rect 46296 17206 46348 17212
rect 46400 17202 46428 18391
rect 46388 17196 46440 17202
rect 46388 17138 46440 17144
rect 46204 17128 46256 17134
rect 46204 17070 46256 17076
rect 46216 5710 46244 17070
rect 46480 11552 46532 11558
rect 46480 11494 46532 11500
rect 46492 11218 46520 11494
rect 46480 11212 46532 11218
rect 46480 11154 46532 11160
rect 46388 10600 46440 10606
rect 46388 10542 46440 10548
rect 46400 8974 46428 10542
rect 46388 8968 46440 8974
rect 46388 8910 46440 8916
rect 46584 7954 46612 21286
rect 46768 20482 46796 23598
rect 46860 23186 46888 25871
rect 46848 23180 46900 23186
rect 46848 23122 46900 23128
rect 47308 20868 47360 20874
rect 47308 20810 47360 20816
rect 46676 20454 46796 20482
rect 46676 20398 46704 20454
rect 46664 20392 46716 20398
rect 46664 20334 46716 20340
rect 46676 19786 46704 20334
rect 46664 19780 46716 19786
rect 46664 19722 46716 19728
rect 46676 7954 46704 19722
rect 47032 19712 47084 19718
rect 47032 19654 47084 19660
rect 47044 19446 47072 19654
rect 47320 19514 47348 20810
rect 47308 19508 47360 19514
rect 47308 19450 47360 19456
rect 47032 19440 47084 19446
rect 47032 19382 47084 19388
rect 46756 19372 46808 19378
rect 46756 19314 46808 19320
rect 46768 10606 46796 19314
rect 47044 16794 47072 19382
rect 47412 18290 47440 42162
rect 47492 35080 47544 35086
rect 47492 35022 47544 35028
rect 47504 33930 47532 35022
rect 47492 33924 47544 33930
rect 47492 33866 47544 33872
rect 47596 32434 47624 44950
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47688 43858 47716 44134
rect 47676 43852 47728 43858
rect 47676 43794 47728 43800
rect 47780 43314 47808 46378
rect 47872 46345 47900 46514
rect 48044 46368 48096 46374
rect 47858 46336 47914 46345
rect 48044 46310 48096 46316
rect 47858 46271 47914 46280
rect 47768 43308 47820 43314
rect 47768 43250 47820 43256
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47676 38956 47728 38962
rect 47676 38898 47728 38904
rect 47688 38865 47716 38898
rect 47860 38888 47912 38894
rect 47674 38856 47730 38865
rect 47860 38830 47912 38836
rect 47674 38791 47730 38800
rect 47676 38276 47728 38282
rect 47676 38218 47728 38224
rect 47688 38010 47716 38218
rect 47676 38004 47728 38010
rect 47676 37946 47728 37952
rect 47872 35894 47900 38830
rect 47780 35866 47900 35894
rect 47676 32836 47728 32842
rect 47676 32778 47728 32784
rect 47688 32570 47716 32778
rect 47676 32564 47728 32570
rect 47676 32506 47728 32512
rect 47584 32428 47636 32434
rect 47584 32370 47636 32376
rect 47780 26234 47808 35866
rect 47952 34400 48004 34406
rect 47952 34342 48004 34348
rect 47860 34128 47912 34134
rect 47860 34070 47912 34076
rect 47872 33658 47900 34070
rect 47964 34066 47992 34342
rect 47952 34060 48004 34066
rect 47952 34002 48004 34008
rect 47860 33652 47912 33658
rect 47860 33594 47912 33600
rect 47860 33516 47912 33522
rect 47860 33458 47912 33464
rect 47872 33425 47900 33458
rect 47858 33416 47914 33425
rect 47858 33351 47914 33360
rect 47780 26206 47900 26234
rect 47676 25220 47728 25226
rect 47676 25162 47728 25168
rect 47688 24818 47716 25162
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47676 24812 47728 24818
rect 47676 24754 47728 24760
rect 47504 20369 47532 24754
rect 47768 24132 47820 24138
rect 47768 24074 47820 24080
rect 47780 23730 47808 24074
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47676 23044 47728 23050
rect 47676 22986 47728 22992
rect 47688 22778 47716 22986
rect 47676 22772 47728 22778
rect 47676 22714 47728 22720
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47596 20466 47624 22578
rect 47676 21956 47728 21962
rect 47676 21898 47728 21904
rect 47688 20602 47716 21898
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 47872 20534 47900 26206
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47964 21622 47992 21791
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 47860 20528 47912 20534
rect 47860 20470 47912 20476
rect 47584 20460 47636 20466
rect 47584 20402 47636 20408
rect 47490 20360 47546 20369
rect 47490 20295 47546 20304
rect 47400 18284 47452 18290
rect 47400 18226 47452 18232
rect 47400 17536 47452 17542
rect 47400 17478 47452 17484
rect 47412 17202 47440 17478
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 47032 16788 47084 16794
rect 47032 16730 47084 16736
rect 46848 16516 46900 16522
rect 46848 16458 46900 16464
rect 46860 16250 46888 16458
rect 46848 16244 46900 16250
rect 46848 16186 46900 16192
rect 47044 12434 47072 16730
rect 46952 12406 47072 12434
rect 46756 10600 46808 10606
rect 46756 10542 46808 10548
rect 46846 9616 46902 9625
rect 46846 9551 46902 9560
rect 46860 9042 46888 9551
rect 46848 9036 46900 9042
rect 46848 8978 46900 8984
rect 46952 8430 46980 12406
rect 47032 10124 47084 10130
rect 47032 10066 47084 10072
rect 47044 9586 47072 10066
rect 47032 9580 47084 9586
rect 47032 9522 47084 9528
rect 46940 8424 46992 8430
rect 46940 8366 46992 8372
rect 46572 7948 46624 7954
rect 46572 7890 46624 7896
rect 46664 7948 46716 7954
rect 46664 7890 46716 7896
rect 46204 5704 46256 5710
rect 46204 5646 46256 5652
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46112 4140 46164 4146
rect 46112 4082 46164 4088
rect 46308 3194 46336 4626
rect 46676 4570 46704 7890
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 46846 6216 46902 6225
rect 46846 6151 46902 6160
rect 46860 5778 46888 6151
rect 46848 5772 46900 5778
rect 46848 5714 46900 5720
rect 46584 4542 46704 4570
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46492 3602 46520 3878
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46296 3188 46348 3194
rect 46296 3130 46348 3136
rect 46584 2990 46612 4542
rect 46664 4140 46716 4146
rect 46664 4082 46716 4088
rect 46848 4140 46900 4146
rect 46848 4082 46900 4088
rect 46572 2984 46624 2990
rect 46572 2926 46624 2932
rect 46020 2440 46072 2446
rect 46020 2382 46072 2388
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45480 1970 45508 2246
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 46400 800 46428 2314
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46676 105 46704 4082
rect 46860 921 46888 4082
rect 47412 3670 47440 17138
rect 47504 9586 47532 20295
rect 47596 20058 47624 20402
rect 47584 20052 47636 20058
rect 47584 19994 47636 20000
rect 48056 19922 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48148 34610 48176 34711
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48136 25288 48188 25294
rect 48134 25256 48136 25265
rect 48188 25256 48190 25265
rect 48134 25191 48190 25200
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 19916 48096 19922
rect 48044 19858 48096 19864
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 47688 17338 47716 17546
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47780 16114 47808 16594
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47768 12640 47820 12646
rect 47768 12582 47820 12588
rect 47780 12306 47808 12582
rect 48134 12336 48190 12345
rect 47768 12300 47820 12306
rect 48134 12271 48136 12280
rect 47768 12242 47820 12248
rect 48188 12271 48190 12280
rect 48136 12242 48188 12248
rect 47676 12164 47728 12170
rect 47676 12106 47728 12112
rect 47688 11898 47716 12106
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47768 11076 47820 11082
rect 47768 11018 47820 11024
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 47780 10674 47808 11018
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47492 9580 47544 9586
rect 47492 9522 47544 9528
rect 47766 8936 47822 8945
rect 47766 8871 47822 8880
rect 47780 8566 47808 8871
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 47492 7812 47544 7818
rect 47492 7754 47544 7760
rect 47504 6866 47532 7754
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 47492 6860 47544 6866
rect 48134 6831 48190 6840
rect 47492 6802 47544 6808
rect 48136 6316 48188 6322
rect 48136 6258 48188 6264
rect 47952 6112 48004 6118
rect 47952 6054 48004 6060
rect 47964 5302 47992 6054
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 47400 3664 47452 3670
rect 47400 3606 47452 3612
rect 47766 3496 47822 3505
rect 47766 3431 47822 3440
rect 47780 3126 47808 3431
rect 47768 3120 47820 3126
rect 47768 3062 47820 3068
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 46846 912 46902 921
rect 46846 847 46902 856
rect 47044 800 47072 2450
rect 47688 800 47716 2926
rect 47872 1465 47900 5170
rect 48148 4185 48176 6258
rect 48134 4176 48190 4185
rect 48134 4111 48190 4120
rect 48044 3936 48096 3942
rect 48044 3878 48096 3884
rect 48056 3466 48084 3878
rect 48044 3460 48096 3466
rect 48044 3402 48096 3408
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48320 2372 48372 2378
rect 48320 2314 48372 2320
rect 47858 1456 47914 1465
rect 47858 1391 47914 1400
rect 48332 800 48360 2314
rect 48976 800 49004 3402
rect 46662 96 46718 105
rect 46662 31 46718 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3054 46960 3110 47016
rect 1398 42880 1454 42936
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1582 35400 1638 35456
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 32680 1638 32736
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1398 23160 1454 23216
rect 1398 17720 1454 17776
rect 1398 12280 1454 12336
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 2778 46280 2834 46336
rect 3330 44920 3386 44976
rect 2226 19080 2282 19136
rect 2778 36760 2834 36816
rect 3422 43560 3478 43616
rect 3514 39480 3570 39536
rect 2778 32000 2834 32056
rect 3146 28600 3202 28656
rect 3698 31320 3754 31376
rect 3422 19760 3478 19816
rect 3054 18400 3110 18456
rect 3054 17040 3110 17096
rect 2778 16360 2834 16416
rect 2778 15000 2834 15056
rect 3422 13640 3478 13696
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3514 10240 3570 10296
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4986 19896 5042 19952
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4066 7520 4122 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 8022 26152 8078 26208
rect 12346 26288 12402 26344
rect 12622 26152 12678 26208
rect 13174 26308 13230 26344
rect 13174 26288 13176 26308
rect 13176 26288 13228 26308
rect 13228 26288 13230 26308
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3440 4122 3496
rect 3790 1400 3846 1456
rect 3238 856 3294 912
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10690 18420 10746 18456
rect 10690 18400 10692 18420
rect 10692 18400 10744 18420
rect 10744 18400 10746 18420
rect 10782 18284 10838 18320
rect 12438 18420 12494 18456
rect 12438 18400 12440 18420
rect 12440 18400 12492 18420
rect 12492 18400 12494 18420
rect 10782 18264 10784 18284
rect 10784 18264 10836 18284
rect 10836 18264 10838 18284
rect 12806 18264 12862 18320
rect 14554 26288 14610 26344
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20258 35808 20314 35864
rect 20074 35672 20130 35728
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 16302 18808 16358 18864
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19982 30096 20038 30152
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19982 28636 19984 28656
rect 19984 28636 20036 28656
rect 20036 28636 20038 28656
rect 19982 28600 20038 28636
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 17038 20340 17040 20360
rect 17040 20340 17092 20360
rect 17092 20340 17094 20360
rect 17038 20304 17094 20340
rect 18418 18844 18420 18864
rect 18420 18844 18472 18864
rect 18472 18844 18474 18864
rect 18418 18808 18474 18844
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20902 33940 20904 33960
rect 20904 33940 20956 33960
rect 20956 33940 20958 33960
rect 20902 33904 20958 33940
rect 22006 33924 22062 33960
rect 22006 33904 22008 33924
rect 22008 33904 22060 33924
rect 22060 33904 22062 33924
rect 20350 32408 20406 32464
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 20258 16532 20260 16552
rect 20260 16532 20312 16552
rect 20312 16532 20314 16552
rect 20258 16496 20314 16532
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21086 30096 21142 30152
rect 21454 31900 21456 31920
rect 21456 31900 21508 31920
rect 21508 31900 21510 31920
rect 21454 31864 21510 31900
rect 22282 32000 22338 32056
rect 23570 31900 23572 31920
rect 23572 31900 23624 31920
rect 23624 31900 23626 31920
rect 23570 31864 23626 31900
rect 23570 28600 23626 28656
rect 23846 32428 23902 32464
rect 23846 32408 23848 32428
rect 23848 32408 23900 32428
rect 23900 32408 23902 32428
rect 24030 33904 24086 33960
rect 24122 32308 24124 32328
rect 24124 32308 24176 32328
rect 24176 32308 24178 32328
rect 24122 32272 24178 32308
rect 22650 19760 22706 19816
rect 23938 19760 23994 19816
rect 22834 16532 22836 16552
rect 22836 16532 22888 16552
rect 22888 16532 22890 16552
rect 22834 16496 22890 16532
rect 24306 16532 24308 16552
rect 24308 16532 24360 16552
rect 24360 16532 24362 16552
rect 24306 16496 24362 16532
rect 25962 35672 26018 35728
rect 26330 32292 26386 32328
rect 26330 32272 26332 32292
rect 26332 32272 26384 32292
rect 26384 32272 26386 32292
rect 25410 20304 25466 20360
rect 27894 35672 27950 35728
rect 27158 19896 27214 19952
rect 28630 35692 28686 35728
rect 28630 35672 28632 35692
rect 28632 35672 28684 35692
rect 28684 35672 28686 35692
rect 28906 32000 28962 32056
rect 28906 30096 28962 30152
rect 28998 24384 29054 24440
rect 30378 32136 30434 32192
rect 30286 31864 30342 31920
rect 29918 24404 29974 24440
rect 29918 24384 29920 24404
rect 29920 24384 29972 24404
rect 29972 24384 29974 24404
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 32494 32172 32496 32192
rect 32496 32172 32548 32192
rect 32548 32172 32550 32192
rect 32494 32136 32550 32172
rect 32402 31864 32458 31920
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 32678 31864 32734 31920
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 41326 2932 41328 2952
rect 41328 2932 41380 2952
rect 41380 2932 41382 2952
rect 41326 2896 41382 2932
rect 44454 20340 44456 20360
rect 44456 20340 44508 20360
rect 44508 20340 44510 20360
rect 44454 20304 44510 20340
rect 46846 47640 46902 47696
rect 46754 46960 46810 47016
rect 45558 15680 45614 15736
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 44270 2932 44272 2952
rect 44272 2932 44324 2952
rect 44324 2932 44326 2952
rect 44270 2896 44326 2932
rect 46662 39480 46718 39536
rect 46386 29960 46442 30016
rect 46202 23160 46258 23216
rect 46110 22480 46166 22536
rect 47306 34040 47362 34096
rect 46846 32272 46902 32328
rect 46846 31320 46902 31376
rect 47306 29280 47362 29336
rect 46846 28600 46902 28656
rect 46846 26560 46902 26616
rect 46846 25880 46902 25936
rect 46754 23840 46810 23896
rect 46386 18400 46442 18456
rect 47858 46280 47914 46336
rect 47950 40840 48006 40896
rect 47674 38800 47730 38856
rect 47858 33360 47914 33416
rect 47950 21800 48006 21856
rect 47490 20304 47546 20360
rect 46846 9560 46902 9616
rect 47306 7520 47362 7576
rect 46846 6160 46902 6216
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48134 32680 48190 32736
rect 48134 27920 48190 27976
rect 48134 25236 48136 25256
rect 48136 25236 48188 25256
rect 48188 25236 48190 25256
rect 48134 25200 48190 25236
rect 48134 24520 48190 24576
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12300 48190 12336
rect 48134 12280 48136 12300
rect 48136 12280 48188 12300
rect 48188 12280 48190 12300
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 47766 8880 47822 8936
rect 48134 6840 48190 6896
rect 47766 3440 47822 3496
rect 46846 856 46902 912
rect 48134 4120 48190 4176
rect 47858 1400 47914 1456
rect 46662 40 46718 96
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3049 47018 3115 47021
rect 0 47016 3115 47018
rect 0 46960 3054 47016
rect 3110 46960 3115 47016
rect 0 46958 3115 46960
rect 0 46868 800 46958
rect 3049 46955 3115 46958
rect 46749 47018 46815 47021
rect 49200 47018 50000 47108
rect 46749 47016 50000 47018
rect 46749 46960 46754 47016
rect 46810 46960 50000 47016
rect 46749 46958 50000 46960
rect 46749 46955 46815 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47853 46338 47919 46341
rect 49200 46338 50000 46428
rect 47853 46336 50000 46338
rect 47853 46280 47858 46336
rect 47914 46280 50000 46336
rect 47853 46278 50000 46280
rect 47853 46275 47919 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3325 44978 3391 44981
rect 0 44976 3391 44978
rect 0 44920 3330 44976
rect 3386 44920 3391 44976
rect 0 44918 3391 44920
rect 0 44828 800 44918
rect 3325 44915 3391 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3417 43618 3483 43621
rect 0 43616 3483 43618
rect 0 43560 3422 43616
rect 3478 43560 3483 43616
rect 0 43558 3483 43560
rect 0 43468 800 43558
rect 3417 43555 3483 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3509 39538 3575 39541
rect 0 39536 3575 39538
rect 0 39480 3514 39536
rect 3570 39480 3575 39536
rect 0 39478 3575 39480
rect 0 39388 800 39478
rect 3509 39475 3575 39478
rect 46657 39538 46723 39541
rect 49200 39538 50000 39628
rect 46657 39536 50000 39538
rect 46657 39480 46662 39536
rect 46718 39480 50000 39536
rect 46657 39478 50000 39480
rect 46657 39475 46723 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47669 38858 47735 38861
rect 49200 38858 50000 38948
rect 47669 38856 50000 38858
rect 47669 38800 47674 38856
rect 47730 38800 50000 38856
rect 47669 38798 50000 38800
rect 47669 38795 47735 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 20253 35866 20319 35869
rect 20118 35864 20319 35866
rect 20118 35808 20258 35864
rect 20314 35808 20319 35864
rect 20118 35806 20319 35808
rect 20118 35733 20178 35806
rect 20253 35803 20319 35806
rect 20069 35728 20178 35733
rect 20069 35672 20074 35728
rect 20130 35672 20178 35728
rect 20069 35670 20178 35672
rect 25957 35730 26023 35733
rect 27889 35730 27955 35733
rect 28625 35730 28691 35733
rect 25957 35728 28691 35730
rect 25957 35672 25962 35728
rect 26018 35672 27894 35728
rect 27950 35672 28630 35728
rect 28686 35672 28691 35728
rect 25957 35670 28691 35672
rect 20069 35667 20135 35670
rect 25957 35667 26023 35670
rect 27889 35667 27955 35670
rect 28625 35667 28691 35670
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 47301 34098 47367 34101
rect 49200 34098 50000 34188
rect 47301 34096 50000 34098
rect 47301 34040 47306 34096
rect 47362 34040 50000 34096
rect 47301 34038 50000 34040
rect 47301 34035 47367 34038
rect 20897 33962 20963 33965
rect 22001 33962 22067 33965
rect 24025 33962 24091 33965
rect 20897 33960 24091 33962
rect 20897 33904 20902 33960
rect 20958 33904 22006 33960
rect 22062 33904 24030 33960
rect 24086 33904 24091 33960
rect 49200 33948 50000 34038
rect 20897 33902 24091 33904
rect 20897 33899 20963 33902
rect 22001 33899 22067 33902
rect 24025 33899 24091 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47853 33418 47919 33421
rect 49200 33418 50000 33508
rect 47853 33416 50000 33418
rect 47853 33360 47858 33416
rect 47914 33360 50000 33416
rect 47853 33358 50000 33360
rect 47853 33355 47919 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 20345 32466 20411 32469
rect 23841 32466 23907 32469
rect 20345 32464 23907 32466
rect 20345 32408 20350 32464
rect 20406 32408 23846 32464
rect 23902 32408 23907 32464
rect 20345 32406 23907 32408
rect 20345 32403 20411 32406
rect 23841 32403 23907 32406
rect 24117 32330 24183 32333
rect 26325 32330 26391 32333
rect 24117 32328 26391 32330
rect 24117 32272 24122 32328
rect 24178 32272 26330 32328
rect 26386 32272 26391 32328
rect 24117 32270 26391 32272
rect 24117 32267 24183 32270
rect 26325 32267 26391 32270
rect 46841 32328 46907 32333
rect 46841 32272 46846 32328
rect 46902 32272 46907 32328
rect 46841 32267 46907 32272
rect 30373 32194 30439 32197
rect 32489 32194 32555 32197
rect 30373 32192 32555 32194
rect 0 32058 800 32148
rect 30373 32136 30378 32192
rect 30434 32136 32494 32192
rect 32550 32136 32555 32192
rect 30373 32134 32555 32136
rect 30373 32131 30439 32134
rect 32489 32131 32555 32134
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31908 800 31998
rect 2773 31995 2839 31998
rect 22277 32058 22343 32061
rect 28901 32058 28967 32061
rect 22277 32056 28967 32058
rect 22277 32000 22282 32056
rect 22338 32000 28906 32056
rect 28962 32000 28967 32056
rect 22277 31998 28967 32000
rect 46844 32058 46904 32267
rect 49200 32058 50000 32148
rect 46844 31998 50000 32058
rect 22277 31995 22343 31998
rect 28901 31995 28967 31998
rect 21449 31922 21515 31925
rect 23565 31922 23631 31925
rect 21449 31920 23631 31922
rect 21449 31864 21454 31920
rect 21510 31864 23570 31920
rect 23626 31864 23631 31920
rect 21449 31862 23631 31864
rect 21449 31859 21515 31862
rect 23565 31859 23631 31862
rect 30281 31922 30347 31925
rect 32397 31922 32463 31925
rect 32673 31922 32739 31925
rect 30281 31920 32739 31922
rect 30281 31864 30286 31920
rect 30342 31864 32402 31920
rect 32458 31864 32678 31920
rect 32734 31864 32739 31920
rect 49200 31908 50000 31998
rect 30281 31862 32739 31864
rect 30281 31859 30347 31862
rect 32397 31859 32463 31862
rect 32673 31859 32739 31862
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3693 31378 3759 31381
rect 0 31376 3759 31378
rect 0 31320 3698 31376
rect 3754 31320 3759 31376
rect 0 31318 3759 31320
rect 0 31228 800 31318
rect 3693 31315 3759 31318
rect 46841 31378 46907 31381
rect 49200 31378 50000 31468
rect 46841 31376 50000 31378
rect 46841 31320 46846 31376
rect 46902 31320 50000 31376
rect 46841 31318 50000 31320
rect 46841 31315 46907 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 19977 30154 20043 30157
rect 21081 30154 21147 30157
rect 28901 30154 28967 30157
rect 19977 30152 28967 30154
rect 0 29868 800 30108
rect 19977 30096 19982 30152
rect 20038 30096 21086 30152
rect 21142 30096 28906 30152
rect 28962 30096 28967 30152
rect 19977 30094 28967 30096
rect 19977 30091 20043 30094
rect 21081 30091 21147 30094
rect 28901 30091 28967 30094
rect 46381 30018 46447 30021
rect 49200 30018 50000 30108
rect 46381 30016 50000 30018
rect 46381 29960 46386 30016
rect 46442 29960 50000 30016
rect 46381 29958 50000 29960
rect 46381 29955 46447 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3141 28658 3207 28661
rect 0 28656 3207 28658
rect 0 28600 3146 28656
rect 3202 28600 3207 28656
rect 0 28598 3207 28600
rect 0 28508 800 28598
rect 3141 28595 3207 28598
rect 19977 28658 20043 28661
rect 23565 28658 23631 28661
rect 19977 28656 23631 28658
rect 19977 28600 19982 28656
rect 20038 28600 23570 28656
rect 23626 28600 23631 28656
rect 19977 28598 23631 28600
rect 19977 28595 20043 28598
rect 23565 28595 23631 28598
rect 46841 28658 46907 28661
rect 49200 28658 50000 28748
rect 46841 28656 50000 28658
rect 46841 28600 46846 28656
rect 46902 28600 50000 28656
rect 46841 28598 50000 28600
rect 46841 28595 46907 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 46841 26618 46907 26621
rect 49200 26618 50000 26708
rect 46841 26616 50000 26618
rect 46841 26560 46846 26616
rect 46902 26560 50000 26616
rect 46841 26558 50000 26560
rect 46841 26555 46907 26558
rect 49200 26468 50000 26558
rect 12341 26346 12407 26349
rect 13169 26346 13235 26349
rect 14549 26346 14615 26349
rect 12341 26344 14615 26346
rect 12341 26288 12346 26344
rect 12402 26288 13174 26344
rect 13230 26288 14554 26344
rect 14610 26288 14615 26344
rect 12341 26286 14615 26288
rect 12341 26283 12407 26286
rect 13169 26283 13235 26286
rect 14549 26283 14615 26286
rect 8017 26210 8083 26213
rect 12617 26210 12683 26213
rect 8017 26208 12683 26210
rect 8017 26152 8022 26208
rect 8078 26152 12622 26208
rect 12678 26152 12683 26208
rect 8017 26150 12683 26152
rect 8017 26147 8083 26150
rect 12617 26147 12683 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46841 25938 46907 25941
rect 49200 25938 50000 26028
rect 46841 25936 50000 25938
rect 46841 25880 46846 25936
rect 46902 25880 50000 25936
rect 46841 25878 50000 25880
rect 46841 25875 46907 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 48129 25258 48195 25261
rect 49200 25258 50000 25348
rect 48129 25256 50000 25258
rect 48129 25200 48134 25256
rect 48190 25200 50000 25256
rect 48129 25198 50000 25200
rect 48129 25195 48195 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 28993 24442 29059 24445
rect 29913 24442 29979 24445
rect 28993 24440 29979 24442
rect 28993 24384 28998 24440
rect 29054 24384 29918 24440
rect 29974 24384 29979 24440
rect 49200 24428 50000 24518
rect 28993 24382 29979 24384
rect 28993 24379 29059 24382
rect 29913 24379 29979 24382
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46749 23898 46815 23901
rect 49200 23898 50000 23988
rect 46749 23896 50000 23898
rect 46749 23840 46754 23896
rect 46810 23840 50000 23896
rect 46749 23838 50000 23840
rect 46749 23835 46815 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23068 800 23158
rect 1393 23155 1459 23158
rect 46197 23218 46263 23221
rect 49200 23218 50000 23308
rect 46197 23216 50000 23218
rect 46197 23160 46202 23216
rect 46258 23160 50000 23216
rect 46197 23158 50000 23160
rect 46197 23155 46263 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46105 22538 46171 22541
rect 49200 22538 50000 22628
rect 46105 22536 50000 22538
rect 46105 22480 46110 22536
rect 46166 22480 50000 22536
rect 46105 22478 50000 22480
rect 46105 22475 46171 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 47945 21858 48011 21861
rect 49200 21858 50000 21948
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 17033 20362 17099 20365
rect 25405 20362 25471 20365
rect 17033 20360 25471 20362
rect 17033 20304 17038 20360
rect 17094 20304 25410 20360
rect 25466 20304 25471 20360
rect 17033 20302 25471 20304
rect 17033 20299 17099 20302
rect 25405 20299 25471 20302
rect 44449 20362 44515 20365
rect 47485 20362 47551 20365
rect 44449 20360 47551 20362
rect 44449 20304 44454 20360
rect 44510 20304 47490 20360
rect 47546 20304 47551 20360
rect 44449 20302 47551 20304
rect 44449 20299 44515 20302
rect 47485 20299 47551 20302
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 4981 19954 5047 19957
rect 27153 19954 27219 19957
rect 4981 19952 27219 19954
rect 0 19818 800 19908
rect 4981 19896 4986 19952
rect 5042 19896 27158 19952
rect 27214 19896 27219 19952
rect 4981 19894 27219 19896
rect 4981 19891 5047 19894
rect 27153 19891 27219 19894
rect 3417 19818 3483 19821
rect 0 19816 3483 19818
rect 0 19760 3422 19816
rect 3478 19760 3483 19816
rect 0 19758 3483 19760
rect 0 19668 800 19758
rect 3417 19755 3483 19758
rect 22645 19818 22711 19821
rect 23933 19818 23999 19821
rect 22645 19816 23999 19818
rect 22645 19760 22650 19816
rect 22706 19760 23938 19816
rect 23994 19760 23999 19816
rect 22645 19758 23999 19760
rect 22645 19755 22711 19758
rect 23933 19755 23999 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 16297 18866 16363 18869
rect 18413 18866 18479 18869
rect 16297 18864 18479 18866
rect 16297 18808 16302 18864
rect 16358 18808 18418 18864
rect 18474 18808 18479 18864
rect 16297 18806 18479 18808
rect 16297 18803 16363 18806
rect 18413 18803 18479 18806
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3049 18458 3115 18461
rect 0 18456 3115 18458
rect 0 18400 3054 18456
rect 3110 18400 3115 18456
rect 0 18398 3115 18400
rect 0 18308 800 18398
rect 3049 18395 3115 18398
rect 10685 18458 10751 18461
rect 12433 18458 12499 18461
rect 10685 18456 12499 18458
rect 10685 18400 10690 18456
rect 10746 18400 12438 18456
rect 12494 18400 12499 18456
rect 10685 18398 12499 18400
rect 10685 18395 10751 18398
rect 12433 18395 12499 18398
rect 46381 18458 46447 18461
rect 49200 18458 50000 18548
rect 46381 18456 50000 18458
rect 46381 18400 46386 18456
rect 46442 18400 50000 18456
rect 46381 18398 50000 18400
rect 46381 18395 46447 18398
rect 10777 18322 10843 18325
rect 12801 18322 12867 18325
rect 10777 18320 12867 18322
rect 10777 18264 10782 18320
rect 10838 18264 12806 18320
rect 12862 18264 12867 18320
rect 49200 18308 50000 18398
rect 10777 18262 12867 18264
rect 10777 18259 10843 18262
rect 12801 18259 12867 18262
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3049 17098 3115 17101
rect 0 17096 3115 17098
rect 0 17040 3054 17096
rect 3110 17040 3115 17096
rect 0 17038 3115 17040
rect 0 16948 800 17038
rect 3049 17035 3115 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 20253 16554 20319 16557
rect 22829 16554 22895 16557
rect 24301 16554 24367 16557
rect 20253 16552 24367 16554
rect 0 16418 800 16508
rect 20253 16496 20258 16552
rect 20314 16496 22834 16552
rect 22890 16496 24306 16552
rect 24362 16496 24367 16552
rect 20253 16494 24367 16496
rect 20253 16491 20319 16494
rect 22829 16491 22895 16494
rect 24301 16491 24367 16494
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16268 800 16358
rect 2773 16355 2839 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13548 800 13638
rect 3417 13635 3483 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3509 10298 3575 10301
rect 0 10296 3575 10298
rect 0 10240 3514 10296
rect 3570 10240 3575 10296
rect 0 10238 3575 10240
rect 0 10148 800 10238
rect 3509 10235 3575 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 46841 9618 46907 9621
rect 49200 9618 50000 9708
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7428 800 7518
rect 4061 7515 4127 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6748 800 6838
rect 4061 6835 4127 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 46841 6218 46907 6221
rect 49200 6218 50000 6308
rect 46841 6216 50000 6218
rect 46841 6160 46846 6216
rect 46902 6160 50000 6216
rect 46841 6158 50000 6160
rect 46841 6155 46907 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 48129 4178 48195 4181
rect 49200 4178 50000 4268
rect 48129 4176 50000 4178
rect 48129 4120 48134 4176
rect 48190 4120 50000 4176
rect 48129 4118 50000 4120
rect 48129 4115 48195 4118
rect 49200 4028 50000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3348 800 3438
rect 4061 3435 4127 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 41321 2954 41387 2957
rect 44265 2954 44331 2957
rect 41321 2952 44331 2954
rect 0 2668 800 2908
rect 41321 2896 41326 2952
rect 41382 2896 44270 2952
rect 44326 2896 44331 2952
rect 41321 2894 44331 2896
rect 41321 2891 41387 2894
rect 44265 2891 44331 2894
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3785 1458 3851 1461
rect 0 1456 3851 1458
rect 0 1400 3790 1456
rect 3846 1400 3851 1456
rect 0 1398 3851 1400
rect 0 1308 800 1398
rect 3785 1395 3851 1398
rect 47853 1458 47919 1461
rect 49200 1458 50000 1548
rect 47853 1456 50000 1458
rect 47853 1400 47858 1456
rect 47914 1400 50000 1456
rect 47853 1398 50000 1400
rect 47853 1395 47919 1398
rect 49200 1308 50000 1398
rect 3233 914 3299 917
rect 2086 912 3299 914
rect 0 778 800 868
rect 2086 856 3238 912
rect 3294 856 3299 912
rect 2086 854 3299 856
rect 2086 778 2146 854
rect 3233 851 3299 854
rect 46841 914 46907 917
rect 46841 912 47042 914
rect 46841 856 46846 912
rect 46902 856 47042 912
rect 46841 854 47042 856
rect 46841 851 46907 854
rect 0 718 2146 778
rect 46982 778 47042 854
rect 49200 778 50000 868
rect 46982 718 50000 778
rect 0 628 800 718
rect 49200 628 50000 718
rect 46657 98 46723 101
rect 49200 98 50000 188
rect 46657 96 50000 98
rect 46657 40 46662 96
rect 46718 40 50000 96
rect 46657 38 50000 40
rect 46657 35 46723 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1644511149
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_269
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_186
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_194
timestamp 1644511149
transform 1 0 18952 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_319
timestamp 1644511149
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_368
timestamp 1644511149
transform 1 0 34960 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_380
timestamp 1644511149
transform 1 0 36064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_401
timestamp 1644511149
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_413
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1644511149
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1644511149
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1644511149
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_111
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_118
timestamp 1644511149
transform 1 0 11960 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1644511149
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1644511149
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_257
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_282
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1644511149
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_351
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_400
timestamp 1644511149
transform 1 0 37904 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_412
timestamp 1644511149
transform 1 0 39008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1644511149
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_239
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_251
timestamp 1644511149
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp 1644511149
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1644511149
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_345
timestamp 1644511149
transform 1 0 32844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_351
timestamp 1644511149
transform 1 0 33396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_363
timestamp 1644511149
transform 1 0 34500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_375
timestamp 1644511149
transform 1 0 35604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_423
timestamp 1644511149
transform 1 0 40020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_435
timestamp 1644511149
transform 1 0 41124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_454
timestamp 1644511149
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_479
timestamp 1644511149
transform 1 0 45172 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_487
timestamp 1644511149
transform 1 0 45908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1644511149
transform 1 0 46368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1644511149
transform 1 0 9660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1644511149
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1644511149
transform 1 0 11868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1644511149
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1644511149
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1644511149
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1644511149
transform 1 0 21528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_229
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1644511149
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_451
timestamp 1644511149
transform 1 0 42596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_455
timestamp 1644511149
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_467
timestamp 1644511149
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_482
timestamp 1644511149
transform 1 0 45448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_507
timestamp 1644511149
transform 1 0 47748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_515
timestamp 1644511149
transform 1 0 48484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1644511149
transform 1 0 16928 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1644511149
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_204
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1644511149
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1644511149
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_481
timestamp 1644511149
transform 1 0 45356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_495
timestamp 1644511149
transform 1 0 46644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_488
timestamp 1644511149
transform 1 0 46000 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_500
timestamp 1644511149
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_118
timestamp 1644511149
transform 1 0 11960 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1644511149
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1644511149
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1644511149
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_155
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_179
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1644511149
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1644511149
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1644511149
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1644511149
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1644511149
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1644511149
transform 1 0 16928 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1644511149
transform 1 0 18032 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1644511149
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1644511149
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1644511149
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1644511149
transform 1 0 16928 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_142
timestamp 1644511149
transform 1 0 14168 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_148
timestamp 1644511149
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_153
timestamp 1644511149
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1644511149
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_124
timestamp 1644511149
transform 1 0 12512 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_170
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_182
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1644511149
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1644511149
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_130
timestamp 1644511149
transform 1 0 13064 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_136
timestamp 1644511149
transform 1 0 13616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_140
timestamp 1644511149
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1644511149
transform 1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1644511149
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_180
timestamp 1644511149
transform 1 0 17664 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_197
timestamp 1644511149
transform 1 0 19228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_209
timestamp 1644511149
transform 1 0 20332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1644511149
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_493
timestamp 1644511149
transform 1 0 46460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_499
timestamp 1644511149
transform 1 0 47012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_128
timestamp 1644511149
transform 1 0 12880 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1644511149
transform 1 0 14352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_152
timestamp 1644511149
transform 1 0 15088 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_166
timestamp 1644511149
transform 1 0 16376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1644511149
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1644511149
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1644511149
transform 1 0 12420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 1644511149
transform 1 0 15088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_156
timestamp 1644511149
transform 1 0 15456 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1644511149
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_161
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_167
timestamp 1644511149
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_179
timestamp 1644511149
transform 1 0 17572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1644511149
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1644511149
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1644511149
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1644511149
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp 1644511149
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1644511149
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1644511149
transform 1 0 19688 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_214
timestamp 1644511149
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_226
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1644511149
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1644511149
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_176
timestamp 1644511149
transform 1 0 17296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1644511149
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1644511149
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1644511149
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1644511149
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1644511149
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1644511149
transform 1 0 11868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_124
timestamp 1644511149
transform 1 0 12512 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_136
timestamp 1644511149
transform 1 0 13616 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_144
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_152
timestamp 1644511149
transform 1 0 15088 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_174
timestamp 1644511149
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_194
timestamp 1644511149
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_198
timestamp 1644511149
transform 1 0 19320 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_233
timestamp 1644511149
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_265
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_269
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_315
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_327
timestamp 1644511149
transform 1 0 31188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_493
timestamp 1644511149
transform 1 0 46460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_499
timestamp 1644511149
transform 1 0 47012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_120
timestamp 1644511149
transform 1 0 12144 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1644511149
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_169
timestamp 1644511149
transform 1 0 16652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_181
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_202
timestamp 1644511149
transform 1 0 19688 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_208
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1644511149
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_256
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_268
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_290
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_298
timestamp 1644511149
transform 1 0 28520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_330
timestamp 1644511149
transform 1 0 31464 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_342
timestamp 1644511149
transform 1 0 32568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_354
timestamp 1644511149
transform 1 0 33672 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1644511149
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1644511149
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1644511149
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_191
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_242
timestamp 1644511149
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_250
timestamp 1644511149
transform 1 0 24104 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_262
timestamp 1644511149
transform 1 0 25208 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1644511149
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_284
timestamp 1644511149
transform 1 0 27232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_308
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_320
timestamp 1644511149
transform 1 0 30544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_472
timestamp 1644511149
transform 1 0 44528 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_484
timestamp 1644511149
transform 1 0 45632 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_493
timestamp 1644511149
transform 1 0 46460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_11
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1644511149
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1644511149
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_181
timestamp 1644511149
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_276
timestamp 1644511149
transform 1 0 26496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_292
timestamp 1644511149
transform 1 0 27968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_300
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1644511149
transform 1 0 31188 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1644511149
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_465
timestamp 1644511149
transform 1 0 43884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_482
timestamp 1644511149
transform 1 0 45448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_490
timestamp 1644511149
transform 1 0 46184 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_14
timestamp 1644511149
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1644511149
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_100
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_104
timestamp 1644511149
transform 1 0 10672 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1644511149
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_173
timestamp 1644511149
transform 1 0 17020 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1644511149
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_187
timestamp 1644511149
transform 1 0 18308 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_199
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_207
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1644511149
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_228
timestamp 1644511149
transform 1 0 22080 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_240
timestamp 1644511149
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_252
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_268
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_304
timestamp 1644511149
transform 1 0 29072 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1644511149
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_358
timestamp 1644511149
transform 1 0 34040 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_370
timestamp 1644511149
transform 1 0 35144 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_382
timestamp 1644511149
transform 1 0 36248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1644511149
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_465
timestamp 1644511149
transform 1 0 43884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_483
timestamp 1644511149
transform 1 0 45540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_492
timestamp 1644511149
transform 1 0 46368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_496
timestamp 1644511149
transform 1 0 46736 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_162
timestamp 1644511149
transform 1 0 16008 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1644511149
transform 1 0 25300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_327
timestamp 1644511149
transform 1 0 31188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_353
timestamp 1644511149
transform 1 0 33580 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1644511149
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_462
timestamp 1644511149
transform 1 0 43608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1644511149
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_482
timestamp 1644511149
transform 1 0 45448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_490
timestamp 1644511149
transform 1 0 46184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_96
timestamp 1644511149
transform 1 0 9936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_127
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_134
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1644511149
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_260
timestamp 1644511149
transform 1 0 25024 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_266
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_288
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_318
timestamp 1644511149
transform 1 0 30360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_352
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_364
timestamp 1644511149
transform 1 0 34592 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_376
timestamp 1644511149
transform 1 0 35696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1644511149
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_434
timestamp 1644511149
transform 1 0 41032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1644511149
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_468
timestamp 1644511149
transform 1 0 44160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_492
timestamp 1644511149
transform 1 0 46368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_496
timestamp 1644511149
transform 1 0 46736 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1644511149
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_89
timestamp 1644511149
transform 1 0 9292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_113
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1644511149
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1644511149
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1644511149
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1644511149
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_263
timestamp 1644511149
transform 1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_279
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_317
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_429
timestamp 1644511149
transform 1 0 40572 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_452
timestamp 1644511149
transform 1 0 42688 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_458
timestamp 1644511149
transform 1 0 43240 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_483
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1644511149
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1644511149
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_124
timestamp 1644511149
transform 1 0 12512 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_146
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_152
timestamp 1644511149
transform 1 0 15088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_207
timestamp 1644511149
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1644511149
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1644511149
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_260
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1644511149
transform 1 0 25760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1644511149
transform 1 0 29624 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1644511149
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_475
timestamp 1644511149
transform 1 0 44804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_114
timestamp 1644511149
transform 1 0 11592 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_126
timestamp 1644511149
transform 1 0 12696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1644511149
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_162
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_206
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1644511149
transform 1 0 21988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1644511149
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_256
timestamp 1644511149
transform 1 0 24656 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1644511149
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 1644511149
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_330
timestamp 1644511149
transform 1 0 31464 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_342
timestamp 1644511149
transform 1 0 32568 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_486
timestamp 1644511149
transform 1 0 45816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_490
timestamp 1644511149
transform 1 0 46184 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1644511149
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_104
timestamp 1644511149
transform 1 0 10672 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_121
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_133
timestamp 1644511149
transform 1 0 13340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_141
timestamp 1644511149
transform 1 0 14076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_151
timestamp 1644511149
transform 1 0 14996 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_172
timestamp 1644511149
transform 1 0 16928 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_179
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_191
timestamp 1644511149
transform 1 0 18676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_257
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_298
timestamp 1644511149
transform 1 0 28520 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_315
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_434
timestamp 1644511149
transform 1 0 41032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1644511149
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_465
timestamp 1644511149
transform 1 0 43884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_474
timestamp 1644511149
transform 1 0 44712 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1644511149
transform 1 0 12420 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1644511149
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_173
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_232
timestamp 1644511149
transform 1 0 22448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_257
timestamp 1644511149
transform 1 0 24748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_286
timestamp 1644511149
transform 1 0 27416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_296
timestamp 1644511149
transform 1 0 28336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1644511149
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_330
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_342
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_485
timestamp 1644511149
transform 1 0 45724 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_119
timestamp 1644511149
transform 1 0 12052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1644511149
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_197
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1644511149
transform 1 0 19596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_309
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1644511149
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_486
timestamp 1644511149
transform 1 0 45816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_102
timestamp 1644511149
transform 1 0 10488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_110
timestamp 1644511149
transform 1 0 11224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_174
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1644511149
transform 1 0 19596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_225
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1644511149
transform 1 0 22356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_238
timestamp 1644511149
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1644511149
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_484
timestamp 1644511149
transform 1 0 45632 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_490
timestamp 1644511149
transform 1 0 46184 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_77
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_82
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_94
timestamp 1644511149
transform 1 0 9752 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1644511149
transform 1 0 11960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_122
timestamp 1644511149
transform 1 0 12328 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_150
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1644511149
transform 1 0 19136 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_263
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_325
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1644511149
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_98
timestamp 1644511149
transform 1 0 10120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_110
timestamp 1644511149
transform 1 0 11224 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_126
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1644511149
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_159
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_276
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_284
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1644511149
transform 1 0 30084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1644511149
transform 1 0 31188 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1644511149
transform 1 0 32292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_75
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1644511149
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_104
timestamp 1644511149
transform 1 0 10672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1644511149
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1644511149
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_148
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_156
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_173
timestamp 1644511149
transform 1 0 17020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_215
timestamp 1644511149
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_325
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1644511149
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_100
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_116
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_154
timestamp 1644511149
transform 1 0 15272 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_216
timestamp 1644511149
transform 1 0 20976 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1644511149
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_235
timestamp 1644511149
transform 1 0 22724 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_269
timestamp 1644511149
transform 1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_282
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_316
timestamp 1644511149
transform 1 0 30176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_323
timestamp 1644511149
transform 1 0 30820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_335
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_347
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_359
timestamp 1644511149
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_96
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_100
timestamp 1644511149
transform 1 0 10304 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1644511149
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_135
timestamp 1644511149
transform 1 0 13524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 1644511149
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_265
timestamp 1644511149
transform 1 0 25484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_288
timestamp 1644511149
transform 1 0 27600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_300
timestamp 1644511149
transform 1 0 28704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1644511149
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1644511149
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_111
timestamp 1644511149
transform 1 0 11316 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_119
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1644511149
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_150
timestamp 1644511149
transform 1 0 14904 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_162
timestamp 1644511149
transform 1 0 16008 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_174
timestamp 1644511149
transform 1 0 17112 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_186
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_238
timestamp 1644511149
transform 1 0 23000 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_273
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_328
timestamp 1644511149
transform 1 0 31280 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_340
timestamp 1644511149
transform 1 0 32384 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_352
timestamp 1644511149
transform 1 0 33488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1644511149
transform 1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1644511149
transform 1 0 12788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_139
timestamp 1644511149
transform 1 0 13892 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_147
timestamp 1644511149
transform 1 0 14628 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1644511149
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_209
timestamp 1644511149
transform 1 0 20332 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_244
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_260
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_268
timestamp 1644511149
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1644511149
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_308
timestamp 1644511149
transform 1 0 29440 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_340
timestamp 1644511149
transform 1 0 32384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_352
timestamp 1644511149
transform 1 0 33488 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_364
timestamp 1644511149
transform 1 0 34592 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_376
timestamp 1644511149
transform 1 0 35696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1644511149
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_115
timestamp 1644511149
transform 1 0 11684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1644511149
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_144
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_148
timestamp 1644511149
transform 1 0 14720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_170
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_200
timestamp 1644511149
transform 1 0 19504 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_208
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1644511149
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1644511149
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp 1644511149
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_316
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_324
timestamp 1644511149
transform 1 0 30912 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_142
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_154
timestamp 1644511149
transform 1 0 15272 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_214
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_238
timestamp 1644511149
transform 1 0 23000 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_246
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1644511149
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_265
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_285
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_294
timestamp 1644511149
transform 1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_304
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_313
timestamp 1644511149
transform 1 0 29900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_342
timestamp 1644511149
transform 1 0 32568 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_354
timestamp 1644511149
transform 1 0 33672 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_366
timestamp 1644511149
transform 1 0 34776 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_378
timestamp 1644511149
transform 1 0 35880 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1644511149
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_493
timestamp 1644511149
transform 1 0 46460 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_499
timestamp 1644511149
transform 1 0 47012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_150
timestamp 1644511149
transform 1 0 14904 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_154
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_176
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_203
timestamp 1644511149
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_211
timestamp 1644511149
transform 1 0 20516 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_239
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1644511149
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_262
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_281
timestamp 1644511149
transform 1 0 26956 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_330
timestamp 1644511149
transform 1 0 31464 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_342
timestamp 1644511149
transform 1 0 32568 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_354
timestamp 1644511149
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1644511149
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_213
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1644511149
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1644511149
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_247
timestamp 1644511149
transform 1 0 23828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_267
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1644511149
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_288
timestamp 1644511149
transform 1 0 27600 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_296
timestamp 1644511149
transform 1 0 28336 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_306
timestamp 1644511149
transform 1 0 29256 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_230
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_242
timestamp 1644511149
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1644511149
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_256
timestamp 1644511149
transform 1 0 24656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_264
timestamp 1644511149
transform 1 0 25392 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_272
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_276
timestamp 1644511149
transform 1 0 26496 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_288
timestamp 1644511149
transform 1 0 27600 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_299
timestamp 1644511149
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_325
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_337
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_202
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_228
timestamp 1644511149
transform 1 0 22080 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_260
timestamp 1644511149
transform 1 0 25024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_291
timestamp 1644511149
transform 1 0 27876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_303
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_319
timestamp 1644511149
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1644511149
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1644511149
transform 1 0 33764 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1644511149
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_185
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1644511149
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_203
timestamp 1644511149
transform 1 0 19780 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_207
timestamp 1644511149
transform 1 0 20148 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1644511149
transform 1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_256
timestamp 1644511149
transform 1 0 24656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_268
timestamp 1644511149
transform 1 0 25760 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_290
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1644511149
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_325
timestamp 1644511149
transform 1 0 31004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_344
timestamp 1644511149
transform 1 0 32752 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_350
timestamp 1644511149
transform 1 0 33304 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_175
timestamp 1644511149
transform 1 0 17204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_207
timestamp 1644511149
transform 1 0 20148 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_211
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1644511149
transform 1 0 22172 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_236
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_259
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_269
timestamp 1644511149
transform 1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1644511149
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1644511149
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_308
timestamp 1644511149
transform 1 0 29440 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_320
timestamp 1644511149
transform 1 0 30544 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 1644511149
transform 1 0 32476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1644511149
transform 1 0 34408 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_371
timestamp 1644511149
transform 1 0 35236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_378
timestamp 1644511149
transform 1 0 35880 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1644511149
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_10
timestamp 1644511149
transform 1 0 2024 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_14
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1644511149
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_216
timestamp 1644511149
transform 1 0 20976 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_228
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_232
timestamp 1644511149
transform 1 0 22448 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_267
timestamp 1644511149
transform 1 0 25668 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_273
timestamp 1644511149
transform 1 0 26220 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_331
timestamp 1644511149
transform 1 0 31556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_337
timestamp 1644511149
transform 1 0 32108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_347
timestamp 1644511149
transform 1 0 33028 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1644511149
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_372
timestamp 1644511149
transform 1 0 35328 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_383
timestamp 1644511149
transform 1 0 36340 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_395
timestamp 1644511149
transform 1 0 37444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_407
timestamp 1644511149
transform 1 0 38548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_507
timestamp 1644511149
transform 1 0 47748 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_515
timestamp 1644511149
transform 1 0 48484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1644511149
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1644511149
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1644511149
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_190
timestamp 1644511149
transform 1 0 18584 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_214
timestamp 1644511149
transform 1 0 20792 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1644511149
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_241
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_251
timestamp 1644511149
transform 1 0 24196 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1644511149
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_287
timestamp 1644511149
transform 1 0 27508 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1644511149
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_303
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_311
timestamp 1644511149
transform 1 0 29716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_347
timestamp 1644511149
transform 1 0 33028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_356
timestamp 1644511149
transform 1 0 33856 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_364
timestamp 1644511149
transform 1 0 34592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1644511149
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_171
timestamp 1644511149
transform 1 0 16836 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_200
timestamp 1644511149
transform 1 0 19504 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_208
timestamp 1644511149
transform 1 0 20240 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1644511149
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_224
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_232
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 1644511149
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1644511149
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_266
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_274
timestamp 1644511149
transform 1 0 26312 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_286
timestamp 1644511149
transform 1 0 27416 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_313
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_324
timestamp 1644511149
transform 1 0 30912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_334
timestamp 1644511149
transform 1 0 31832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_341
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1644511149
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1644511149
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_373
timestamp 1644511149
transform 1 0 35420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_380
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_392
timestamp 1644511149
transform 1 0 37168 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_404
timestamp 1644511149
transform 1 0 38272 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_416
timestamp 1644511149
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_209
timestamp 1644511149
transform 1 0 20332 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_245
timestamp 1644511149
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_256
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_268
timestamp 1644511149
transform 1 0 25760 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1644511149
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_301
timestamp 1644511149
transform 1 0 28796 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_313
timestamp 1644511149
transform 1 0 29900 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_325
timestamp 1644511149
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1644511149
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_369
timestamp 1644511149
transform 1 0 35052 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_381
timestamp 1644511149
transform 1 0 36156 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1644511149
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_201
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_220
timestamp 1644511149
transform 1 0 21344 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_232
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_270
timestamp 1644511149
transform 1 0 25944 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_278
timestamp 1644511149
transform 1 0 26680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_284
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_296
timestamp 1644511149
transform 1 0 28336 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_372
timestamp 1644511149
transform 1 0 35328 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_383
timestamp 1644511149
transform 1 0 36340 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_395
timestamp 1644511149
transform 1 0 37444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_407
timestamp 1644511149
transform 1 0 38548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_189
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1644511149
transform 1 0 19136 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1644511149
transform 1 0 20240 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_246
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_250
timestamp 1644511149
transform 1 0 24104 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_290
timestamp 1644511149
transform 1 0 27784 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_294
timestamp 1644511149
transform 1 0 28152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1644511149
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1644511149
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_356
timestamp 1644511149
transform 1 0 33856 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_377
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1644511149
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_10
timestamp 1644511149
transform 1 0 2024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_14
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_203
timestamp 1644511149
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_207
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_219
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_246
timestamp 1644511149
transform 1 0 23736 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_298
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1644511149
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_330
timestamp 1644511149
transform 1 0 31464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_341
timestamp 1644511149
transform 1 0 32476 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1644511149
transform 1 0 33396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_371
timestamp 1644511149
transform 1 0 35236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_378
timestamp 1644511149
transform 1 0 35880 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_390
timestamp 1644511149
transform 1 0 36984 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_402
timestamp 1644511149
transform 1 0 38088 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_414
timestamp 1644511149
transform 1 0 39192 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1644511149
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1644511149
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1644511149
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1644511149
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_232
timestamp 1644511149
transform 1 0 22448 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_244
timestamp 1644511149
transform 1 0 23552 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_256
timestamp 1644511149
transform 1 0 24656 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1644511149
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_302
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_312
timestamp 1644511149
transform 1 0 29808 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_324
timestamp 1644511149
transform 1 0 30912 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_328
timestamp 1644511149
transform 1 0 31280 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_358
timestamp 1644511149
transform 1 0 34040 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_370
timestamp 1644511149
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_382
timestamp 1644511149
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1644511149
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_213
timestamp 1644511149
transform 1 0 20700 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_217
timestamp 1644511149
transform 1 0 21068 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_225
timestamp 1644511149
transform 1 0 21804 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_236
timestamp 1644511149
transform 1 0 22816 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_263
timestamp 1644511149
transform 1 0 25300 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_283
timestamp 1644511149
transform 1 0 27140 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_291
timestamp 1644511149
transform 1 0 27876 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_313
timestamp 1644511149
transform 1 0 29900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1644511149
transform 1 0 32108 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1644511149
transform 1 0 33212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_361
timestamp 1644511149
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_253
timestamp 1644511149
transform 1 0 24380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1644511149
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1644511149
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_229
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_267
timestamp 1644511149
transform 1 0 25668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1644511149
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1644511149
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_507
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_253
timestamp 1644511149
transform 1 0 24380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_265
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_277
timestamp 1644511149
transform 1 0 26588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_301
timestamp 1644511149
transform 1 0 28796 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_313
timestamp 1644511149
transform 1 0 29900 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_325
timestamp 1644511149
transform 1 0 31004 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_333
timestamp 1644511149
transform 1 0 31740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_229
timestamp 1644511149
transform 1 0 22172 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_235
timestamp 1644511149
transform 1 0 22724 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_271
timestamp 1644511149
transform 1 0 26036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_275
timestamp 1644511149
transform 1 0 26404 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_279
timestamp 1644511149
transform 1 0 26772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_290
timestamp 1644511149
transform 1 0 27784 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_302
timestamp 1644511149
transform 1 0 28888 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1644511149
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_451
timestamp 1644511149
transform 1 0 42596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_455
timestamp 1644511149
transform 1 0 42964 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_467
timestamp 1644511149
transform 1 0 44068 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1644511149
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1644511149
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1644511149
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_140
timestamp 1644511149
transform 1 0 13984 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_152
timestamp 1644511149
transform 1 0 15088 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_209
timestamp 1644511149
transform 1 0 20332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_265
timestamp 1644511149
transform 1 0 25484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_277
timestamp 1644511149
transform 1 0 26588 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_340
timestamp 1644511149
transform 1 0 32384 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_455
timestamp 1644511149
transform 1 0 42964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_463
timestamp 1644511149
transform 1 0 43700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_468
timestamp 1644511149
transform 1 0 44160 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1644511149
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1644511149
transform 1 0 5152 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1644511149
transform 1 0 6256 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1644511149
transform 1 0 7360 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1644511149
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_112
timestamp 1644511149
transform 1 0 11408 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_124
timestamp 1644511149
transform 1 0 12512 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_205
timestamp 1644511149
transform 1 0 19964 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1644511149
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_14
timestamp 1644511149
transform 1 0 2392 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_21
timestamp 1644511149
transform 1 0 3036 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1644511149
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1644511149
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_316
timestamp 1644511149
transform 1 0 30176 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_328
timestamp 1644511149
transform 1 0 31280 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_9
timestamp 1644511149
transform 1 0 1932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_16
timestamp 1644511149
transform 1 0 2576 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_91
timestamp 1644511149
transform 1 0 9476 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_103
timestamp 1644511149
transform 1 0 10580 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_157
timestamp 1644511149
transform 1 0 15548 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1644511149
transform 1 0 24840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1644511149
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0567_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27416 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0573_
timestamp 1644511149
transform 1 0 26036 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0574_
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0575_
timestamp 1644511149
transform 1 0 27232 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0576_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0577_
timestamp 1644511149
transform 1 0 22816 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0579_
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0581_
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0582_
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0583_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0584_
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0589_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0590_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0591_
timestamp 1644511149
transform 1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0592_
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0594_
timestamp 1644511149
transform 1 0 14260 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0595_
timestamp 1644511149
transform 1 0 15272 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0596_
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0599_
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0602_
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0603_
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0608_
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0610_
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0611_
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0612_
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0613_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0615_
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1644511149
transform 1 0 22724 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0617_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0618_
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0620_
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1644511149
transform 1 0 18216 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0622_
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0624_
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0625_
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0628_
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0631_
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0633_
timestamp 1644511149
transform 1 0 15088 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1644511149
transform 1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13800 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12972 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1644511149
transform 1 0 14996 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0638_
timestamp 1644511149
transform 1 0 12972 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0639_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1644511149
transform 1 0 12512 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0644_
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0645_
timestamp 1644511149
transform 1 0 12052 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0646_
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0648_
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1644511149
transform 1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0650_
timestamp 1644511149
transform 1 0 11592 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0651_
timestamp 1644511149
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0652_
timestamp 1644511149
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0653_
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1644511149
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0655_
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0658_
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9752 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0662_
timestamp 1644511149
transform 1 0 7820 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0665_
timestamp 1644511149
transform 1 0 12328 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0666_
timestamp 1644511149
transform 1 0 10764 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0669_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0670_
timestamp 1644511149
transform 1 0 12512 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0672_
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 1644511149
transform 1 0 11868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1644511149
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0675_
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0677_
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0678_
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0679_
timestamp 1644511149
transform 1 0 12420 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0680_
timestamp 1644511149
transform 1 0 11868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0682_
timestamp 1644511149
transform 1 0 19320 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1644511149
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0685_
timestamp 1644511149
transform 1 0 11868 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1644511149
transform 1 0 11776 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0689_
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0690_
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1644511149
transform 1 0 15180 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0693_
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0695_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0696_
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0700_
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0701_
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0703_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1644511149
transform 1 0 17480 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0705_
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0706_
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0707_
timestamp 1644511149
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0708_
timestamp 1644511149
transform 1 0 22264 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1644511149
transform 1 0 26036 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0712_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0715_
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0717_
timestamp 1644511149
transform 1 0 22448 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0718_
timestamp 1644511149
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1644511149
transform 1 0 21344 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0721_
timestamp 1644511149
transform 1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_1  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0723_
timestamp 1644511149
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0725_
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0726_
timestamp 1644511149
transform 1 0 28336 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0728_
timestamp 1644511149
transform 1 0 20884 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0730_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0733_
timestamp 1644511149
transform 1 0 25024 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0734_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0735_
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0736_
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0737_
timestamp 1644511149
transform 1 0 22448 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0738_
timestamp 1644511149
transform 1 0 25576 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0739_
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0741_
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0743_
timestamp 1644511149
transform 1 0 20884 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0746_
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0747_
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1644511149
transform 1 0 20976 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0750_
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0751_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0752_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0753_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0754_
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0755_
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0756_
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0758_
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0759_
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0760_
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0762_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0766_
timestamp 1644511149
transform 1 0 21712 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0767_
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0771_
timestamp 1644511149
transform 1 0 30084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0772_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0773_
timestamp 1644511149
transform 1 0 32200 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0774_
timestamp 1644511149
transform 1 0 30912 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0775_
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0776_
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0778_
timestamp 1644511149
transform 1 0 31280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1644511149
transform 1 0 27876 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0780_
timestamp 1644511149
transform 1 0 34776 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0781_
timestamp 1644511149
transform 1 0 33396 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0782_
timestamp 1644511149
transform 1 0 32108 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0783_
timestamp 1644511149
transform 1 0 32384 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0784_
timestamp 1644511149
transform 1 0 33396 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0785_
timestamp 1644511149
transform 1 0 32384 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0786_
timestamp 1644511149
transform 1 0 32200 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0788_
timestamp 1644511149
transform 1 0 35604 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0789_
timestamp 1644511149
transform 1 0 35696 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0790_
timestamp 1644511149
transform 1 0 34868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0792_
timestamp 1644511149
transform 1 0 35696 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0793_
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0794_
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1644511149
transform 1 0 27048 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0796_
timestamp 1644511149
transform 1 0 26772 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0797_
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0798_
timestamp 1644511149
transform 1 0 24840 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1644511149
transform 1 0 26956 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 1644511149
transform 1 0 26128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0802_
timestamp 1644511149
transform 1 0 23092 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0804_
timestamp 1644511149
transform 1 0 23184 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0805_
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1644511149
transform 1 0 29256 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0807_
timestamp 1644511149
transform 1 0 28060 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0808_
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1644511149
transform 1 0 31832 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0810_
timestamp 1644511149
transform 1 0 32844 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0811_
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0812_
timestamp 1644511149
transform 1 0 27508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0813_
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0814_
timestamp 1644511149
transform 1 0 27232 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0815_
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0816_
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0817_
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0818_
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0819_
timestamp 1644511149
transform 1 0 25668 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0820_
timestamp 1644511149
transform 1 0 25392 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0821_
timestamp 1644511149
transform 1 0 24472 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0822_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1644511149
transform 1 0 22448 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0825_
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0827_
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 1644511149
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1644511149
transform 1 0 29440 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0831_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0832_
timestamp 1644511149
transform 1 0 28612 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0833_
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0835_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0836_
timestamp 1644511149
transform 1 0 26404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0837_
timestamp 1644511149
transform 1 0 28612 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0838_
timestamp 1644511149
transform 1 0 28152 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0839_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1644511149
transform 1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0842_
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0843_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0844_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0845_
timestamp 1644511149
transform 1 0 27416 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0846_
timestamp 1644511149
transform 1 0 27508 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0847_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1644511149
transform 1 0 27232 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0849_
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0852_
timestamp 1644511149
transform 1 0 25576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1644511149
transform 1 0 23184 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0856_
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1644511149
transform 1 0 8004 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1644511149
transform 1 0 7360 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 12696 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0868_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0874_
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0880_
timestamp 1644511149
transform 1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0881_
timestamp 1644511149
transform 1 0 25668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0893_
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0899_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 46736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 25944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1644511149
transform 1 0 24932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 25484 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0912_
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0918_
timestamp 1644511149
transform 1 0 27784 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 28704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0924_
timestamp 1644511149
transform 1 0 28888 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 40756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0930_
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0936_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 46736 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0942_
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  _0943_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 25208 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 46736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 2760 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 33120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0949_
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 2944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 42596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0955_
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 25208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0961_
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 14352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0967_
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0975_
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _0978_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0980_
timestamp 1644511149
transform 1 0 25852 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0981_
timestamp 1644511149
transform 1 0 26864 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26680 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0985_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _0987_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0988_
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0989_
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1644511149
transform 1 0 44252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0994_
timestamp 1644511149
transform 1 0 45908 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _0995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1644511149
transform 1 0 44160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0997_
timestamp 1644511149
transform 1 0 44528 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0998_
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1644511149
transform 1 0 46092 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1000_
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _1001_
timestamp 1644511149
transform 1 0 43976 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1002_
timestamp 1644511149
transform 1 0 43332 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1644511149
transform 1 0 45356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1644511149
transform 1 0 45356 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1005_
timestamp 1644511149
transform 1 0 45264 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43608 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1007_
timestamp 1644511149
transform 1 0 45080 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__a21bo_1  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1009_
timestamp 1644511149
transform 1 0 43332 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1010_
timestamp 1644511149
transform 1 0 43792 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1011_
timestamp 1644511149
transform 1 0 27140 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1012_
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1013_
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1014_
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1018_
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform 1 0 30544 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1024_
timestamp 1644511149
transform 1 0 25944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 25392 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1030_
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 29624 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 25668 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 35604 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1036_
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 33488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 31096 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1042_
timestamp 1644511149
transform 1 0 18768 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 18400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 19320 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 19504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1048_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 20056 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1054_
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1055_
timestamp 1644511149
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1644511149
transform 1 0 16560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1057_
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1058_
timestamp 1644511149
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1059_
timestamp 1644511149
transform 1 0 12512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1060_
timestamp 1644511149
transform 1 0 12052 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1061_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1062_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1063_
timestamp 1644511149
transform 1 0 11776 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1065_
timestamp 1644511149
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1066_
timestamp 1644511149
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1067_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1068_
timestamp 1644511149
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1069_
timestamp 1644511149
transform 1 0 11684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1070_
timestamp 1644511149
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1071_
timestamp 1644511149
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1072_
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1644511149
transform 1 0 11408 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1074_
timestamp 1644511149
transform 1 0 11408 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1077_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1078_
timestamp 1644511149
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1079_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1080_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1081_
timestamp 1644511149
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1082_
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1083_
timestamp 1644511149
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1084_
timestamp 1644511149
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1085_
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1644511149
transform 1 0 21988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1644511149
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1088_
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1089_
timestamp 1644511149
transform 1 0 19320 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1092_
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1093_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1644511149
transform 1 0 29808 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1098_
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1099_
timestamp 1644511149
transform 1 0 22540 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1100_
timestamp 1644511149
transform 1 0 24472 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1101_
timestamp 1644511149
transform 1 0 29624 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1644511149
transform 1 0 24196 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1644511149
transform 1 0 33948 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1644511149
transform 1 0 34776 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1644511149
transform 1 0 32568 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1644511149
transform 1 0 23184 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1644511149
transform 1 0 19504 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1644511149
transform 1 0 16928 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1116_
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1117_
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1644511149
transform 1 0 17848 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1644511149
transform 1 0 18952 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1644511149
transform 1 0 19504 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1644511149
transform 1 0 16836 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1124_
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1125_
timestamp 1644511149
transform 1 0 17296 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1126_
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1644511149
transform 1 0 14904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1128_
timestamp 1644511149
transform 1 0 12788 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1129_
timestamp 1644511149
transform 1 0 12236 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1644511149
transform 1 0 11408 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1644511149
transform 1 0 11776 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1133_
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1644511149
transform 1 0 9108 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1135_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1644511149
transform 1 0 10580 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1644511149
transform 1 0 8004 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1644511149
transform 1 0 8832 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1139_
timestamp 1644511149
transform 1 0 9384 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1140_
timestamp 1644511149
transform 1 0 12236 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1644511149
transform 1 0 11684 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1143_
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1147_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1151_
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1644511149
transform 1 0 21068 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1155_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1156__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1157__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1158__83
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1159__84
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1160__85
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1161__86
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1162__87
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1163__88
timestamp 1644511149
transform 1 0 24564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1164__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__90
timestamp 1644511149
transform 1 0 25208 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__91
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__92
timestamp 1644511149
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__93
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__94
timestamp 1644511149
transform 1 0 2760 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__95
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__96
timestamp 1644511149
transform 1 0 42688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__98
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__99
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__101
timestamp 1644511149
transform 1 0 38088 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__102
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__103
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__104
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__105
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__106
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__108
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1184__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185__110
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1186__111
timestamp 1644511149
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1187__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1188__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1189__114
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1190__115
timestamp 1644511149
transform 1 0 24472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1191__116
timestamp 1644511149
transform 1 0 42688 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1192__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1193__118
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1194__119
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1195__120
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1196__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1197__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1198__123
timestamp 1644511149
transform 1 0 47472 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1199__124
timestamp 1644511149
transform 1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200__125
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1201__126
timestamp 1644511149
transform 1 0 20056 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1202__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1203__128
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1204__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1205__130
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1206__131
timestamp 1644511149
transform 1 0 1840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1207__132
timestamp 1644511149
transform 1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1208__133
timestamp 1644511149
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1209__134
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1210__135
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1212_
timestamp 1644511149
transform 1 0 27140 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1213_
timestamp 1644511149
transform 1 0 29624 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1214_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1215_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1216_
timestamp 1644511149
transform 1 0 40756 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1217_
timestamp 1644511149
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1218_
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1219_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1220_
timestamp 1644511149
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1224_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1225_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1226_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1227_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1228_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1229_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1231_
timestamp 1644511149
transform 1 0 1932 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1232_
timestamp 1644511149
transform 1 0 33028 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1233_
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1234_
timestamp 1644511149
transform 1 0 2024 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1235_
timestamp 1644511149
transform 1 0 42596 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1236_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1237_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1238_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1239_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1240_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1241_
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1242_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1243_
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1244_
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1245_
timestamp 1644511149
transform 1 0 14260 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1246_
timestamp 1644511149
transform 1 0 14260 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1247_
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1248_
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1249_
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1250_
timestamp 1644511149
transform 1 0 11684 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1251_
timestamp 1644511149
transform 1 0 11684 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1252_
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1253_
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1254_
timestamp 1644511149
transform 1 0 8004 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1255_
timestamp 1644511149
transform 1 0 7544 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1256_
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1257_
timestamp 1644511149
transform 1 0 8004 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1258_
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1259_
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1260_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1261_
timestamp 1644511149
transform 1 0 14168 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1262_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1263_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1264_
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1265_
timestamp 1644511149
transform 1 0 18952 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1266_
timestamp 1644511149
transform 1 0 15364 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1267_
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1268_
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1269_
timestamp 1644511149
transform 1 0 19504 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1270_
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1271_
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1272_
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1273_
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1274_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1275_
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1276_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 25116 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22080 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 2944 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 47288 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 47932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1644511149
transform 1 0 47288 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 46184 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 2024 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1644511149
transform 1 0 47840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1644511149
transform 1 0 9108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1644511149
transform 1 0 43792 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 11684 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 46184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 47288 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 39100 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 24380 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44804 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 28244 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 29532 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 15272 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1932 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45448 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35972 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 45816 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 43240 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 28520 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
