magic
tech sky130A
magscale 1 2
timestamp 1654519615
<< viali >>
rect 13369 47209 13403 47243
rect 21833 47141 21867 47175
rect 28641 47141 28675 47175
rect 43867 47141 43901 47175
rect 47961 47141 47995 47175
rect 6653 47073 6687 47107
rect 30757 47073 30791 47107
rect 39865 47073 39899 47107
rect 43637 47073 43671 47107
rect 47041 47073 47075 47107
rect 1777 47005 1811 47039
rect 3801 47005 3835 47039
rect 4813 47005 4847 47039
rect 6377 47005 6411 47039
rect 7389 47005 7423 47039
rect 9413 47005 9447 47039
rect 11621 47005 11655 47039
rect 12357 47005 12391 47039
rect 13093 47005 13127 47039
rect 14105 47005 14139 47039
rect 14381 47005 14415 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 21005 47005 21039 47039
rect 22017 47005 22051 47039
rect 24777 47005 24811 47039
rect 25421 47005 25455 47039
rect 28457 47005 28491 47039
rect 30021 47005 30055 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 40141 47005 40175 47039
rect 41889 47005 41923 47039
rect 42993 47005 43027 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2053 46937 2087 46971
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 7573 46937 7607 46971
rect 9597 46937 9631 46971
rect 11805 46937 11839 46971
rect 12541 46937 12575 46971
rect 19717 46937 19751 46971
rect 20085 46937 20119 46971
rect 30205 46937 30239 46971
rect 43177 46937 43211 46971
rect 45385 46937 45419 46971
rect 2881 46869 2915 46903
rect 4905 46869 4939 46903
rect 1869 46597 1903 46631
rect 24593 46529 24627 46563
rect 38117 46529 38151 46563
rect 47961 46529 47995 46563
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 12173 46461 12207 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19257 46461 19291 46495
rect 19441 46461 19475 46495
rect 20453 46461 20487 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 34437 46461 34471 46495
rect 34621 46461 34655 46495
rect 34897 46461 34931 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46765 46461 46799 46495
rect 2145 46325 2179 46359
rect 2881 46325 2915 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 12081 46121 12115 46155
rect 13553 46121 13587 46155
rect 14197 46121 14231 46155
rect 18613 46121 18647 46155
rect 19441 46121 19475 46155
rect 24685 46121 24719 46155
rect 32045 46121 32079 46155
rect 33609 46121 33643 46155
rect 34805 46121 34839 46155
rect 38301 46121 38335 46155
rect 43821 46121 43855 46155
rect 1409 45985 1443 46019
rect 2789 45985 2823 46019
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41245 45985 41279 46019
rect 41981 45985 42015 46019
rect 44465 45985 44499 46019
rect 46305 45985 46339 46019
rect 47041 45985 47075 46019
rect 11989 45917 12023 45951
rect 14105 45917 14139 45951
rect 18521 45917 18555 45951
rect 24593 45917 24627 45951
rect 31953 45917 31987 45951
rect 34713 45917 34747 45951
rect 38209 45917 38243 45951
rect 45661 45917 45695 45951
rect 1593 45849 1627 45883
rect 20913 45849 20947 45883
rect 25421 45849 25455 45883
rect 41429 45849 41463 45883
rect 46489 45849 46523 45883
rect 45753 45781 45787 45815
rect 2237 45577 2271 45611
rect 20913 45577 20947 45611
rect 41797 45577 41831 45611
rect 25421 45509 25455 45543
rect 41153 45509 41187 45543
rect 47961 45509 47995 45543
rect 2145 45441 2179 45475
rect 20821 45441 20855 45475
rect 25329 45441 25363 45475
rect 41061 45441 41095 45475
rect 41705 45441 41739 45475
rect 42717 45441 42751 45475
rect 42901 45373 42935 45407
rect 44097 45373 44131 45407
rect 45017 45373 45051 45407
rect 45201 45373 45235 45407
rect 45753 45373 45787 45407
rect 48053 45237 48087 45271
rect 42901 45033 42935 45067
rect 44465 45033 44499 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 42809 44829 42843 44863
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 46397 44489 46431 44523
rect 47685 44489 47719 44523
rect 44925 44353 44959 44387
rect 45661 44353 45695 44387
rect 46305 44353 46339 44387
rect 47593 44353 47627 44387
rect 45753 44149 45787 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 47685 43401 47719 43435
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 47593 43265 47627 43299
rect 1593 43197 1627 43231
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 48145 41497 48179 41531
rect 2145 41225 2179 41259
rect 46857 41225 46891 41259
rect 2053 41089 2087 41123
rect 46765 41089 46799 41123
rect 47961 41089 47995 41123
rect 48145 40953 48179 40987
rect 47685 40681 47719 40715
rect 26893 40545 26927 40579
rect 26709 40477 26743 40511
rect 47041 40477 47075 40511
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 26249 40341 26283 40375
rect 26617 40341 26651 40375
rect 25881 40137 25915 40171
rect 19901 40001 19935 40035
rect 47593 40001 47627 40035
rect 24133 39933 24167 39967
rect 24409 39933 24443 39967
rect 19993 39797 20027 39831
rect 47685 39797 47719 39831
rect 22937 39593 22971 39627
rect 25145 39593 25179 39627
rect 26617 39593 26651 39627
rect 26341 39457 26375 39491
rect 46305 39457 46339 39491
rect 46489 39457 46523 39491
rect 48145 39457 48179 39491
rect 19257 39389 19291 39423
rect 22845 39389 22879 39423
rect 25329 39389 25363 39423
rect 26249 39389 26283 39423
rect 19533 39321 19567 39355
rect 21005 39253 21039 39287
rect 18981 39049 19015 39083
rect 19625 39049 19659 39083
rect 19993 39049 20027 39083
rect 26341 38981 26375 39015
rect 19165 38913 19199 38947
rect 21925 38913 21959 38947
rect 23213 38913 23247 38947
rect 26249 38913 26283 38947
rect 29929 38913 29963 38947
rect 46121 38913 46155 38947
rect 47869 38913 47903 38947
rect 20085 38845 20119 38879
rect 20177 38845 20211 38879
rect 23857 38845 23891 38879
rect 24133 38845 24167 38879
rect 26985 38845 27019 38879
rect 27261 38845 27295 38879
rect 28733 38845 28767 38879
rect 30021 38845 30055 38879
rect 30113 38845 30147 38879
rect 22109 38709 22143 38743
rect 23305 38709 23339 38743
rect 25605 38709 25639 38743
rect 29561 38709 29595 38743
rect 46213 38709 46247 38743
rect 48053 38709 48087 38743
rect 20177 38505 20211 38539
rect 24409 38505 24443 38539
rect 25145 38505 25179 38539
rect 25973 38505 26007 38539
rect 31309 38505 31343 38539
rect 20729 38369 20763 38403
rect 26157 38369 26191 38403
rect 27537 38369 27571 38403
rect 29561 38369 29595 38403
rect 46397 38369 46431 38403
rect 48053 38369 48087 38403
rect 19257 38301 19291 38335
rect 20545 38301 20579 38335
rect 22017 38301 22051 38335
rect 24593 38301 24627 38335
rect 25053 38301 25087 38335
rect 26249 38301 26283 38335
rect 27261 38301 27295 38335
rect 29009 38301 29043 38335
rect 46213 38301 46247 38335
rect 22293 38233 22327 38267
rect 25973 38233 26007 38267
rect 29837 38233 29871 38267
rect 19349 38165 19383 38199
rect 20637 38165 20671 38199
rect 23765 38165 23799 38199
rect 26433 38165 26467 38199
rect 26893 38165 26927 38199
rect 27353 38165 27387 38199
rect 28825 38165 28859 38199
rect 22385 37961 22419 37995
rect 24961 37961 24995 37995
rect 26985 37961 27019 37995
rect 29837 37961 29871 37995
rect 31125 37961 31159 37995
rect 20177 37825 20211 37859
rect 22569 37825 22603 37859
rect 23029 37825 23063 37859
rect 25329 37825 25363 37859
rect 27169 37825 27203 37859
rect 30205 37825 30239 37859
rect 31033 37825 31067 37859
rect 33149 37825 33183 37859
rect 46673 37825 46707 37859
rect 17601 37757 17635 37791
rect 17877 37757 17911 37791
rect 20085 37757 20119 37791
rect 25421 37757 25455 37791
rect 25605 37757 25639 37791
rect 30297 37757 30331 37791
rect 30481 37757 30515 37791
rect 20545 37689 20579 37723
rect 29469 37689 29503 37723
rect 19349 37621 19383 37655
rect 23213 37621 23247 37655
rect 32965 37621 32999 37655
rect 46765 37621 46799 37655
rect 47777 37621 47811 37655
rect 18245 37417 18279 37451
rect 23121 37417 23155 37451
rect 27353 37417 27387 37451
rect 30021 37417 30055 37451
rect 26893 37349 26927 37383
rect 19901 37281 19935 37315
rect 23673 37281 23707 37315
rect 26617 37281 26651 37315
rect 27905 37281 27939 37315
rect 29653 37281 29687 37315
rect 32689 37281 32723 37315
rect 35265 37281 35299 37315
rect 46489 37281 46523 37315
rect 48145 37281 48179 37315
rect 2053 37213 2087 37247
rect 18429 37213 18463 37247
rect 19625 37213 19659 37247
rect 23489 37213 23523 37247
rect 24685 37213 24719 37247
rect 24869 37213 24903 37247
rect 26525 37213 26559 37247
rect 27813 37213 27847 37247
rect 29745 37213 29779 37247
rect 32413 37213 32447 37247
rect 35081 37213 35115 37247
rect 46305 37213 46339 37247
rect 19257 37077 19291 37111
rect 19717 37077 19751 37111
rect 23581 37077 23615 37111
rect 24777 37077 24811 37111
rect 27721 37077 27755 37111
rect 34161 37077 34195 37111
rect 34713 37077 34747 37111
rect 35173 37077 35207 37111
rect 19901 36873 19935 36907
rect 23489 36873 23523 36907
rect 23949 36873 23983 36907
rect 33149 36873 33183 36907
rect 33609 36873 33643 36907
rect 34897 36873 34931 36907
rect 24961 36805 24995 36839
rect 25145 36805 25179 36839
rect 1777 36737 1811 36771
rect 19257 36737 19291 36771
rect 19441 36737 19475 36771
rect 20269 36737 20303 36771
rect 22109 36737 22143 36771
rect 23857 36737 23891 36771
rect 24777 36737 24811 36771
rect 25697 36737 25731 36771
rect 25881 36737 25915 36771
rect 26065 36737 26099 36771
rect 26249 36737 26283 36771
rect 27169 36737 27203 36771
rect 27353 36737 27387 36771
rect 29193 36737 29227 36771
rect 29377 36737 29411 36771
rect 33517 36737 33551 36771
rect 34529 36737 34563 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 19349 36669 19383 36703
rect 20361 36669 20395 36703
rect 20545 36669 20579 36703
rect 24041 36669 24075 36703
rect 26433 36669 26467 36703
rect 27445 36669 27479 36703
rect 29837 36669 29871 36703
rect 30113 36669 30147 36703
rect 31585 36669 31619 36703
rect 33701 36669 33735 36703
rect 34621 36669 34655 36703
rect 22201 36533 22235 36567
rect 26985 36533 27019 36567
rect 29193 36533 29227 36567
rect 2237 36329 2271 36363
rect 24777 36329 24811 36363
rect 25789 36329 25823 36363
rect 28917 36329 28951 36363
rect 30297 36329 30331 36363
rect 31033 36329 31067 36363
rect 33609 36329 33643 36363
rect 19441 36261 19475 36295
rect 20637 36261 20671 36295
rect 26157 36261 26191 36295
rect 19533 36193 19567 36227
rect 20729 36193 20763 36227
rect 21465 36193 21499 36227
rect 29929 36193 29963 36227
rect 2145 36125 2179 36159
rect 18521 36125 18555 36159
rect 19257 36125 19291 36159
rect 19349 36125 19383 36159
rect 20453 36125 20487 36159
rect 21189 36125 21223 36159
rect 24685 36125 24719 36159
rect 24869 36125 24903 36159
rect 25973 36125 26007 36159
rect 26065 36125 26099 36159
rect 26249 36125 26283 36159
rect 27169 36125 27203 36159
rect 28733 36125 28767 36159
rect 29009 36125 29043 36159
rect 29561 36125 29595 36159
rect 29745 36125 29779 36159
rect 29837 36125 29871 36159
rect 30113 36125 30147 36159
rect 30941 36125 30975 36159
rect 33517 36125 33551 36159
rect 26801 36057 26835 36091
rect 26985 36057 27019 36091
rect 18613 35989 18647 36023
rect 20269 35989 20303 36023
rect 22937 35989 22971 36023
rect 28549 35989 28583 36023
rect 22569 35785 22603 35819
rect 30481 35785 30515 35819
rect 31309 35785 31343 35819
rect 17785 35717 17819 35751
rect 30113 35717 30147 35751
rect 1593 35649 1627 35683
rect 17969 35649 18003 35683
rect 18613 35649 18647 35683
rect 18797 35649 18831 35683
rect 19349 35649 19383 35683
rect 19441 35649 19475 35683
rect 20177 35649 20211 35683
rect 20361 35649 20395 35683
rect 21833 35649 21867 35683
rect 22017 35649 22051 35683
rect 22385 35649 22419 35683
rect 30297 35649 30331 35683
rect 30941 35649 30975 35683
rect 48145 35649 48179 35683
rect 22109 35581 22143 35615
rect 22201 35581 22235 35615
rect 28825 35581 28859 35615
rect 29101 35581 29135 35615
rect 31033 35581 31067 35615
rect 18705 35513 18739 35547
rect 19717 35513 19751 35547
rect 1409 35445 1443 35479
rect 18153 35445 18187 35479
rect 19349 35445 19383 35479
rect 20361 35445 20395 35479
rect 20545 35445 20579 35479
rect 30941 35445 30975 35479
rect 47961 35445 47995 35479
rect 20637 35241 20671 35275
rect 22569 35241 22603 35275
rect 29009 35241 29043 35275
rect 33885 35241 33919 35275
rect 17693 35105 17727 35139
rect 19349 35105 19383 35139
rect 20729 35105 20763 35139
rect 28181 35105 28215 35139
rect 31309 35105 31343 35139
rect 33977 35105 34011 35139
rect 35357 35105 35391 35139
rect 16681 35037 16715 35071
rect 16957 35037 16991 35071
rect 17417 35037 17451 35071
rect 17601 35037 17635 35071
rect 17785 35037 17819 35071
rect 17969 35037 18003 35071
rect 19625 35037 19659 35071
rect 20637 35037 20671 35071
rect 23581 35037 23615 35071
rect 28825 35037 28859 35071
rect 30021 35037 30055 35071
rect 30205 35037 30239 35071
rect 30297 35037 30331 35071
rect 30389 35037 30423 35071
rect 30573 35037 30607 35071
rect 33701 35037 33735 35071
rect 35081 35037 35115 35071
rect 48145 35037 48179 35071
rect 16865 34969 16899 35003
rect 22477 34969 22511 35003
rect 27997 34969 28031 35003
rect 28641 34969 28675 35003
rect 30757 34969 30791 35003
rect 31585 34969 31619 35003
rect 16957 34901 16991 34935
rect 18153 34901 18187 34935
rect 21005 34901 21039 34935
rect 23673 34901 23707 34935
rect 33057 34901 33091 34935
rect 33517 34901 33551 34935
rect 34713 34901 34747 34935
rect 35173 34901 35207 34935
rect 47961 34901 47995 34935
rect 19257 34697 19291 34731
rect 28457 34697 28491 34731
rect 30297 34697 30331 34731
rect 31401 34697 31435 34731
rect 32597 34697 32631 34731
rect 34253 34697 34287 34731
rect 35081 34697 35115 34731
rect 35633 34697 35667 34731
rect 17785 34629 17819 34663
rect 21925 34629 21959 34663
rect 26985 34629 27019 34663
rect 33793 34629 33827 34663
rect 17509 34561 17543 34595
rect 20453 34561 20487 34595
rect 22569 34561 22603 34595
rect 24777 34561 24811 34595
rect 25053 34561 25087 34595
rect 26157 34561 26191 34595
rect 27169 34561 27203 34595
rect 28273 34561 28307 34595
rect 29101 34561 29135 34595
rect 29745 34561 29779 34595
rect 30941 34561 30975 34595
rect 31585 34561 31619 34595
rect 32505 34561 32539 34595
rect 34069 34561 34103 34595
rect 34713 34561 34747 34595
rect 34897 34561 34931 34595
rect 35541 34561 35575 34595
rect 35725 34561 35759 34595
rect 47777 34561 47811 34595
rect 20177 34493 20211 34527
rect 22845 34493 22879 34527
rect 25145 34493 25179 34527
rect 26249 34493 26283 34527
rect 29285 34493 29319 34527
rect 30021 34493 30055 34527
rect 33977 34493 34011 34527
rect 22109 34425 22143 34459
rect 24869 34425 24903 34459
rect 24317 34357 24351 34391
rect 24961 34357 24995 34391
rect 27353 34357 27387 34391
rect 30113 34357 30147 34391
rect 30757 34357 30791 34391
rect 33977 34357 34011 34391
rect 47593 34357 47627 34391
rect 20545 34153 20579 34187
rect 21373 34153 21407 34187
rect 23489 34153 23523 34187
rect 24593 34153 24627 34187
rect 27353 34153 27387 34187
rect 27813 34153 27847 34187
rect 34805 34153 34839 34187
rect 20453 34017 20487 34051
rect 23121 34017 23155 34051
rect 25145 34017 25179 34051
rect 27537 34017 27571 34051
rect 28641 34017 28675 34051
rect 30205 34017 30239 34051
rect 33977 34017 34011 34051
rect 47133 34017 47167 34051
rect 47593 34017 47627 34051
rect 1593 33949 1627 33983
rect 20545 33949 20579 33983
rect 21281 33949 21315 33983
rect 21465 33949 21499 33983
rect 22753 33949 22787 33983
rect 22937 33949 22971 33983
rect 23029 33949 23063 33983
rect 23305 33949 23339 33983
rect 24501 33949 24535 33983
rect 27629 33949 27663 33983
rect 28825 33949 28859 33983
rect 29929 33949 29963 33983
rect 30113 33949 30147 33983
rect 30297 33949 30331 33983
rect 30481 33949 30515 33983
rect 32965 33949 32999 33983
rect 33885 33949 33919 33983
rect 34713 33949 34747 33983
rect 34897 33949 34931 33983
rect 20269 33881 20303 33915
rect 25421 33881 25455 33915
rect 27353 33881 27387 33915
rect 33793 33881 33827 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 20729 33813 20763 33847
rect 26893 33813 26927 33847
rect 29009 33813 29043 33847
rect 30665 33813 30699 33847
rect 32781 33813 32815 33847
rect 33425 33813 33459 33847
rect 23489 33609 23523 33643
rect 30021 33609 30055 33643
rect 35173 33609 35207 33643
rect 48053 33609 48087 33643
rect 22845 33541 22879 33575
rect 27169 33541 27203 33575
rect 28641 33541 28675 33575
rect 28825 33541 28859 33575
rect 29009 33541 29043 33575
rect 33701 33541 33735 33575
rect 20453 33473 20487 33507
rect 20545 33473 20579 33507
rect 23673 33473 23707 33507
rect 23765 33473 23799 33507
rect 23949 33473 23983 33507
rect 24041 33473 24075 33507
rect 24685 33473 24719 33507
rect 27445 33473 27479 33507
rect 29469 33473 29503 33507
rect 32321 33473 32355 33507
rect 46765 33473 46799 33507
rect 47593 33473 47627 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 20729 33405 20763 33439
rect 27353 33405 27387 33439
rect 29745 33405 29779 33439
rect 33425 33405 33459 33439
rect 27629 33337 27663 33371
rect 20085 33269 20119 33303
rect 22937 33269 22971 33303
rect 25973 33269 26007 33303
rect 27169 33269 27203 33303
rect 29561 33269 29595 33303
rect 32413 33269 32447 33303
rect 46949 33269 46983 33303
rect 47869 33269 47903 33303
rect 1961 33065 1995 33099
rect 21005 33065 21039 33099
rect 23673 33065 23707 33099
rect 25605 33065 25639 33099
rect 26065 33065 26099 33099
rect 26525 33065 26559 33099
rect 27629 33065 27663 33099
rect 28641 33065 28675 33099
rect 32781 33065 32815 33099
rect 34805 33065 34839 33099
rect 21925 32997 21959 33031
rect 2329 32929 2363 32963
rect 19809 32929 19843 32963
rect 19993 32929 20027 32963
rect 20821 32929 20855 32963
rect 25237 32929 25271 32963
rect 25881 32929 25915 32963
rect 26157 32929 26191 32963
rect 29837 32929 29871 32963
rect 31033 32929 31067 32963
rect 31309 32929 31343 32963
rect 1869 32861 1903 32895
rect 2973 32861 3007 32895
rect 18705 32861 18739 32895
rect 19717 32861 19751 32895
rect 20729 32861 20763 32895
rect 21557 32861 21591 32895
rect 23673 32861 23707 32895
rect 23857 32861 23891 32895
rect 24869 32861 24903 32895
rect 25053 32861 25087 32895
rect 25145 32861 25179 32895
rect 25421 32861 25455 32895
rect 26341 32861 26375 32895
rect 27445 32861 27479 32895
rect 28457 32861 28491 32895
rect 28641 32861 28675 32895
rect 29561 32861 29595 32895
rect 29653 32861 29687 32895
rect 34713 32861 34747 32895
rect 45845 32861 45879 32895
rect 46305 32861 46339 32895
rect 21741 32793 21775 32827
rect 26065 32793 26099 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 2789 32725 2823 32759
rect 18521 32725 18555 32759
rect 19349 32725 19383 32759
rect 28825 32725 28859 32759
rect 29837 32725 29871 32759
rect 25053 32521 25087 32555
rect 26341 32521 26375 32555
rect 46949 32521 46983 32555
rect 2237 32453 2271 32487
rect 18153 32453 18187 32487
rect 2053 32385 2087 32419
rect 20269 32385 20303 32419
rect 20545 32385 20579 32419
rect 21005 32385 21039 32419
rect 21189 32385 21223 32419
rect 24685 32385 24719 32419
rect 25513 32385 25547 32419
rect 25697 32385 25731 32419
rect 26249 32385 26283 32419
rect 27445 32385 27479 32419
rect 28365 32385 28399 32419
rect 28641 32385 28675 32419
rect 29745 32385 29779 32419
rect 31033 32385 31067 32419
rect 32137 32385 32171 32419
rect 46857 32385 46891 32419
rect 47961 32385 47995 32419
rect 3893 32317 3927 32351
rect 17877 32317 17911 32351
rect 19625 32317 19659 32351
rect 24777 32317 24811 32351
rect 28549 32317 28583 32351
rect 29837 32317 29871 32351
rect 29929 32317 29963 32351
rect 20453 32249 20487 32283
rect 48145 32249 48179 32283
rect 1593 32181 1627 32215
rect 20085 32181 20119 32215
rect 21005 32181 21039 32215
rect 24869 32181 24903 32215
rect 25513 32181 25547 32215
rect 27629 32181 27663 32215
rect 28549 32181 28583 32215
rect 28825 32181 28859 32215
rect 29377 32181 29411 32215
rect 31125 32181 31159 32215
rect 32321 32181 32355 32215
rect 19349 31977 19383 32011
rect 20453 31977 20487 32011
rect 27261 31977 27295 32011
rect 28825 31977 28859 32011
rect 31861 31977 31895 32011
rect 20821 31909 20855 31943
rect 23765 31909 23799 31943
rect 26525 31909 26559 31943
rect 32505 31909 32539 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 3801 31841 3835 31875
rect 3985 31841 4019 31875
rect 4629 31841 4663 31875
rect 12449 31841 12483 31875
rect 14841 31841 14875 31875
rect 15301 31841 15335 31875
rect 17969 31841 18003 31875
rect 24133 31841 24167 31875
rect 25697 31841 25731 31875
rect 35265 31841 35299 31875
rect 46765 31841 46799 31875
rect 47593 31841 47627 31875
rect 11713 31773 11747 31807
rect 17601 31773 17635 31807
rect 17785 31773 17819 31807
rect 17877 31773 17911 31807
rect 18153 31773 18187 31807
rect 19257 31773 19291 31807
rect 20453 31773 20487 31807
rect 20637 31773 20671 31807
rect 21373 31773 21407 31807
rect 21557 31773 21591 31807
rect 22017 31773 22051 31807
rect 24041 31773 24075 31807
rect 24225 31773 24259 31807
rect 24869 31773 24903 31807
rect 25513 31773 25547 31807
rect 26341 31773 26375 31807
rect 27169 31773 27203 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 28825 31773 28859 31807
rect 30113 31773 30147 31807
rect 32321 31773 32355 31807
rect 1593 31705 1627 31739
rect 11897 31705 11931 31739
rect 15025 31705 15059 31739
rect 22293 31705 22327 31739
rect 30389 31705 30423 31739
rect 35173 31705 35207 31739
rect 46857 31705 46891 31739
rect 18337 31637 18371 31671
rect 25145 31637 25179 31671
rect 25605 31637 25639 31671
rect 29009 31637 29043 31671
rect 34713 31637 34747 31671
rect 35081 31637 35115 31671
rect 2237 31433 2271 31467
rect 12909 31433 12943 31467
rect 14841 31433 14875 31467
rect 19073 31433 19107 31467
rect 22661 31433 22695 31467
rect 23305 31433 23339 31467
rect 23765 31433 23799 31467
rect 27629 31433 27663 31467
rect 28825 31433 28859 31467
rect 29377 31433 29411 31467
rect 30573 31433 30607 31467
rect 31493 31433 31527 31467
rect 19625 31365 19659 31399
rect 35817 31365 35851 31399
rect 2145 31297 2179 31331
rect 12817 31297 12851 31331
rect 14749 31297 14783 31331
rect 19533 31297 19567 31331
rect 22845 31297 22879 31331
rect 23673 31297 23707 31331
rect 24961 31297 24995 31331
rect 25789 31297 25823 31331
rect 27445 31297 27479 31331
rect 28641 31297 28675 31331
rect 29745 31297 29779 31331
rect 30757 31297 30791 31331
rect 31401 31297 31435 31331
rect 32321 31297 32355 31331
rect 35725 31297 35759 31331
rect 17325 31229 17359 31263
rect 17601 31229 17635 31263
rect 23949 31229 23983 31263
rect 25053 31229 25087 31263
rect 25329 31229 25363 31263
rect 29837 31229 29871 31263
rect 30021 31229 30055 31263
rect 32137 31229 32171 31263
rect 33517 31229 33551 31263
rect 33793 31229 33827 31263
rect 25881 31093 25915 31127
rect 26249 31093 26283 31127
rect 32505 31093 32539 31127
rect 35265 31093 35299 31127
rect 23489 30889 23523 30923
rect 26985 30889 27019 30923
rect 29653 30889 29687 30923
rect 31677 30889 31711 30923
rect 33885 30889 33919 30923
rect 34713 30889 34747 30923
rect 17877 30753 17911 30787
rect 35357 30753 35391 30787
rect 12541 30685 12575 30719
rect 13001 30685 13035 30719
rect 14749 30685 14783 30719
rect 16313 30685 16347 30719
rect 19809 30685 19843 30719
rect 20269 30685 20303 30719
rect 23397 30685 23431 30719
rect 25789 30685 25823 30719
rect 25937 30685 25971 30719
rect 26157 30685 26191 30719
rect 26295 30685 26329 30719
rect 27169 30685 27203 30719
rect 27445 30685 27479 30719
rect 28365 30685 28399 30719
rect 29561 30685 29595 30719
rect 29745 30685 29779 30719
rect 31493 30685 31527 30719
rect 34069 30685 34103 30719
rect 35081 30685 35115 30719
rect 15025 30617 15059 30651
rect 16497 30617 16531 30651
rect 26065 30617 26099 30651
rect 28549 30617 28583 30651
rect 32321 30617 32355 30651
rect 12357 30549 12391 30583
rect 13093 30549 13127 30583
rect 19625 30549 19659 30583
rect 20361 30549 20395 30583
rect 26433 30549 26467 30583
rect 27353 30549 27387 30583
rect 32413 30549 32447 30583
rect 35173 30549 35207 30583
rect 13921 30345 13955 30379
rect 25145 30345 25179 30379
rect 34713 30345 34747 30379
rect 12449 30277 12483 30311
rect 19257 30277 19291 30311
rect 27445 30277 27479 30311
rect 27629 30277 27663 30311
rect 28273 30277 28307 30311
rect 29377 30277 29411 30311
rect 9781 30209 9815 30243
rect 10241 30209 10275 30243
rect 14841 30209 14875 30243
rect 15669 30209 15703 30243
rect 22293 30209 22327 30243
rect 28089 30209 28123 30243
rect 28365 30209 28399 30243
rect 29193 30209 29227 30243
rect 34529 30209 34563 30243
rect 34713 30209 34747 30243
rect 12173 30141 12207 30175
rect 14933 30141 14967 30175
rect 16681 30141 16715 30175
rect 16865 30141 16899 30175
rect 17601 30141 17635 30175
rect 18981 30141 19015 30175
rect 23397 30141 23431 30175
rect 23673 30141 23707 30175
rect 28089 30073 28123 30107
rect 9597 30005 9631 30039
rect 10333 30005 10367 30039
rect 15209 30005 15243 30039
rect 15761 30005 15795 30039
rect 20729 30005 20763 30039
rect 22385 30005 22419 30039
rect 13001 29801 13035 29835
rect 16865 29801 16899 29835
rect 17509 29801 17543 29835
rect 20453 29801 20487 29835
rect 24501 29801 24535 29835
rect 25973 29801 26007 29835
rect 27077 29801 27111 29835
rect 28549 29801 28583 29835
rect 30205 29801 30239 29835
rect 30941 29801 30975 29835
rect 14197 29733 14231 29767
rect 9689 29665 9723 29699
rect 11161 29665 11195 29699
rect 12081 29665 12115 29699
rect 15117 29665 15151 29699
rect 15393 29665 15427 29699
rect 21097 29665 21131 29699
rect 21833 29665 21867 29699
rect 22753 29665 22787 29699
rect 33241 29665 33275 29699
rect 9413 29597 9447 29631
rect 12173 29597 12207 29631
rect 12541 29597 12575 29631
rect 13231 29597 13265 29631
rect 13461 29597 13495 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 17417 29597 17451 29631
rect 19257 29597 19291 29631
rect 21925 29597 21959 29631
rect 22017 29597 22051 29631
rect 22109 29597 22143 29631
rect 22661 29597 22695 29631
rect 22845 29597 22879 29631
rect 23397 29597 23431 29631
rect 24409 29597 24443 29631
rect 26203 29597 26237 29631
rect 26338 29597 26372 29631
rect 26438 29597 26472 29631
rect 26617 29597 26651 29631
rect 27077 29597 27111 29631
rect 27261 29597 27295 29631
rect 29561 29597 29595 29631
rect 29709 29597 29743 29631
rect 30026 29597 30060 29631
rect 30757 29597 30791 29631
rect 48145 29597 48179 29631
rect 13369 29529 13403 29563
rect 14105 29529 14139 29563
rect 28457 29529 28491 29563
rect 29837 29529 29871 29563
rect 29929 29529 29963 29563
rect 33149 29529 33183 29563
rect 11897 29461 11931 29495
rect 12357 29461 12391 29495
rect 12449 29461 12483 29495
rect 19441 29461 19475 29495
rect 20177 29461 20211 29495
rect 20821 29461 20855 29495
rect 20913 29461 20947 29495
rect 21649 29461 21683 29495
rect 23489 29461 23523 29495
rect 27445 29461 27479 29495
rect 32689 29461 32723 29495
rect 33057 29461 33091 29495
rect 47961 29461 47995 29495
rect 9321 29257 9355 29291
rect 10517 29257 10551 29291
rect 12265 29257 12299 29291
rect 13093 29257 13127 29291
rect 16773 29257 16807 29291
rect 21833 29257 21867 29291
rect 22937 29257 22971 29291
rect 32689 29257 32723 29291
rect 33149 29257 33183 29291
rect 34437 29257 34471 29291
rect 35173 29257 35207 29291
rect 12725 29189 12759 29223
rect 13001 29189 13035 29223
rect 14473 29189 14507 29223
rect 16129 29189 16163 29223
rect 20913 29189 20947 29223
rect 21097 29189 21131 29223
rect 30021 29189 30055 29223
rect 9229 29121 9263 29155
rect 11897 29121 11931 29155
rect 12081 29121 12115 29155
rect 12909 29121 12943 29155
rect 16681 29121 16715 29155
rect 19073 29121 19107 29155
rect 22017 29121 22051 29155
rect 22753 29121 22787 29155
rect 27077 29121 27111 29155
rect 27353 29121 27387 29155
rect 27813 29121 27847 29155
rect 28089 29121 28123 29155
rect 29101 29121 29135 29155
rect 29745 29121 29779 29155
rect 33057 29121 33091 29155
rect 34069 29121 34103 29155
rect 34897 29121 34931 29155
rect 10057 29053 10091 29087
rect 14289 29053 14323 29087
rect 22293 29053 22327 29087
rect 28457 29053 28491 29087
rect 28917 29053 28951 29087
rect 31493 29053 31527 29087
rect 33241 29053 33275 29087
rect 34161 29053 34195 29087
rect 34989 29053 35023 29087
rect 35173 29053 35207 29087
rect 10425 28985 10459 29019
rect 13277 28985 13311 29019
rect 19257 28985 19291 29019
rect 22201 28985 22235 29019
rect 29285 28985 29319 29019
rect 21281 28917 21315 28951
rect 12541 28713 12575 28747
rect 18245 28713 18279 28747
rect 18613 28713 18647 28747
rect 19809 28713 19843 28747
rect 26433 28713 26467 28747
rect 30113 28713 30147 28747
rect 30941 28713 30975 28747
rect 34161 28713 34195 28747
rect 34713 28713 34747 28747
rect 35173 28713 35207 28747
rect 21465 28645 21499 28679
rect 9781 28577 9815 28611
rect 15945 28577 15979 28611
rect 16589 28577 16623 28611
rect 18705 28577 18739 28611
rect 23213 28577 23247 28611
rect 26525 28577 26559 28611
rect 28917 28577 28951 28611
rect 29653 28577 29687 28611
rect 32413 28577 32447 28611
rect 34805 28577 34839 28611
rect 9321 28509 9355 28543
rect 12541 28509 12575 28543
rect 18429 28509 18463 28543
rect 20361 28509 20395 28543
rect 21373 28509 21407 28543
rect 21557 28509 21591 28543
rect 21649 28509 21683 28543
rect 22845 28509 22879 28543
rect 23033 28511 23067 28545
rect 23130 28509 23164 28543
rect 23397 28509 23431 28543
rect 24409 28509 24443 28543
rect 26065 28509 26099 28543
rect 27445 28509 27479 28543
rect 27721 28509 27755 28543
rect 27997 28509 28031 28543
rect 28181 28509 28215 28543
rect 28825 28509 28859 28543
rect 29009 28509 29043 28543
rect 29745 28509 29779 28543
rect 30849 28509 30883 28543
rect 31769 28509 31803 28543
rect 34989 28509 35023 28543
rect 47685 28509 47719 28543
rect 9505 28441 9539 28475
rect 14565 28441 14599 28475
rect 16129 28441 16163 28475
rect 19717 28441 19751 28475
rect 26157 28441 26191 28475
rect 32689 28441 32723 28475
rect 34713 28441 34747 28475
rect 14657 28373 14691 28407
rect 20453 28373 20487 28407
rect 21189 28373 21223 28407
rect 23581 28373 23615 28407
rect 24501 28373 24535 28407
rect 25789 28373 25823 28407
rect 26249 28373 26283 28407
rect 27537 28373 27571 28407
rect 31861 28373 31895 28407
rect 10057 28169 10091 28203
rect 16037 28169 16071 28203
rect 16773 28169 16807 28203
rect 17969 28169 18003 28203
rect 24409 28169 24443 28203
rect 28273 28169 28307 28203
rect 32597 28169 32631 28203
rect 21833 28101 21867 28135
rect 22201 28101 22235 28135
rect 22937 28101 22971 28135
rect 24869 28101 24903 28135
rect 25513 28101 25547 28135
rect 8217 28033 8251 28067
rect 9321 28033 9355 28067
rect 9965 28033 9999 28067
rect 11897 28033 11931 28067
rect 12909 28033 12943 28067
rect 13461 28033 13495 28067
rect 15945 28033 15979 28067
rect 16681 28033 16715 28067
rect 18245 28033 18279 28067
rect 18429 28033 18463 28067
rect 19257 28033 19291 28067
rect 22017 28033 22051 28067
rect 27445 28033 27479 28067
rect 27537 28033 27571 28067
rect 27629 28033 27663 28067
rect 27813 28033 27847 28067
rect 28457 28033 28491 28067
rect 28733 28033 28767 28067
rect 32781 28033 32815 28067
rect 47593 28033 47627 28067
rect 11989 27965 12023 27999
rect 17877 27965 17911 27999
rect 18153 27965 18187 27999
rect 19533 27965 19567 27999
rect 21005 27965 21039 27999
rect 22661 27965 22695 27999
rect 25605 27965 25639 27999
rect 25697 27965 25731 27999
rect 28549 27897 28583 27931
rect 28641 27897 28675 27931
rect 8309 27829 8343 27863
rect 9413 27829 9447 27863
rect 12173 27829 12207 27863
rect 12725 27829 12759 27863
rect 13553 27829 13587 27863
rect 17693 27829 17727 27863
rect 25145 27829 25179 27863
rect 27169 27829 27203 27863
rect 47685 27829 47719 27863
rect 11976 27625 12010 27659
rect 19993 27625 20027 27659
rect 25605 27625 25639 27659
rect 27261 27625 27295 27659
rect 26341 27557 26375 27591
rect 27721 27557 27755 27591
rect 28733 27557 28767 27591
rect 33057 27557 33091 27591
rect 8953 27489 8987 27523
rect 11713 27489 11747 27523
rect 21281 27489 21315 27523
rect 21465 27489 21499 27523
rect 25329 27489 25363 27523
rect 27353 27489 27387 27523
rect 28825 27489 28859 27523
rect 30573 27489 30607 27523
rect 33977 27489 34011 27523
rect 36185 27489 36219 27523
rect 39865 27489 39899 27523
rect 40325 27489 40359 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 48145 27489 48179 27523
rect 8401 27421 8435 27455
rect 14197 27421 14231 27455
rect 14381 27421 14415 27455
rect 14841 27421 14875 27455
rect 17049 27421 17083 27455
rect 18245 27421 18279 27455
rect 18337 27421 18371 27455
rect 18429 27421 18463 27455
rect 18613 27421 18647 27455
rect 19349 27421 19383 27455
rect 20177 27421 20211 27455
rect 22109 27421 22143 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 26249 27421 26283 27455
rect 27537 27421 27571 27455
rect 28549 27421 28583 27455
rect 30757 27421 30791 27455
rect 32965 27421 32999 27455
rect 33793 27421 33827 27455
rect 35357 27421 35391 27455
rect 9229 27353 9263 27387
rect 15117 27353 15151 27387
rect 17141 27353 17175 27387
rect 22293 27353 22327 27387
rect 27261 27353 27295 27387
rect 33609 27353 33643 27387
rect 40049 27353 40083 27387
rect 8217 27285 8251 27319
rect 10701 27285 10735 27319
rect 13461 27285 13495 27319
rect 16589 27285 16623 27319
rect 17969 27285 18003 27319
rect 19441 27285 19475 27319
rect 20821 27285 20855 27319
rect 21189 27285 21223 27319
rect 24409 27285 24443 27319
rect 28365 27285 28399 27319
rect 30941 27285 30975 27319
rect 9689 27081 9723 27115
rect 10701 27081 10735 27115
rect 13185 27081 13219 27115
rect 15301 27081 15335 27115
rect 18429 27081 18463 27115
rect 25329 27081 25363 27115
rect 33425 27081 33459 27115
rect 39957 27081 39991 27115
rect 10425 27013 10459 27047
rect 23857 27013 23891 27047
rect 33241 27013 33275 27047
rect 8677 26945 8711 26979
rect 9505 26945 9539 26979
rect 10609 26945 10643 26979
rect 10793 26945 10827 26979
rect 13001 26945 13035 26979
rect 15485 26945 15519 26979
rect 15761 26945 15795 26979
rect 15945 26945 15979 26979
rect 18245 26945 18279 26979
rect 23581 26945 23615 26979
rect 29285 26945 29319 26979
rect 30297 26945 30331 26979
rect 31125 26945 31159 26979
rect 31249 26945 31283 26979
rect 31401 26945 31435 26979
rect 31503 26951 31537 26985
rect 32137 26945 32171 26979
rect 32321 26945 32355 26979
rect 33517 26945 33551 26979
rect 33977 26945 34011 26979
rect 34161 26945 34195 26979
rect 35265 26945 35299 26979
rect 39865 26945 39899 26979
rect 9321 26877 9355 26911
rect 11529 26877 11563 26911
rect 11805 26877 11839 26911
rect 29009 26877 29043 26911
rect 32229 26877 32263 26911
rect 34069 26877 34103 26911
rect 10977 26809 11011 26843
rect 8769 26741 8803 26775
rect 30389 26741 30423 26775
rect 30941 26741 30975 26775
rect 33241 26741 33275 26775
rect 35357 26741 35391 26775
rect 24593 26537 24627 26571
rect 25237 26537 25271 26571
rect 10333 26469 10367 26503
rect 11621 26469 11655 26503
rect 16405 26469 16439 26503
rect 26985 26469 27019 26503
rect 14105 26401 14139 26435
rect 15485 26401 15519 26435
rect 26525 26401 26559 26435
rect 35541 26401 35575 26435
rect 8217 26333 8251 26367
rect 9229 26333 9263 26367
rect 9505 26333 9539 26367
rect 9965 26333 9999 26367
rect 10149 26333 10183 26367
rect 11069 26333 11103 26367
rect 11529 26333 11563 26367
rect 11713 26333 11747 26367
rect 13369 26333 13403 26367
rect 16405 26333 16439 26367
rect 16681 26333 16715 26367
rect 24409 26333 24443 26367
rect 25145 26333 25179 26367
rect 26617 26333 26651 26367
rect 27445 26333 27479 26367
rect 27629 26333 27663 26367
rect 28089 26333 28123 26367
rect 28237 26333 28271 26367
rect 28554 26333 28588 26367
rect 30665 26333 30699 26367
rect 33057 26333 33091 26367
rect 33149 26333 33183 26367
rect 33333 26333 33367 26367
rect 33425 26333 33459 26367
rect 33885 26333 33919 26367
rect 35357 26333 35391 26367
rect 45017 26333 45051 26367
rect 47685 26333 47719 26367
rect 10793 26265 10827 26299
rect 10977 26265 11011 26299
rect 13461 26265 13495 26299
rect 14289 26265 14323 26299
rect 28365 26265 28399 26299
rect 28457 26265 28491 26299
rect 30941 26265 30975 26299
rect 33977 26265 34011 26299
rect 8217 26197 8251 26231
rect 9045 26197 9079 26231
rect 9413 26197 9447 26231
rect 11069 26197 11103 26231
rect 16589 26197 16623 26231
rect 27537 26197 27571 26231
rect 28733 26197 28767 26231
rect 32413 26197 32447 26231
rect 32873 26197 32907 26231
rect 45109 26197 45143 26231
rect 10793 25993 10827 26027
rect 16129 25993 16163 26027
rect 16957 25993 16991 26027
rect 23489 25993 23523 26027
rect 30297 25993 30331 26027
rect 31493 25993 31527 26027
rect 34253 25993 34287 26027
rect 8217 25925 8251 25959
rect 10609 25925 10643 25959
rect 15761 25925 15795 25959
rect 15977 25925 16011 25959
rect 16773 25925 16807 25959
rect 17325 25925 17359 25959
rect 23305 25925 23339 25959
rect 28825 25925 28859 25959
rect 32781 25925 32815 25959
rect 35541 25925 35575 25959
rect 45293 25925 45327 25959
rect 7941 25857 7975 25891
rect 11713 25857 11747 25891
rect 14657 25857 14691 25891
rect 17049 25857 17083 25891
rect 17141 25857 17175 25891
rect 17785 25857 17819 25891
rect 19073 25857 19107 25891
rect 19901 25857 19935 25891
rect 22063 25857 22097 25891
rect 22198 25857 22232 25891
rect 22293 25857 22327 25891
rect 22477 25857 22511 25891
rect 22937 25857 22971 25891
rect 23121 25857 23155 25891
rect 23213 25857 23247 25891
rect 24685 25857 24719 25891
rect 26985 25857 27019 25891
rect 27078 25857 27112 25891
rect 27261 25857 27295 25891
rect 27353 25857 27387 25891
rect 27450 25857 27484 25891
rect 28549 25857 28583 25891
rect 31401 25857 31435 25891
rect 32505 25857 32539 25891
rect 35265 25857 35299 25891
rect 36185 25857 36219 25891
rect 19993 25789 20027 25823
rect 24961 25789 24995 25823
rect 45109 25789 45143 25823
rect 46857 25789 46891 25823
rect 9689 25721 9723 25755
rect 10241 25721 10275 25755
rect 17877 25721 17911 25755
rect 19165 25721 19199 25755
rect 21833 25721 21867 25755
rect 26433 25721 26467 25755
rect 27629 25721 27663 25755
rect 10609 25653 10643 25687
rect 11529 25653 11563 25687
rect 14841 25653 14875 25687
rect 15945 25653 15979 25687
rect 20269 25653 20303 25687
rect 36277 25653 36311 25687
rect 47777 25653 47811 25687
rect 14289 25449 14323 25483
rect 16773 25449 16807 25483
rect 22017 25449 22051 25483
rect 22661 25449 22695 25483
rect 25145 25449 25179 25483
rect 29929 25449 29963 25483
rect 33609 25449 33643 25483
rect 21005 25381 21039 25415
rect 22845 25381 22879 25415
rect 10425 25313 10459 25347
rect 10517 25313 10551 25347
rect 10885 25313 10919 25347
rect 11437 25313 11471 25347
rect 15025 25313 15059 25347
rect 17509 25313 17543 25347
rect 17785 25313 17819 25347
rect 19533 25313 19567 25347
rect 29561 25313 29595 25347
rect 33241 25313 33275 25347
rect 35909 25313 35943 25347
rect 46305 25313 46339 25347
rect 10793 25245 10827 25279
rect 11529 25245 11563 25279
rect 12449 25245 12483 25279
rect 14105 25245 14139 25279
rect 17417 25245 17451 25279
rect 18521 25245 18555 25279
rect 19257 25245 19291 25279
rect 21741 25245 21775 25279
rect 21833 25245 21867 25279
rect 25053 25245 25087 25279
rect 29745 25245 29779 25279
rect 33425 25245 33459 25279
rect 34897 25245 34931 25279
rect 35725 25245 35759 25279
rect 1869 25177 1903 25211
rect 15301 25177 15335 25211
rect 22477 25177 22511 25211
rect 37565 25177 37599 25211
rect 46489 25177 46523 25211
rect 48145 25177 48179 25211
rect 1961 25109 1995 25143
rect 10241 25109 10275 25143
rect 10701 25109 10735 25143
rect 11897 25109 11931 25143
rect 12541 25109 12575 25143
rect 18613 25109 18647 25143
rect 22687 25109 22721 25143
rect 34989 25109 35023 25143
rect 13553 24905 13587 24939
rect 15945 24905 15979 24939
rect 23581 24905 23615 24939
rect 12081 24837 12115 24871
rect 34437 24837 34471 24871
rect 14105 24769 14139 24803
rect 14933 24769 14967 24803
rect 15853 24769 15887 24803
rect 16037 24769 16071 24803
rect 20085 24769 20119 24803
rect 21281 24769 21315 24803
rect 25053 24769 25087 24803
rect 26985 24769 27019 24803
rect 28641 24769 28675 24803
rect 28825 24769 28859 24803
rect 32137 24769 32171 24803
rect 33609 24769 33643 24803
rect 33701 24769 33735 24803
rect 36093 24769 36127 24803
rect 46397 24769 46431 24803
rect 46857 24769 46891 24803
rect 46949 24769 46983 24803
rect 47593 24769 47627 24803
rect 11805 24701 11839 24735
rect 17785 24701 17819 24735
rect 18061 24701 18095 24735
rect 21833 24701 21867 24735
rect 22109 24701 22143 24735
rect 34253 24701 34287 24735
rect 20177 24633 20211 24667
rect 21097 24633 21131 24667
rect 46213 24633 46247 24667
rect 14197 24565 14231 24599
rect 15117 24565 15151 24599
rect 19533 24565 19567 24599
rect 25145 24565 25179 24599
rect 27169 24565 27203 24599
rect 28733 24565 28767 24599
rect 32321 24565 32355 24599
rect 47685 24565 47719 24599
rect 13277 24361 13311 24395
rect 19441 24361 19475 24395
rect 21189 24361 21223 24395
rect 22477 24361 22511 24395
rect 33609 24361 33643 24395
rect 10057 24293 10091 24327
rect 12633 24293 12667 24327
rect 22385 24293 22419 24327
rect 23029 24293 23063 24327
rect 29561 24293 29595 24327
rect 14105 24225 14139 24259
rect 14289 24225 14323 24259
rect 15577 24225 15611 24259
rect 18245 24225 18279 24259
rect 23397 24225 23431 24259
rect 25145 24225 25179 24259
rect 26801 24225 26835 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 9137 24157 9171 24191
rect 10609 24157 10643 24191
rect 12449 24157 12483 24191
rect 13185 24157 13219 24191
rect 16405 24157 16439 24191
rect 19441 24157 19475 24191
rect 21189 24157 21223 24191
rect 22017 24157 22051 24191
rect 23213 24157 23247 24191
rect 23305 24157 23339 24191
rect 23489 24157 23523 24191
rect 24961 24157 24995 24191
rect 27261 24157 27295 24191
rect 27537 24157 27571 24191
rect 29745 24157 29779 24191
rect 29846 24157 29880 24191
rect 30481 24157 30515 24191
rect 31677 24157 31711 24191
rect 33517 24157 33551 24191
rect 35081 24157 35115 24191
rect 36921 24157 36955 24191
rect 43085 24157 43119 24191
rect 43269 24157 43303 24191
rect 43913 24157 43947 24191
rect 44097 24157 44131 24191
rect 45661 24157 45695 24191
rect 45845 24157 45879 24191
rect 9689 24089 9723 24123
rect 16589 24089 16623 24123
rect 28641 24089 28675 24123
rect 28825 24089 28859 24123
rect 29561 24089 29595 24123
rect 35265 24089 35299 24123
rect 43453 24089 43487 24123
rect 9137 24021 9171 24055
rect 10149 24021 10183 24055
rect 10701 24021 10735 24055
rect 29009 24021 29043 24055
rect 30297 24021 30331 24055
rect 31769 24021 31803 24055
rect 44005 24021 44039 24055
rect 45845 24021 45879 24055
rect 15853 23817 15887 23851
rect 16773 23817 16807 23851
rect 22385 23817 22419 23851
rect 31493 23817 31527 23851
rect 35817 23817 35851 23851
rect 8493 23749 8527 23783
rect 9229 23749 9263 23783
rect 15761 23749 15795 23783
rect 25605 23749 25639 23783
rect 30021 23749 30055 23783
rect 32229 23749 32263 23783
rect 35265 23749 35299 23783
rect 42441 23749 42475 23783
rect 42625 23749 42659 23783
rect 45109 23749 45143 23783
rect 1869 23681 1903 23715
rect 8401 23681 8435 23715
rect 13093 23681 13127 23715
rect 16681 23681 16715 23715
rect 17509 23681 17543 23715
rect 19533 23681 19567 23715
rect 22293 23681 22327 23715
rect 23029 23681 23063 23715
rect 23949 23681 23983 23715
rect 27445 23681 27479 23715
rect 28365 23681 28399 23715
rect 29745 23681 29779 23715
rect 32137 23681 32171 23715
rect 33517 23681 33551 23715
rect 35725 23681 35759 23715
rect 39221 23681 39255 23715
rect 40049 23681 40083 23715
rect 42717 23681 42751 23715
rect 43269 23681 43303 23715
rect 44005 23681 44039 23715
rect 45753 23681 45787 23715
rect 47593 23681 47627 23715
rect 9045 23613 9079 23647
rect 10885 23613 10919 23647
rect 13277 23613 13311 23647
rect 14013 23613 14047 23647
rect 17877 23613 17911 23647
rect 23673 23613 23707 23647
rect 27537 23613 27571 23647
rect 28641 23613 28675 23647
rect 39129 23613 39163 23647
rect 40233 23613 40267 23647
rect 41889 23613 41923 23647
rect 46213 23613 46247 23647
rect 46489 23613 46523 23647
rect 48053 23613 48087 23647
rect 2053 23545 2087 23579
rect 25789 23545 25823 23579
rect 19625 23477 19659 23511
rect 23121 23477 23155 23511
rect 27813 23477 27847 23511
rect 39497 23477 39531 23511
rect 42441 23477 42475 23511
rect 45569 23477 45603 23511
rect 47685 23477 47719 23511
rect 10793 23273 10827 23307
rect 13093 23273 13127 23307
rect 18429 23273 18463 23307
rect 25513 23273 25547 23307
rect 28733 23273 28767 23307
rect 29929 23273 29963 23307
rect 32137 23273 32171 23307
rect 24777 23205 24811 23239
rect 25697 23205 25731 23239
rect 28917 23205 28951 23239
rect 43269 23205 43303 23239
rect 44281 23205 44315 23239
rect 9045 23137 9079 23171
rect 19533 23137 19567 23171
rect 22109 23137 22143 23171
rect 24409 23137 24443 23171
rect 24869 23137 24903 23171
rect 26525 23137 26559 23171
rect 29561 23137 29595 23171
rect 30665 23137 30699 23171
rect 40049 23137 40083 23171
rect 40877 23137 40911 23171
rect 42625 23137 42659 23171
rect 45753 23137 45787 23171
rect 45937 23137 45971 23171
rect 46949 23137 46983 23171
rect 11345 23069 11379 23103
rect 12909 23069 12943 23103
rect 15761 23069 15795 23103
rect 17601 23069 17635 23103
rect 18153 23069 18187 23103
rect 19257 23069 19291 23103
rect 21833 23069 21867 23103
rect 24593 23069 24627 23103
rect 26249 23069 26283 23103
rect 29745 23069 29779 23103
rect 30389 23069 30423 23103
rect 33977 23069 34011 23103
rect 34713 23069 34747 23103
rect 40325 23069 40359 23103
rect 42349 23069 42383 23103
rect 43269 23069 43303 23103
rect 43453 23069 43487 23103
rect 44465 23069 44499 23103
rect 9321 23001 9355 23035
rect 14565 23001 14599 23035
rect 15945 23001 15979 23035
rect 25329 23001 25363 23035
rect 28549 23001 28583 23035
rect 33241 23001 33275 23035
rect 41521 23001 41555 23035
rect 45109 23001 45143 23035
rect 45293 23001 45327 23035
rect 11437 22933 11471 22967
rect 14657 22933 14691 22967
rect 21005 22933 21039 22967
rect 23581 22933 23615 22967
rect 25529 22933 25563 22967
rect 27997 22933 28031 22967
rect 28749 22933 28783 22967
rect 34897 22933 34931 22967
rect 41613 22933 41647 22967
rect 9597 22729 9631 22763
rect 13921 22729 13955 22763
rect 21097 22729 21131 22763
rect 22017 22729 22051 22763
rect 22845 22729 22879 22763
rect 23397 22729 23431 22763
rect 23857 22729 23891 22763
rect 23949 22729 23983 22763
rect 26341 22729 26375 22763
rect 27267 22729 27301 22763
rect 27445 22729 27479 22763
rect 29193 22729 29227 22763
rect 30113 22729 30147 22763
rect 40877 22729 40911 22763
rect 43085 22729 43119 22763
rect 48145 22729 48179 22763
rect 11713 22661 11747 22695
rect 24501 22661 24535 22695
rect 45385 22661 45419 22695
rect 24731 22627 24765 22661
rect 9781 22593 9815 22627
rect 11529 22593 11563 22627
rect 13829 22593 13863 22627
rect 15025 22593 15059 22627
rect 15853 22593 15887 22627
rect 19165 22593 19199 22627
rect 19901 22593 19935 22627
rect 20913 22593 20947 22627
rect 21833 22593 21867 22627
rect 22753 22593 22787 22627
rect 23581 22593 23615 22627
rect 24041 22593 24075 22627
rect 25513 22593 25547 22627
rect 25697 22593 25731 22627
rect 26249 22593 26283 22627
rect 27353 22593 27387 22627
rect 29101 22593 29135 22627
rect 29285 22593 29319 22627
rect 29929 22593 29963 22627
rect 39957 22593 39991 22627
rect 41061 22593 41095 22627
rect 42993 22593 43027 22627
rect 43177 22593 43211 22627
rect 45201 22593 45235 22627
rect 47593 22593 47627 22627
rect 13369 22525 13403 22559
rect 16957 22525 16991 22559
rect 17233 22525 17267 22559
rect 23673 22525 23707 22559
rect 25789 22525 25823 22559
rect 27721 22525 27755 22559
rect 40417 22525 40451 22559
rect 43913 22525 43947 22559
rect 44189 22525 44223 22559
rect 46949 22525 46983 22559
rect 47869 22525 47903 22559
rect 15209 22457 15243 22491
rect 19349 22457 19383 22491
rect 25329 22457 25363 22491
rect 16037 22389 16071 22423
rect 18705 22389 18739 22423
rect 20085 22389 20119 22423
rect 24685 22389 24719 22423
rect 24869 22389 24903 22423
rect 26985 22389 27019 22423
rect 27629 22389 27663 22423
rect 40049 22389 40083 22423
rect 47685 22389 47719 22423
rect 15485 22185 15519 22219
rect 16865 22185 16899 22219
rect 26341 22185 26375 22219
rect 27721 22185 27755 22219
rect 29929 22185 29963 22219
rect 9597 22049 9631 22083
rect 16589 22049 16623 22083
rect 18613 22049 18647 22083
rect 21833 22049 21867 22083
rect 47133 22049 47167 22083
rect 12449 21981 12483 22015
rect 13093 21981 13127 22015
rect 14105 21981 14139 22015
rect 15393 21981 15427 22015
rect 16497 21981 16531 22015
rect 17417 21981 17451 22015
rect 18521 21981 18555 22015
rect 19257 21981 19291 22015
rect 19993 21981 20027 22015
rect 23673 21981 23707 22015
rect 23857 21981 23891 22015
rect 24685 21981 24719 22015
rect 26157 21981 26191 22015
rect 29745 21981 29779 22015
rect 39957 21981 39991 22015
rect 40141 21981 40175 22015
rect 42533 21981 42567 22015
rect 42717 21981 42751 22015
rect 43821 21981 43855 22015
rect 45385 21981 45419 22015
rect 46857 21981 46891 22015
rect 9781 21913 9815 21947
rect 11437 21913 11471 21947
rect 17877 21913 17911 21947
rect 20177 21913 20211 21947
rect 24409 21913 24443 21947
rect 24593 21913 24627 21947
rect 27537 21913 27571 21947
rect 40325 21913 40359 21947
rect 44281 21913 44315 21947
rect 46213 21913 46247 21947
rect 12541 21845 12575 21879
rect 13277 21845 13311 21879
rect 14289 21845 14323 21879
rect 19441 21845 19475 21879
rect 23765 21845 23799 21879
rect 24507 21845 24541 21879
rect 27737 21845 27771 21879
rect 27905 21845 27939 21879
rect 42901 21845 42935 21879
rect 9965 21641 9999 21675
rect 27553 21641 27587 21675
rect 27721 21641 27755 21675
rect 42809 21641 42843 21675
rect 47777 21641 47811 21675
rect 17509 21573 17543 21607
rect 21005 21573 21039 21607
rect 27353 21573 27387 21607
rect 30941 21573 30975 21607
rect 31033 21573 31067 21607
rect 41797 21573 41831 21607
rect 47593 21573 47627 21607
rect 9229 21505 9263 21539
rect 9873 21505 9907 21539
rect 10701 21505 10735 21539
rect 14289 21505 14323 21539
rect 17417 21505 17451 21539
rect 20085 21505 20119 21539
rect 20913 21505 20947 21539
rect 21833 21505 21867 21539
rect 22753 21505 22787 21539
rect 23581 21505 23615 21539
rect 23765 21505 23799 21539
rect 26249 21505 26283 21539
rect 41705 21505 41739 21539
rect 41889 21505 41923 21539
rect 42993 21505 43027 21539
rect 43177 21505 43211 21539
rect 43269 21505 43303 21539
rect 44005 21505 44039 21539
rect 44557 21505 44591 21539
rect 45477 21505 45511 21539
rect 47869 21505 47903 21539
rect 47961 21505 47995 21539
rect 10977 21437 11011 21471
rect 11621 21437 11655 21471
rect 11897 21437 11931 21471
rect 14565 21437 14599 21471
rect 22845 21437 22879 21471
rect 32137 21437 32171 21471
rect 32321 21437 32355 21471
rect 32597 21437 32631 21471
rect 44097 21437 44131 21471
rect 44833 21437 44867 21471
rect 46213 21437 46247 21471
rect 20361 21369 20395 21403
rect 31493 21369 31527 21403
rect 48145 21369 48179 21403
rect 9321 21301 9355 21335
rect 13369 21301 13403 21335
rect 16037 21301 16071 21335
rect 21925 21301 21959 21335
rect 23121 21301 23155 21335
rect 23581 21301 23615 21335
rect 26341 21301 26375 21335
rect 27537 21301 27571 21335
rect 11437 21097 11471 21131
rect 30941 21097 30975 21131
rect 31217 21097 31251 21131
rect 32045 21097 32079 21131
rect 34805 21097 34839 21131
rect 35449 21097 35483 21131
rect 12081 21029 12115 21063
rect 13369 21029 13403 21063
rect 15761 21029 15795 21063
rect 41705 21029 41739 21063
rect 9597 20961 9631 20995
rect 9873 20961 9907 20995
rect 14657 20961 14691 20995
rect 21097 20961 21131 20995
rect 21373 20961 21407 20995
rect 26157 20961 26191 20995
rect 26433 20961 26467 20995
rect 27169 20961 27203 20995
rect 30021 20961 30055 20995
rect 30389 20961 30423 20995
rect 31585 20961 31619 20995
rect 35173 20961 35207 20995
rect 42257 20961 42291 20995
rect 42993 20961 43027 20995
rect 46305 20961 46339 20995
rect 48145 20961 48179 20995
rect 9505 20893 9539 20927
rect 11437 20893 11471 20927
rect 11621 20893 11655 20927
rect 12357 20893 12391 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 14473 20893 14507 20927
rect 15669 20893 15703 20927
rect 19257 20893 19291 20927
rect 26065 20893 26099 20927
rect 26893 20893 26927 20927
rect 31125 20893 31159 20927
rect 32229 20893 32263 20927
rect 34713 20893 34747 20927
rect 42165 20893 42199 20927
rect 42349 20893 42383 20927
rect 43269 20893 43303 20927
rect 45385 20893 45419 20927
rect 12081 20825 12115 20859
rect 30113 20825 30147 20859
rect 45661 20825 45695 20859
rect 46489 20825 46523 20859
rect 12265 20757 12299 20791
rect 19349 20757 19383 20791
rect 22845 20757 22879 20791
rect 28641 20757 28675 20791
rect 43913 20757 43947 20791
rect 12725 20553 12759 20587
rect 14289 20553 14323 20587
rect 14749 20553 14783 20587
rect 17325 20553 17359 20587
rect 22109 20553 22143 20587
rect 27169 20553 27203 20587
rect 27813 20553 27847 20587
rect 36185 20553 36219 20587
rect 47961 20553 47995 20587
rect 9321 20485 9355 20519
rect 12357 20485 12391 20519
rect 12557 20485 12591 20519
rect 18889 20485 18923 20519
rect 23213 20485 23247 20519
rect 34713 20485 34747 20519
rect 34805 20485 34839 20519
rect 45385 20485 45419 20519
rect 47593 20485 47627 20519
rect 9137 20417 9171 20451
rect 11529 20417 11563 20451
rect 13645 20417 13679 20451
rect 13829 20417 13863 20451
rect 16957 20417 16991 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 22017 20417 22051 20451
rect 25697 20417 25731 20451
rect 25881 20417 25915 20451
rect 26985 20417 27019 20451
rect 27261 20417 27295 20451
rect 27721 20417 27755 20451
rect 31493 20417 31527 20451
rect 32321 20417 32355 20451
rect 36369 20417 36403 20451
rect 42717 20417 42751 20451
rect 42901 20417 42935 20451
rect 43821 20417 43855 20451
rect 44465 20417 44499 20451
rect 44649 20417 44683 20451
rect 47777 20417 47811 20451
rect 9597 20349 9631 20383
rect 14473 20349 14507 20383
rect 14565 20349 14599 20383
rect 14841 20349 14875 20383
rect 14933 20349 14967 20383
rect 18705 20349 18739 20383
rect 19349 20349 19383 20383
rect 22937 20349 22971 20383
rect 24961 20349 24995 20383
rect 32505 20349 32539 20383
rect 34161 20349 34195 20383
rect 35725 20349 35759 20383
rect 43637 20349 43671 20383
rect 45201 20349 45235 20383
rect 47041 20349 47075 20383
rect 16773 20281 16807 20315
rect 26985 20281 27019 20315
rect 31309 20281 31343 20315
rect 42717 20281 42751 20315
rect 44465 20281 44499 20315
rect 11621 20213 11655 20247
rect 12541 20213 12575 20247
rect 13737 20213 13771 20247
rect 25697 20213 25731 20247
rect 44005 20213 44039 20247
rect 11621 20009 11655 20043
rect 15025 20009 15059 20043
rect 16313 20009 16347 20043
rect 22937 20009 22971 20043
rect 23581 20009 23615 20043
rect 43637 20009 43671 20043
rect 45385 20009 45419 20043
rect 14473 19941 14507 19975
rect 16497 19941 16531 19975
rect 30941 19941 30975 19975
rect 10149 19873 10183 19907
rect 17233 19873 17267 19907
rect 17509 19873 17543 19907
rect 25697 19873 25731 19907
rect 30113 19873 30147 19907
rect 35173 19873 35207 19907
rect 36185 19873 36219 19907
rect 47041 19873 47075 19907
rect 2053 19805 2087 19839
rect 9873 19805 9907 19839
rect 12173 19805 12207 19839
rect 14841 19805 14875 19839
rect 17141 19805 17175 19839
rect 18153 19805 18187 19839
rect 20729 19805 20763 19839
rect 22753 19805 22787 19839
rect 23489 19805 23523 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 25421 19805 25455 19839
rect 29745 19805 29779 19839
rect 30573 19805 30607 19839
rect 30757 19805 30791 19839
rect 33793 19805 33827 19839
rect 42993 19805 43027 19839
rect 43177 19805 43211 19839
rect 43821 19805 43855 19839
rect 44097 19805 44131 19839
rect 45293 19805 45327 19839
rect 45937 19805 45971 19839
rect 14749 19737 14783 19771
rect 16129 19737 16163 19771
rect 16345 19737 16379 19771
rect 29929 19737 29963 19771
rect 35265 19737 35299 19771
rect 43085 19737 43119 19771
rect 44005 19737 44039 19771
rect 46121 19737 46155 19771
rect 12357 19669 12391 19703
rect 14657 19669 14691 19703
rect 18153 19669 18187 19703
rect 20821 19669 20855 19703
rect 27169 19669 27203 19703
rect 33885 19669 33919 19703
rect 10517 19465 10551 19499
rect 27077 19465 27111 19499
rect 29929 19465 29963 19499
rect 33241 19465 33275 19499
rect 47961 19465 47995 19499
rect 16129 19397 16163 19431
rect 33885 19397 33919 19431
rect 46305 19397 46339 19431
rect 47869 19397 47903 19431
rect 1777 19329 1811 19363
rect 10425 19329 10459 19363
rect 12173 19329 12207 19363
rect 13001 19329 13035 19363
rect 14473 19329 14507 19363
rect 15945 19329 15979 19363
rect 16957 19329 16991 19363
rect 17785 19329 17819 19363
rect 20729 19329 20763 19363
rect 24317 19329 24351 19363
rect 24501 19329 24535 19363
rect 26985 19329 27019 19363
rect 29745 19329 29779 19363
rect 29929 19329 29963 19363
rect 32321 19329 32355 19363
rect 32781 19329 32815 19363
rect 33701 19329 33735 19363
rect 35541 19329 35575 19363
rect 37289 19329 37323 19363
rect 39129 19329 39163 19363
rect 44557 19329 44591 19363
rect 46397 19329 46431 19363
rect 46765 19329 46799 19363
rect 47041 19329 47075 19363
rect 47777 19329 47811 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 12265 19261 12299 19295
rect 14381 19261 14415 19295
rect 15761 19261 15795 19295
rect 16865 19261 16899 19295
rect 17049 19261 17083 19295
rect 17141 19261 17175 19295
rect 18061 19261 18095 19295
rect 19533 19261 19567 19295
rect 21833 19261 21867 19295
rect 22109 19261 22143 19295
rect 37473 19261 37507 19295
rect 44281 19261 44315 19295
rect 45109 19261 45143 19295
rect 46029 19261 46063 19295
rect 48145 19261 48179 19295
rect 23581 19193 23615 19227
rect 47593 19193 47627 19227
rect 12541 19125 12575 19159
rect 13093 19125 13127 19159
rect 14749 19125 14783 19159
rect 16681 19125 16715 19159
rect 20913 19125 20947 19159
rect 24317 19125 24351 19159
rect 32137 19125 32171 19159
rect 33057 19125 33091 19159
rect 43637 19125 43671 19159
rect 2237 18921 2271 18955
rect 16221 18853 16255 18887
rect 17325 18853 17359 18887
rect 19349 18853 19383 18887
rect 23029 18853 23063 18887
rect 24501 18853 24535 18887
rect 37197 18853 37231 18887
rect 11713 18785 11747 18819
rect 11989 18785 12023 18819
rect 14749 18785 14783 18819
rect 20637 18785 20671 18819
rect 20821 18785 20855 18819
rect 26525 18785 26559 18819
rect 28917 18785 28951 18819
rect 29837 18785 29871 18819
rect 30297 18785 30331 18819
rect 31033 18785 31067 18819
rect 46305 18785 46339 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 14473 18717 14507 18751
rect 17049 18717 17083 18751
rect 18337 18717 18371 18751
rect 19257 18717 19291 18751
rect 19901 18717 19935 18751
rect 22937 18717 22971 18751
rect 23673 18717 23707 18751
rect 24777 18717 24811 18751
rect 25881 18717 25915 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29929 18717 29963 18751
rect 30573 18717 30607 18751
rect 32781 18717 32815 18751
rect 33149 18717 33183 18751
rect 33333 18717 33367 18751
rect 33609 18717 33643 18751
rect 37105 18717 37139 18751
rect 44005 18717 44039 18751
rect 44189 18717 44223 18751
rect 45201 18717 45235 18751
rect 45385 18717 45419 18751
rect 22477 18649 22511 18683
rect 24501 18649 24535 18683
rect 25973 18649 26007 18683
rect 26709 18649 26743 18683
rect 28365 18649 28399 18683
rect 30757 18649 30791 18683
rect 33793 18649 33827 18683
rect 44097 18649 44131 18683
rect 46489 18649 46523 18683
rect 13461 18581 13495 18615
rect 17509 18581 17543 18615
rect 18337 18581 18371 18615
rect 19993 18581 20027 18615
rect 23765 18581 23799 18615
rect 24685 18581 24719 18615
rect 45293 18581 45327 18615
rect 14105 18377 14139 18411
rect 15853 18377 15887 18411
rect 22017 18377 22051 18411
rect 30021 18377 30055 18411
rect 31033 18377 31067 18411
rect 44005 18377 44039 18411
rect 47685 18377 47719 18411
rect 23305 18309 23339 18343
rect 29653 18309 29687 18343
rect 32321 18309 32355 18343
rect 34621 18309 34655 18343
rect 46397 18309 46431 18343
rect 1409 18241 1443 18275
rect 14013 18241 14047 18275
rect 15761 18241 15795 18275
rect 17601 18241 17635 18275
rect 18061 18241 18095 18275
rect 21833 18241 21867 18275
rect 25421 18241 25455 18275
rect 26157 18241 26191 18275
rect 28089 18241 28123 18275
rect 28733 18241 28767 18275
rect 29837 18241 29871 18275
rect 30941 18241 30975 18275
rect 32137 18241 32171 18275
rect 34437 18241 34471 18275
rect 44189 18241 44223 18275
rect 44741 18241 44775 18275
rect 46213 18241 46247 18275
rect 47593 18241 47627 18275
rect 18337 18173 18371 18207
rect 23121 18173 23155 18207
rect 23581 18173 23615 18207
rect 29009 18173 29043 18207
rect 29101 18173 29135 18207
rect 33977 18173 34011 18207
rect 36277 18173 36311 18207
rect 45661 18173 45695 18207
rect 1593 18105 1627 18139
rect 17417 18105 17451 18139
rect 28181 18105 28215 18139
rect 46581 18105 46615 18139
rect 19809 18037 19843 18071
rect 25421 18037 25455 18071
rect 26249 18037 26283 18071
rect 28825 18037 28859 18071
rect 29101 18037 29135 18071
rect 22937 17833 22971 17867
rect 24961 17833 24995 17867
rect 45661 17833 45695 17867
rect 28457 17765 28491 17799
rect 19993 17697 20027 17731
rect 23397 17697 23431 17731
rect 24409 17697 24443 17731
rect 25697 17697 25731 17731
rect 25973 17697 26007 17731
rect 44373 17697 44407 17731
rect 45385 17697 45419 17731
rect 45477 17697 45511 17731
rect 23121 17629 23155 17663
rect 23305 17629 23339 17663
rect 25605 17629 25639 17663
rect 26433 17629 26467 17663
rect 27077 17629 27111 17663
rect 27813 17629 27847 17663
rect 27997 17629 28031 17663
rect 28641 17629 28675 17663
rect 29653 17629 29687 17663
rect 29837 17629 29871 17663
rect 44281 17629 44315 17663
rect 44465 17629 44499 17663
rect 45017 17629 45051 17663
rect 46305 17629 46339 17663
rect 20177 17561 20211 17595
rect 21833 17561 21867 17595
rect 24685 17561 24719 17595
rect 27905 17561 27939 17595
rect 29009 17561 29043 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 24593 17493 24627 17527
rect 24777 17493 24811 17527
rect 26525 17493 26559 17527
rect 27169 17493 27203 17527
rect 28733 17493 28767 17527
rect 28825 17493 28859 17527
rect 30665 17493 30699 17527
rect 20177 17289 20211 17323
rect 28825 17289 28859 17323
rect 29653 17289 29687 17323
rect 47685 17289 47719 17323
rect 21189 17221 21223 17255
rect 22017 17221 22051 17255
rect 24409 17221 24443 17255
rect 20085 17153 20119 17187
rect 21097 17153 21131 17187
rect 27905 17153 27939 17187
rect 28089 17153 28123 17187
rect 28641 17153 28675 17187
rect 28825 17153 28859 17187
rect 29469 17153 29503 17187
rect 33609 17153 33643 17187
rect 47593 17153 47627 17187
rect 21833 17085 21867 17119
rect 22293 17085 22327 17119
rect 24133 17085 24167 17119
rect 29285 17085 29319 17119
rect 33793 17085 33827 17119
rect 35449 17085 35483 17119
rect 45201 17085 45235 17119
rect 45385 17085 45419 17119
rect 46857 17085 46891 17119
rect 27905 17017 27939 17051
rect 2053 16949 2087 16983
rect 25881 16949 25915 16983
rect 24593 16745 24627 16779
rect 24777 16745 24811 16779
rect 29561 16745 29595 16779
rect 33793 16745 33827 16779
rect 48145 16745 48179 16779
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 20177 16609 20211 16643
rect 25973 16609 26007 16643
rect 26249 16609 26283 16643
rect 45017 16609 45051 16643
rect 45477 16609 45511 16643
rect 19533 16541 19567 16575
rect 22477 16541 22511 16575
rect 29561 16541 29595 16575
rect 29745 16541 29779 16575
rect 33701 16541 33735 16575
rect 47317 16541 47351 16575
rect 1593 16473 1627 16507
rect 19625 16473 19659 16507
rect 20361 16473 20395 16507
rect 22017 16473 22051 16507
rect 24409 16473 24443 16507
rect 24625 16473 24659 16507
rect 45201 16473 45235 16507
rect 47409 16473 47443 16507
rect 22569 16405 22603 16439
rect 27721 16405 27755 16439
rect 2145 16201 2179 16235
rect 45201 16201 45235 16235
rect 2053 16065 2087 16099
rect 18521 16065 18555 16099
rect 22753 16065 22787 16099
rect 29745 16065 29779 16099
rect 45109 16065 45143 16099
rect 47777 16065 47811 16099
rect 18705 15997 18739 16031
rect 19993 15997 20027 16031
rect 22937 15997 22971 16031
rect 24593 15997 24627 16031
rect 29929 15997 29963 16031
rect 31401 15997 31435 16031
rect 19349 15657 19383 15691
rect 29929 15657 29963 15691
rect 2053 15453 2087 15487
rect 19257 15453 19291 15487
rect 29837 15453 29871 15487
rect 1777 14977 1811 15011
rect 21005 14977 21039 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 21097 14773 21131 14807
rect 2329 14569 2363 14603
rect 21741 14433 21775 14467
rect 22661 14433 22695 14467
rect 26709 14433 26743 14467
rect 2237 14365 2271 14399
rect 21097 14365 21131 14399
rect 21557 14365 21591 14399
rect 26893 14297 26927 14331
rect 28549 14297 28583 14331
rect 27077 14025 27111 14059
rect 8769 13889 8803 13923
rect 26985 13889 27019 13923
rect 46673 13889 46707 13923
rect 8861 13821 8895 13855
rect 46765 13685 46799 13719
rect 46489 13345 46523 13379
rect 46305 13277 46339 13311
rect 48145 13209 48179 13243
rect 1869 12801 1903 12835
rect 47777 12801 47811 12835
rect 2145 12597 2179 12631
rect 47777 11509 47811 11543
rect 46305 11169 46339 11203
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 47685 10761 47719 10795
rect 47593 10625 47627 10659
rect 47041 10421 47075 10455
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 46489 9945 46523 9979
rect 46949 9605 46983 9639
rect 46857 9537 46891 9571
rect 47869 9537 47903 9571
rect 48053 9401 48087 9435
rect 47869 8925 47903 8959
rect 48053 8789 48087 8823
rect 46121 8449 46155 8483
rect 45845 8245 45879 8279
rect 46213 8245 46247 8279
rect 46581 8245 46615 8279
rect 47225 7905 47259 7939
rect 46397 7837 46431 7871
rect 46949 7769 46983 7803
rect 47041 7769 47075 7803
rect 46213 7701 46247 7735
rect 47961 7497 47995 7531
rect 46121 7429 46155 7463
rect 48145 7361 48179 7395
rect 46029 7293 46063 7327
rect 46305 7293 46339 7327
rect 47317 6817 47351 6851
rect 47593 6749 47627 6783
rect 48053 6409 48087 6443
rect 47961 6273 47995 6307
rect 40233 5661 40267 5695
rect 40325 5525 40359 5559
rect 38669 5321 38703 5355
rect 48053 5321 48087 5355
rect 37473 5253 37507 5287
rect 42625 5253 42659 5287
rect 19625 5185 19659 5219
rect 22569 5185 22603 5219
rect 23489 5185 23523 5219
rect 40049 5185 40083 5219
rect 43821 5185 43855 5219
rect 47869 5185 47903 5219
rect 37381 5117 37415 5151
rect 38301 5117 38335 5151
rect 40233 5117 40267 5151
rect 41889 5117 41923 5151
rect 42533 5117 42567 5151
rect 43545 5117 43579 5151
rect 22661 5049 22695 5083
rect 19717 4981 19751 5015
rect 23305 4981 23339 5015
rect 40233 4777 40267 4811
rect 42349 4777 42383 4811
rect 39221 4709 39255 4743
rect 47593 4641 47627 4675
rect 19349 4573 19383 4607
rect 20361 4573 20395 4607
rect 21005 4573 21039 4607
rect 21649 4573 21683 4607
rect 22293 4573 22327 4607
rect 22937 4573 22971 4607
rect 23581 4573 23615 4607
rect 39129 4573 39163 4607
rect 40417 4573 40451 4607
rect 40877 4573 40911 4607
rect 40969 4573 41003 4607
rect 41521 4573 41555 4607
rect 42533 4573 42567 4607
rect 46673 4573 46707 4607
rect 47317 4573 47351 4607
rect 23029 4505 23063 4539
rect 41613 4505 41647 4539
rect 19441 4437 19475 4471
rect 20453 4437 20487 4471
rect 21097 4437 21131 4471
rect 21741 4437 21775 4471
rect 22385 4437 22419 4471
rect 23673 4437 23707 4471
rect 46765 4437 46799 4471
rect 20729 4233 20763 4267
rect 21925 4233 21959 4267
rect 22569 4233 22603 4267
rect 37289 4233 37323 4267
rect 40877 4233 40911 4267
rect 20085 4165 20119 4199
rect 25421 4165 25455 4199
rect 25513 4165 25547 4199
rect 40049 4165 40083 4199
rect 42809 4165 42843 4199
rect 43729 4165 43763 4199
rect 46673 4165 46707 4199
rect 47777 4165 47811 4199
rect 2145 4097 2179 4131
rect 2789 4097 2823 4131
rect 7481 4097 7515 4131
rect 10057 4097 10091 4131
rect 18613 4097 18647 4131
rect 19257 4097 19291 4131
rect 19993 4097 20027 4131
rect 20637 4097 20671 4131
rect 21833 4097 21867 4131
rect 22477 4097 22511 4131
rect 23121 4097 23155 4131
rect 23765 4097 23799 4131
rect 30113 4097 30147 4131
rect 37473 4097 37507 4131
rect 40509 4097 40543 4131
rect 40693 4097 40727 4131
rect 26433 4029 26467 4063
rect 39405 4029 39439 4063
rect 39589 4029 39623 4063
rect 42717 4029 42751 4063
rect 48053 4029 48087 4063
rect 30205 3961 30239 3995
rect 46857 3961 46891 3995
rect 2237 3893 2271 3927
rect 2881 3893 2915 3927
rect 6837 3893 6871 3927
rect 7573 3893 7607 3927
rect 8309 3893 8343 3927
rect 9505 3893 9539 3927
rect 10149 3893 10183 3927
rect 11713 3893 11747 3927
rect 18705 3893 18739 3927
rect 19349 3893 19383 3927
rect 23213 3893 23247 3927
rect 23857 3893 23891 3927
rect 24869 3893 24903 3927
rect 46121 3893 46155 3927
rect 17693 3689 17727 3723
rect 19625 3689 19659 3723
rect 40325 3689 40359 3723
rect 22569 3621 22603 3655
rect 23213 3621 23247 3655
rect 7113 3553 7147 3587
rect 9321 3553 9355 3587
rect 9505 3553 9539 3587
rect 10701 3553 10735 3587
rect 20637 3553 20671 3587
rect 25605 3553 25639 3587
rect 26617 3553 26651 3587
rect 37657 3553 37691 3587
rect 38301 3553 38335 3587
rect 40233 3553 40267 3587
rect 41889 3553 41923 3587
rect 44097 3553 44131 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 2881 3485 2915 3519
rect 3985 3485 4019 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 12081 3485 12115 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 17601 3485 17635 3519
rect 18245 3485 18279 3519
rect 19533 3485 19567 3519
rect 20177 3485 20211 3519
rect 22477 3485 22511 3519
rect 23121 3485 23155 3519
rect 24685 3485 24719 3519
rect 27261 3485 27295 3519
rect 32965 3485 32999 3519
rect 33793 3485 33827 3519
rect 39957 3485 39991 3519
rect 40969 3485 41003 3519
rect 43269 3485 43303 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 1869 3417 1903 3451
rect 6745 3417 6779 3451
rect 20361 3417 20395 3451
rect 25706 3417 25740 3451
rect 37749 3417 37783 3451
rect 41153 3417 41187 3451
rect 48145 3417 48179 3451
rect 2145 3349 2179 3383
rect 12173 3349 12207 3383
rect 14197 3349 14231 3383
rect 18337 3349 18371 3383
rect 24777 3349 24811 3383
rect 27077 3349 27111 3383
rect 33057 3349 33091 3383
rect 40509 3349 40543 3383
rect 43361 3349 43395 3383
rect 45753 3349 45787 3383
rect 6745 3145 6779 3179
rect 18337 3145 18371 3179
rect 18981 3145 19015 3179
rect 37749 3145 37783 3179
rect 39773 3145 39807 3179
rect 41061 3145 41095 3179
rect 47869 3145 47903 3179
rect 1961 3077 1995 3111
rect 8125 3077 8159 3111
rect 11713 3077 11747 3111
rect 14013 3077 14047 3111
rect 21189 3077 21223 3111
rect 24777 3077 24811 3111
rect 33149 3077 33183 3111
rect 42993 3077 43027 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 6653 3009 6687 3043
rect 7941 3009 7975 3043
rect 11529 3009 11563 3043
rect 13829 3009 13863 3043
rect 17417 3009 17451 3043
rect 18245 3009 18279 3043
rect 18889 3009 18923 3043
rect 19533 3009 19567 3043
rect 20361 3009 20395 3043
rect 21097 3009 21131 3043
rect 22385 3009 22419 3043
rect 23121 3009 23155 3043
rect 23765 3009 23799 3043
rect 24593 3009 24627 3043
rect 27169 3009 27203 3043
rect 32965 3009 32999 3043
rect 37289 3009 37323 3043
rect 39957 3009 39991 3043
rect 40417 3009 40451 3043
rect 42809 3009 42843 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 8401 2941 8435 2975
rect 11989 2941 12023 2975
rect 14289 2941 14323 2975
rect 17325 2941 17359 2975
rect 17785 2941 17819 2975
rect 23029 2941 23063 2975
rect 25145 2941 25179 2975
rect 33517 2941 33551 2975
rect 40601 2941 40635 2975
rect 43269 2941 43303 2975
rect 47041 2941 47075 2975
rect 19625 2805 19659 2839
rect 23857 2805 23891 2839
rect 27353 2805 27387 2839
rect 37381 2805 37415 2839
rect 19993 2601 20027 2635
rect 20913 2601 20947 2635
rect 22385 2601 22419 2635
rect 23029 2601 23063 2635
rect 25973 2601 26007 2635
rect 28641 2601 28675 2635
rect 36369 2601 36403 2635
rect 39129 2601 39163 2635
rect 41705 2601 41739 2635
rect 42533 2601 42567 2635
rect 42901 2601 42935 2635
rect 19349 2533 19383 2567
rect 26157 2533 26191 2567
rect 38301 2533 38335 2567
rect 41245 2533 41279 2567
rect 1409 2465 1443 2499
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 7021 2465 7055 2499
rect 15853 2465 15887 2499
rect 27261 2465 27295 2499
rect 40509 2465 40543 2499
rect 46489 2465 46523 2499
rect 47869 2465 47903 2499
rect 4997 2397 5031 2431
rect 6561 2397 6595 2431
rect 16681 2397 16715 2431
rect 19257 2397 19291 2431
rect 19901 2397 19935 2431
rect 20729 2397 20763 2431
rect 22937 2397 22971 2431
rect 23581 2397 23615 2431
rect 25697 2397 25731 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 29929 2397 29963 2431
rect 35725 2397 35759 2431
rect 38117 2397 38151 2431
rect 39313 2397 39347 2431
rect 41889 2397 41923 2431
rect 42441 2397 42475 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46213 2397 46247 2431
rect 47685 2397 47719 2431
rect 1593 2329 1627 2363
rect 4169 2329 4203 2363
rect 6745 2329 6779 2363
rect 9413 2329 9447 2363
rect 15669 2329 15703 2363
rect 22293 2329 22327 2363
rect 24869 2329 24903 2363
rect 36277 2329 36311 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 45385 2329 45419 2363
rect 4445 2261 4479 2295
rect 9689 2261 9723 2295
rect 16865 2261 16899 2295
rect 23673 2261 23707 2295
rect 24961 2261 24995 2295
rect 29745 2261 29779 2295
rect 35541 2261 35575 2295
rect 45477 2261 45511 2295
<< metal1 >>
rect 45554 47880 45560 47932
rect 45612 47920 45618 47932
rect 46106 47920 46112 47932
rect 45612 47892 46112 47920
rect 45612 47880 45618 47892
rect 46106 47880 46112 47892
rect 46164 47880 46170 47932
rect 40034 47404 40040 47456
rect 40092 47444 40098 47456
rect 41230 47444 41236 47456
rect 40092 47416 41236 47444
rect 40092 47404 40098 47416
rect 41230 47404 41236 47416
rect 41288 47404 41294 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 13357 47243 13415 47249
rect 13357 47209 13369 47243
rect 13403 47240 13415 47243
rect 21910 47240 21916 47252
rect 13403 47212 21916 47240
rect 13403 47209 13415 47212
rect 13357 47203 13415 47209
rect 21910 47200 21916 47212
rect 21968 47200 21974 47252
rect 36906 47200 36912 47252
rect 36964 47240 36970 47252
rect 46842 47240 46848 47252
rect 36964 47212 46848 47240
rect 36964 47200 36970 47212
rect 46842 47200 46848 47212
rect 46900 47200 46906 47252
rect 20530 47132 20536 47184
rect 20588 47172 20594 47184
rect 21821 47175 21879 47181
rect 21821 47172 21833 47175
rect 20588 47144 21833 47172
rect 20588 47132 20594 47144
rect 21821 47141 21833 47144
rect 21867 47141 21879 47175
rect 21821 47135 21879 47141
rect 28629 47175 28687 47181
rect 28629 47141 28641 47175
rect 28675 47172 28687 47175
rect 28902 47172 28908 47184
rect 28675 47144 28908 47172
rect 28675 47141 28687 47144
rect 28629 47135 28687 47141
rect 28902 47132 28908 47144
rect 28960 47132 28966 47184
rect 35342 47132 35348 47184
rect 35400 47172 35406 47184
rect 43855 47175 43913 47181
rect 43855 47172 43867 47175
rect 35400 47144 43867 47172
rect 35400 47132 35406 47144
rect 43855 47141 43867 47144
rect 43901 47141 43913 47175
rect 43855 47135 43913 47141
rect 44450 47132 44456 47184
rect 44508 47132 44514 47184
rect 47762 47132 47768 47184
rect 47820 47172 47826 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 47820 47144 47961 47172
rect 47820 47132 47826 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 6641 47107 6699 47113
rect 6641 47073 6653 47107
rect 6687 47104 6699 47107
rect 30742 47104 30748 47116
rect 6687 47076 30604 47104
rect 30703 47076 30748 47104
rect 6687 47073 6699 47076
rect 6641 47067 6699 47073
rect 1765 47039 1823 47045
rect 1765 47005 1777 47039
rect 1811 47036 1823 47039
rect 1946 47036 1952 47048
rect 1811 47008 1952 47036
rect 1811 47005 1823 47008
rect 1765 46999 1823 47005
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4798 47036 4804 47048
rect 4759 47008 4804 47036
rect 3789 46999 3847 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 5868 47008 6377 47036
rect 5868 46996 5874 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7374 47036 7380 47048
rect 7335 47008 7380 47036
rect 6365 46999 6423 47005
rect 7374 46996 7380 47008
rect 7432 46996 7438 47048
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 11606 47036 11612 47048
rect 11567 47008 11612 47036
rect 9401 46999 9459 47005
rect 11606 46996 11612 47008
rect 11664 46996 11670 47048
rect 12250 46996 12256 47048
rect 12308 47036 12314 47048
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 12308 47008 12357 47036
rect 12308 46996 12314 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12345 46999 12403 47005
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 14093 47039 14151 47045
rect 14093 47036 14105 47039
rect 13872 47008 14105 47036
rect 13872 46996 13878 47008
rect 14093 47005 14105 47008
rect 14139 47005 14151 47039
rect 14366 47036 14372 47048
rect 14327 47008 14372 47036
rect 14093 46999 14151 47005
rect 14366 46996 14372 47008
rect 14424 46996 14430 47048
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 16945 47039 17003 47045
rect 16945 47005 16957 47039
rect 16991 47036 17003 47039
rect 17770 47036 17776 47048
rect 16991 47008 17776 47036
rect 16991 47005 17003 47008
rect 16945 46999 17003 47005
rect 17770 46996 17776 47008
rect 17828 46996 17834 47048
rect 20990 47036 20996 47048
rect 20951 47008 20996 47036
rect 20990 46996 20996 47008
rect 21048 46996 21054 47048
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21100 47008 22017 47036
rect 2041 46971 2099 46977
rect 2041 46937 2053 46971
rect 2087 46968 2099 46971
rect 2498 46968 2504 46980
rect 2087 46940 2504 46968
rect 2087 46937 2099 46940
rect 2041 46931 2099 46937
rect 2498 46928 2504 46940
rect 2556 46928 2562 46980
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 2777 46931 2835 46937
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 2792 46900 2820 46931
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 7466 46928 7472 46980
rect 7524 46968 7530 46980
rect 7561 46971 7619 46977
rect 7561 46968 7573 46971
rect 7524 46940 7573 46968
rect 7524 46928 7530 46940
rect 7561 46937 7573 46940
rect 7607 46937 7619 46971
rect 7561 46931 7619 46937
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 11698 46928 11704 46980
rect 11756 46968 11762 46980
rect 11793 46971 11851 46977
rect 11793 46968 11805 46971
rect 11756 46940 11805 46968
rect 11756 46928 11762 46940
rect 11793 46937 11805 46940
rect 11839 46937 11851 46971
rect 11793 46931 11851 46937
rect 12434 46928 12440 46980
rect 12492 46968 12498 46980
rect 12529 46971 12587 46977
rect 12529 46968 12541 46971
rect 12492 46940 12541 46968
rect 12492 46928 12498 46940
rect 12529 46937 12541 46940
rect 12575 46937 12587 46971
rect 12529 46931 12587 46937
rect 19705 46971 19763 46977
rect 19705 46937 19717 46971
rect 19751 46937 19763 46971
rect 19705 46931 19763 46937
rect 20073 46971 20131 46977
rect 20073 46937 20085 46971
rect 20119 46968 20131 46971
rect 20622 46968 20628 46980
rect 20119 46940 20628 46968
rect 20119 46937 20131 46940
rect 20073 46931 20131 46937
rect 2648 46872 2820 46900
rect 2648 46860 2654 46872
rect 2866 46860 2872 46912
rect 2924 46900 2930 46912
rect 4890 46900 4896 46912
rect 2924 46872 2969 46900
rect 4851 46872 4896 46900
rect 2924 46860 2930 46872
rect 4890 46860 4896 46872
rect 4948 46860 4954 46912
rect 18690 46860 18696 46912
rect 18748 46900 18754 46912
rect 19720 46900 19748 46931
rect 20622 46928 20628 46940
rect 20680 46928 20686 46980
rect 18748 46872 19748 46900
rect 18748 46860 18754 46872
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 21100 46900 21128 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 24578 46996 24584 47048
rect 24636 47036 24642 47048
rect 24765 47039 24823 47045
rect 24765 47036 24777 47039
rect 24636 47008 24777 47036
rect 24636 46996 24642 47008
rect 24765 47005 24777 47008
rect 24811 47005 24823 47039
rect 25406 47036 25412 47048
rect 25367 47008 25412 47036
rect 24765 46999 24823 47005
rect 25406 46996 25412 47008
rect 25464 46996 25470 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28445 47039 28503 47045
rect 28445 47036 28457 47039
rect 28408 47008 28457 47036
rect 28408 46996 28414 47008
rect 28445 47005 28457 47008
rect 28491 47005 28503 47039
rect 28445 46999 28503 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 30009 47039 30067 47045
rect 30009 47036 30021 47039
rect 29696 47008 30021 47036
rect 29696 46996 29702 47008
rect 30009 47005 30021 47008
rect 30055 47005 30067 47039
rect 30009 46999 30067 47005
rect 29362 46928 29368 46980
rect 29420 46968 29426 46980
rect 30193 46971 30251 46977
rect 30193 46968 30205 46971
rect 29420 46940 30205 46968
rect 29420 46928 29426 46940
rect 30193 46937 30205 46940
rect 30239 46937 30251 46971
rect 30576 46968 30604 47076
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 39298 47064 39304 47116
rect 39356 47104 39362 47116
rect 39853 47107 39911 47113
rect 39853 47104 39865 47107
rect 39356 47076 39865 47104
rect 39356 47064 39362 47076
rect 39853 47073 39865 47076
rect 39899 47073 39911 47107
rect 39853 47067 39911 47073
rect 43625 47107 43683 47113
rect 43625 47073 43637 47107
rect 43671 47104 43683 47107
rect 44468 47104 44496 47132
rect 43671 47076 44496 47104
rect 47029 47107 47087 47113
rect 43671 47073 43683 47076
rect 43625 47067 43683 47073
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 31021 47039 31079 47045
rect 31021 47005 31033 47039
rect 31067 47036 31079 47039
rect 34698 47036 34704 47048
rect 31067 47008 34704 47036
rect 31067 47005 31079 47008
rect 31021 46999 31079 47005
rect 34698 46996 34704 47008
rect 34756 46996 34762 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 40129 47039 40187 47045
rect 40129 47036 40141 47039
rect 38381 46999 38439 47005
rect 39316 47008 40141 47036
rect 39316 46980 39344 47008
rect 40129 47005 40141 47008
rect 40175 47005 40187 47039
rect 41874 47036 41880 47048
rect 41835 47008 41880 47036
rect 40129 46999 40187 47005
rect 41874 46996 41880 47008
rect 41932 46996 41938 47048
rect 42981 47039 43039 47045
rect 42981 47005 42993 47039
rect 43027 47036 43039 47039
rect 43806 47036 43812 47048
rect 43027 47008 43812 47036
rect 43027 47005 43039 47008
rect 42981 46999 43039 47005
rect 43806 46996 43812 47008
rect 43864 46996 43870 47048
rect 44450 46996 44456 47048
rect 44508 47036 44514 47048
rect 45189 47039 45247 47045
rect 45189 47036 45201 47039
rect 44508 47008 45201 47036
rect 44508 46996 44514 47008
rect 45189 47005 45201 47008
rect 45235 47005 45247 47039
rect 45189 46999 45247 47005
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 37366 46968 37372 46980
rect 30576 46940 37372 46968
rect 30193 46931 30251 46937
rect 37366 46928 37372 46940
rect 37424 46928 37430 46980
rect 39298 46928 39304 46980
rect 39356 46928 39362 46980
rect 43070 46928 43076 46980
rect 43128 46968 43134 46980
rect 43165 46971 43223 46977
rect 43165 46968 43177 46971
rect 43128 46940 43177 46968
rect 43128 46928 43134 46940
rect 43165 46937 43177 46940
rect 43211 46937 43223 46971
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 43165 46931 43223 46937
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 20036 46872 21128 46900
rect 20036 46860 20042 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 3878 46588 3884 46640
rect 3936 46628 3942 46640
rect 3936 46600 33548 46628
rect 3936 46588 3942 46600
rect 24578 46560 24584 46572
rect 24539 46532 24584 46560
rect 24578 46520 24584 46532
rect 24636 46520 24642 46572
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46492 11759 46495
rect 12066 46492 12072 46504
rect 11747 46464 12072 46492
rect 11747 46461 11759 46464
rect 11701 46455 11759 46461
rect 12066 46452 12072 46464
rect 12124 46452 12130 46504
rect 12161 46495 12219 46501
rect 12161 46461 12173 46495
rect 12207 46461 12219 46495
rect 12161 46455 12219 46461
rect 12176 46424 12204 46455
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13817 46495 13875 46501
rect 13817 46492 13829 46495
rect 13596 46464 13829 46492
rect 13596 46452 13602 46464
rect 13817 46461 13829 46464
rect 13863 46461 13875 46495
rect 13817 46455 13875 46461
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46492 14059 46495
rect 14182 46492 14188 46504
rect 14047 46464 14188 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19242 46492 19248 46504
rect 14332 46464 14377 46492
rect 19203 46464 19248 46492
rect 14332 46452 14338 46464
rect 19242 46452 19248 46464
rect 19300 46452 19306 46504
rect 19429 46495 19487 46501
rect 19429 46461 19441 46495
rect 19475 46461 19487 46495
rect 20438 46492 20444 46504
rect 20399 46464 20444 46492
rect 19429 46455 19487 46461
rect 10980 46396 12204 46424
rect 10980 46368 11008 46396
rect 18598 46384 18604 46436
rect 18656 46424 18662 46436
rect 19444 46424 19472 46455
rect 20438 46452 20444 46464
rect 20496 46452 20502 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 32585 46455 32643 46461
rect 18656 46396 19472 46424
rect 18656 46384 18662 46396
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 32272 46396 32628 46424
rect 33520 46424 33548 46600
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47946 46560 47952 46572
rect 47907 46532 47952 46560
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 34422 46492 34428 46504
rect 34383 46464 34428 46492
rect 34422 46452 34428 46464
rect 34480 46452 34486 46504
rect 34609 46495 34667 46501
rect 34609 46461 34621 46495
rect 34655 46492 34667 46495
rect 34790 46492 34796 46504
rect 34655 46464 34796 46492
rect 34655 46461 34667 46464
rect 34609 46455 34667 46461
rect 34790 46452 34796 46464
rect 34848 46452 34854 46504
rect 34885 46495 34943 46501
rect 34885 46461 34897 46495
rect 34931 46461 34943 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 34885 46455 34943 46461
rect 34900 46424 34928 46455
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 45186 46492 45192 46504
rect 45147 46464 45192 46492
rect 42889 46455 42947 46461
rect 33520 46396 34928 46424
rect 32272 46384 32278 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 45186 46452 45192 46464
rect 45244 46452 45250 46504
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46750 46492 46756 46504
rect 45419 46464 45554 46492
rect 46711 46464 46756 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 42576 46396 42932 46424
rect 45526 46424 45554 46464
rect 46750 46452 46756 46464
rect 46808 46452 46814 46504
rect 46658 46424 46664 46436
rect 45526 46396 46664 46424
rect 42576 46384 42582 46396
rect 46658 46384 46664 46396
rect 46716 46384 46722 46436
rect 2133 46359 2191 46365
rect 2133 46325 2145 46359
rect 2179 46356 2191 46359
rect 2314 46356 2320 46368
rect 2179 46328 2320 46356
rect 2179 46325 2191 46328
rect 2133 46319 2191 46325
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 2406 46316 2412 46368
rect 2464 46356 2470 46368
rect 2869 46359 2927 46365
rect 2869 46356 2881 46359
rect 2464 46328 2881 46356
rect 2464 46316 2470 46328
rect 2869 46325 2881 46328
rect 2915 46325 2927 46359
rect 2869 46319 2927 46325
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 38654 46316 38660 46368
rect 38712 46356 38718 46368
rect 39942 46356 39948 46368
rect 38712 46328 39948 46356
rect 38712 46316 38718 46328
rect 39942 46316 39948 46328
rect 40000 46316 40006 46368
rect 41230 46356 41236 46368
rect 41191 46328 41236 46356
rect 41230 46316 41236 46328
rect 41288 46316 41294 46368
rect 47302 46316 47308 46368
rect 47360 46356 47366 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47360 46328 48053 46356
rect 47360 46316 47366 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 12066 46152 12072 46164
rect 12027 46124 12072 46152
rect 12066 46112 12072 46124
rect 12124 46112 12130 46164
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 18598 46152 18604 46164
rect 18559 46124 18604 46152
rect 18598 46112 18604 46124
rect 18656 46112 18662 46164
rect 19242 46112 19248 46164
rect 19300 46152 19306 46164
rect 19429 46155 19487 46161
rect 19429 46152 19441 46155
rect 19300 46124 19441 46152
rect 19300 46112 19306 46124
rect 19429 46121 19441 46124
rect 19475 46121 19487 46155
rect 19429 46115 19487 46121
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 32033 46155 32091 46161
rect 32033 46121 32045 46155
rect 32079 46152 32091 46155
rect 32306 46152 32312 46164
rect 32079 46124 32312 46152
rect 32079 46121 32091 46124
rect 32033 46115 32091 46121
rect 32306 46112 32312 46124
rect 32364 46112 32370 46164
rect 33597 46155 33655 46161
rect 33597 46121 33609 46155
rect 33643 46152 33655 46155
rect 34422 46152 34428 46164
rect 33643 46124 34428 46152
rect 33643 46121 33655 46124
rect 33597 46115 33655 46121
rect 34422 46112 34428 46124
rect 34480 46112 34486 46164
rect 34790 46152 34796 46164
rect 34751 46124 34796 46152
rect 34790 46112 34796 46124
rect 34848 46112 34854 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 43809 46155 43867 46161
rect 43809 46121 43821 46155
rect 43855 46152 43867 46155
rect 45186 46152 45192 46164
rect 43855 46124 45192 46152
rect 43855 46121 43867 46124
rect 43809 46115 43867 46121
rect 45186 46112 45192 46124
rect 45244 46112 45250 46164
rect 38212 46056 42656 46084
rect 1397 46019 1455 46025
rect 1397 45985 1409 46019
rect 1443 46016 1455 46019
rect 2406 46016 2412 46028
rect 1443 45988 2412 46016
rect 1443 45985 1455 45988
rect 1397 45979 1455 45985
rect 2406 45976 2412 45988
rect 2464 45976 2470 46028
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 20717 46019 20775 46025
rect 20717 45985 20729 46019
rect 20763 46016 20775 46019
rect 20990 46016 20996 46028
rect 20763 45988 20996 46016
rect 20763 45985 20775 45988
rect 20717 45979 20775 45985
rect 20990 45976 20996 45988
rect 21048 45976 21054 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25406 46016 25412 46028
rect 25271 45988 25412 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25406 45976 25412 45988
rect 25464 45976 25470 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 11974 45948 11980 45960
rect 11935 45920 11980 45948
rect 11974 45908 11980 45920
rect 12032 45908 12038 45960
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 18509 45951 18567 45957
rect 18509 45948 18521 45951
rect 14148 45920 18521 45948
rect 14148 45908 14154 45920
rect 18509 45917 18521 45920
rect 18555 45948 18567 45951
rect 18690 45948 18696 45960
rect 18555 45920 18696 45948
rect 18555 45917 18567 45920
rect 18509 45911 18567 45917
rect 18690 45908 18696 45920
rect 18748 45908 18754 45960
rect 24578 45948 24584 45960
rect 24539 45920 24584 45948
rect 24578 45908 24584 45920
rect 24636 45908 24642 45960
rect 31941 45951 31999 45957
rect 31941 45917 31953 45951
rect 31987 45948 31999 45951
rect 32582 45948 32588 45960
rect 31987 45920 32588 45948
rect 31987 45917 31999 45920
rect 31941 45911 31999 45917
rect 32582 45908 32588 45920
rect 32640 45908 32646 45960
rect 34701 45951 34759 45957
rect 34701 45917 34713 45951
rect 34747 45948 34759 45951
rect 35434 45948 35440 45960
rect 34747 45920 35440 45948
rect 34747 45917 34759 45920
rect 34701 45911 34759 45917
rect 35434 45908 35440 45920
rect 35492 45948 35498 45960
rect 38212 45957 38240 46056
rect 41230 46016 41236 46028
rect 41191 45988 41236 46016
rect 41230 45976 41236 45988
rect 41288 45976 41294 46028
rect 41966 46016 41972 46028
rect 41927 45988 41972 46016
rect 41966 45976 41972 45988
rect 42024 45976 42030 46028
rect 38197 45951 38255 45957
rect 38197 45948 38209 45951
rect 35492 45920 38209 45948
rect 35492 45908 35498 45920
rect 38197 45917 38209 45920
rect 38243 45917 38255 45951
rect 42628 45948 42656 46056
rect 45094 46044 45100 46096
rect 45152 46084 45158 46096
rect 45646 46084 45652 46096
rect 45152 46056 45652 46084
rect 45152 46044 45158 46056
rect 45646 46044 45652 46056
rect 45704 46044 45710 46096
rect 44453 46019 44511 46025
rect 44453 45985 44465 46019
rect 44499 46016 44511 46019
rect 46293 46019 46351 46025
rect 46293 46016 46305 46019
rect 44499 45988 46305 46016
rect 44499 45985 44511 45988
rect 44453 45979 44511 45985
rect 46293 45985 46305 45988
rect 46339 45985 46351 46019
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 46293 45979 46351 45985
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 45649 45951 45707 45957
rect 42628 45920 45554 45948
rect 38197 45911 38255 45917
rect 1581 45883 1639 45889
rect 1581 45849 1593 45883
rect 1627 45880 1639 45883
rect 2222 45880 2228 45892
rect 1627 45852 2228 45880
rect 1627 45849 1639 45852
rect 1581 45843 1639 45849
rect 2222 45840 2228 45852
rect 2280 45840 2286 45892
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 41414 45880 41420 45892
rect 41375 45852 41420 45880
rect 41414 45840 41420 45852
rect 41472 45840 41478 45892
rect 45526 45880 45554 45920
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 46290 45880 46296 45892
rect 45526 45852 46296 45880
rect 46290 45840 46296 45852
rect 46348 45840 46354 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 26878 45772 26884 45824
rect 26936 45812 26942 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 26936 45784 45753 45812
rect 26936 45772 26942 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 2222 45608 2228 45620
rect 2183 45580 2228 45608
rect 2222 45568 2228 45580
rect 2280 45568 2286 45620
rect 11974 45568 11980 45620
rect 12032 45608 12038 45620
rect 20898 45608 20904 45620
rect 12032 45580 20760 45608
rect 20859 45580 20904 45608
rect 12032 45568 12038 45580
rect 1946 45432 1952 45484
rect 2004 45472 2010 45484
rect 2133 45475 2191 45481
rect 2133 45472 2145 45475
rect 2004 45444 2145 45472
rect 2004 45432 2010 45444
rect 2133 45441 2145 45444
rect 2179 45472 2191 45475
rect 20732 45472 20760 45580
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 24578 45568 24584 45620
rect 24636 45608 24642 45620
rect 36170 45608 36176 45620
rect 24636 45580 36176 45608
rect 24636 45568 24642 45580
rect 36170 45568 36176 45580
rect 36228 45568 36234 45620
rect 41785 45611 41843 45617
rect 41785 45577 41797 45611
rect 41831 45608 41843 45611
rect 42610 45608 42616 45620
rect 41831 45580 42616 45608
rect 41831 45577 41843 45580
rect 41785 45571 41843 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45554 45568 45560 45620
rect 45612 45608 45618 45620
rect 45612 45580 47992 45608
rect 45612 45568 45618 45580
rect 25406 45540 25412 45552
rect 25367 45512 25412 45540
rect 25406 45500 25412 45512
rect 25464 45500 25470 45552
rect 41141 45543 41199 45549
rect 41141 45509 41153 45543
rect 41187 45540 41199 45543
rect 41414 45540 41420 45552
rect 41187 45512 41420 45540
rect 41187 45509 41199 45512
rect 41141 45503 41199 45509
rect 41414 45500 41420 45512
rect 41472 45500 41478 45552
rect 47964 45549 47992 45580
rect 47949 45543 48007 45549
rect 47949 45509 47961 45543
rect 47995 45509 48007 45543
rect 47949 45503 48007 45509
rect 20809 45475 20867 45481
rect 20809 45472 20821 45475
rect 2179 45444 6914 45472
rect 2179 45441 2191 45444
rect 2133 45435 2191 45441
rect 6886 45336 6914 45444
rect 20732 45444 20821 45472
rect 20732 45404 20760 45444
rect 20809 45441 20821 45444
rect 20855 45441 20867 45475
rect 20809 45435 20867 45441
rect 25317 45475 25375 45481
rect 25317 45441 25329 45475
rect 25363 45472 25375 45475
rect 25774 45472 25780 45484
rect 25363 45444 25780 45472
rect 25363 45441 25375 45444
rect 25317 45435 25375 45441
rect 25774 45432 25780 45444
rect 25832 45432 25838 45484
rect 41046 45472 41052 45484
rect 41007 45444 41052 45472
rect 41046 45432 41052 45444
rect 41104 45432 41110 45484
rect 41693 45475 41751 45481
rect 41693 45441 41705 45475
rect 41739 45441 41751 45475
rect 41693 45435 41751 45441
rect 32582 45404 32588 45416
rect 20732 45376 32588 45404
rect 32582 45364 32588 45376
rect 32640 45364 32646 45416
rect 24578 45336 24584 45348
rect 6886 45308 24584 45336
rect 24578 45296 24584 45308
rect 24636 45296 24642 45348
rect 41708 45336 41736 45435
rect 41874 45432 41880 45484
rect 41932 45472 41938 45484
rect 42705 45475 42763 45481
rect 42705 45472 42717 45475
rect 41932 45444 42717 45472
rect 41932 45432 41938 45444
rect 42705 45441 42717 45444
rect 42751 45441 42763 45475
rect 42705 45435 42763 45441
rect 42886 45404 42892 45416
rect 42847 45376 42892 45404
rect 42886 45364 42892 45376
rect 42944 45364 42950 45416
rect 44082 45404 44088 45416
rect 44043 45376 44088 45404
rect 44082 45364 44088 45376
rect 44140 45364 44146 45416
rect 44910 45364 44916 45416
rect 44968 45404 44974 45416
rect 45005 45407 45063 45413
rect 45005 45404 45017 45407
rect 44968 45376 45017 45404
rect 44968 45364 44974 45376
rect 45005 45373 45017 45376
rect 45051 45373 45063 45407
rect 45186 45404 45192 45416
rect 45147 45376 45192 45404
rect 45005 45367 45063 45373
rect 45186 45364 45192 45376
rect 45244 45364 45250 45416
rect 45738 45404 45744 45416
rect 45699 45376 45744 45404
rect 45738 45364 45744 45376
rect 45796 45364 45802 45416
rect 46842 45336 46848 45348
rect 41708 45308 46848 45336
rect 46842 45296 46848 45308
rect 46900 45296 46906 45348
rect 48038 45268 48044 45280
rect 47999 45240 48044 45268
rect 48038 45228 48044 45240
rect 48096 45228 48102 45280
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 42886 45064 42892 45076
rect 42847 45036 42892 45064
rect 42886 45024 42892 45036
rect 42944 45024 42950 45076
rect 44450 45064 44456 45076
rect 44411 45036 44456 45064
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45097 45067 45155 45073
rect 45097 45033 45109 45067
rect 45143 45064 45155 45067
rect 45186 45064 45192 45076
rect 45143 45036 45192 45064
rect 45143 45033 45155 45036
rect 45097 45027 45155 45033
rect 45186 45024 45192 45036
rect 45244 45024 45250 45076
rect 45370 45024 45376 45076
rect 45428 45064 45434 45076
rect 45741 45067 45799 45073
rect 45741 45064 45753 45067
rect 45428 45036 45753 45064
rect 45428 45024 45434 45036
rect 45741 45033 45753 45036
rect 45787 45033 45799 45067
rect 45741 45027 45799 45033
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 42797 44863 42855 44869
rect 42797 44829 42809 44863
rect 42843 44829 42855 44863
rect 42797 44823 42855 44829
rect 45005 44863 45063 44869
rect 45005 44829 45017 44863
rect 45051 44860 45063 44863
rect 45554 44860 45560 44872
rect 45051 44832 45560 44860
rect 45051 44829 45063 44832
rect 45005 44823 45063 44829
rect 42812 44724 42840 44823
rect 45554 44820 45560 44832
rect 45612 44820 45618 44872
rect 45649 44863 45707 44869
rect 45649 44829 45661 44863
rect 45695 44860 45707 44863
rect 45738 44860 45744 44872
rect 45695 44832 45744 44860
rect 45695 44829 45707 44832
rect 45649 44823 45707 44829
rect 45738 44820 45744 44832
rect 45796 44820 45802 44872
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 47854 44724 47860 44736
rect 42812 44696 47860 44724
rect 47854 44684 47860 44696
rect 47912 44684 47918 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 46385 44523 46443 44529
rect 46385 44489 46397 44523
rect 46431 44520 46443 44523
rect 46474 44520 46480 44532
rect 46431 44492 46480 44520
rect 46431 44489 46443 44492
rect 46385 44483 46443 44489
rect 46474 44480 46480 44492
rect 46532 44480 46538 44532
rect 46658 44480 46664 44532
rect 46716 44520 46722 44532
rect 47673 44523 47731 44529
rect 47673 44520 47685 44523
rect 46716 44492 47685 44520
rect 46716 44480 46722 44492
rect 47673 44489 47685 44492
rect 47719 44489 47731 44523
rect 47673 44483 47731 44489
rect 44910 44384 44916 44396
rect 44871 44356 44916 44384
rect 44910 44344 44916 44356
rect 44968 44344 44974 44396
rect 45649 44387 45707 44393
rect 45649 44353 45661 44387
rect 45695 44353 45707 44387
rect 46290 44384 46296 44396
rect 46251 44356 46296 44384
rect 45649 44347 45707 44353
rect 45664 44316 45692 44347
rect 46290 44344 46296 44356
rect 46348 44344 46354 44396
rect 47486 44344 47492 44396
rect 47544 44384 47550 44396
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 47544 44356 47593 44384
rect 47544 44344 47550 44356
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 47394 44316 47400 44328
rect 45664 44288 47400 44316
rect 47394 44276 47400 44288
rect 47452 44276 47458 44328
rect 41046 44208 41052 44260
rect 41104 44248 41110 44260
rect 47578 44248 47584 44260
rect 41104 44220 47584 44248
rect 41104 44208 41110 44220
rect 47578 44208 47584 44220
rect 47636 44208 47642 44260
rect 45741 44183 45799 44189
rect 45741 44149 45753 44183
rect 45787 44180 45799 44183
rect 46474 44180 46480 44192
rect 45787 44152 46480 44180
rect 45787 44149 45799 44152
rect 45741 44143 45799 44149
rect 46474 44140 46480 44152
rect 46532 44140 46538 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46474 43840 46480 43852
rect 46435 43812 46480 43840
rect 46474 43800 46480 43812
rect 46532 43800 46538 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 47670 43432 47676 43444
rect 47631 43404 47676 43432
rect 47670 43392 47676 43404
rect 47728 43392 47734 43444
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47394 43256 47400 43308
rect 47452 43296 47458 43308
rect 47581 43299 47639 43305
rect 47581 43296 47593 43299
rect 47452 43268 47593 43296
rect 47452 43256 47458 43268
rect 47581 43265 47593 43268
rect 47627 43265 47639 43299
rect 47581 43259 47639 43265
rect 1486 43188 1492 43240
rect 1544 43228 1550 43240
rect 1581 43231 1639 43237
rect 1581 43228 1593 43231
rect 1544 43200 1593 43228
rect 1544 43188 1550 43200
rect 1581 43197 1593 43200
rect 1627 43197 1639 43231
rect 1581 43191 1639 43197
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47029 42171 47087 42177
rect 47581 42211 47639 42217
rect 47581 42177 47593 42211
rect 47627 42208 47639 42211
rect 47854 42208 47860 42220
rect 47627 42180 47860 42208
rect 47627 42177 47639 42180
rect 47581 42171 47639 42177
rect 47854 42168 47860 42180
rect 47912 42168 47918 42220
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46845 41259 46903 41265
rect 46845 41256 46857 41259
rect 46532 41228 46857 41256
rect 46532 41216 46538 41228
rect 46845 41225 46857 41228
rect 46891 41225 46903 41259
rect 46845 41219 46903 41225
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 46753 41123 46811 41129
rect 46753 41089 46765 41123
rect 46799 41120 46811 41123
rect 46842 41120 46848 41132
rect 46799 41092 46848 41120
rect 46799 41089 46811 41092
rect 46753 41083 46811 41089
rect 46842 41080 46848 41092
rect 46900 41080 46906 41132
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 45526 40956 48145 40984
rect 39206 40876 39212 40928
rect 39264 40916 39270 40928
rect 45526 40916 45554 40956
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 39264 40888 45554 40916
rect 39264 40876 39270 40888
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 26881 40579 26939 40585
rect 26881 40545 26893 40579
rect 26927 40576 26939 40579
rect 26970 40576 26976 40588
rect 26927 40548 26976 40576
rect 26927 40545 26939 40548
rect 26881 40539 26939 40545
rect 26970 40536 26976 40548
rect 27028 40536 27034 40588
rect 26602 40468 26608 40520
rect 26660 40508 26666 40520
rect 26697 40511 26755 40517
rect 26697 40508 26709 40511
rect 26660 40480 26709 40508
rect 26660 40468 26666 40480
rect 26697 40477 26709 40480
rect 26743 40477 26755 40511
rect 47026 40508 47032 40520
rect 46987 40480 47032 40508
rect 26697 40471 26755 40477
rect 47026 40468 47032 40480
rect 47084 40468 47090 40520
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2038 40440 2044 40452
rect 1999 40412 2044 40440
rect 2038 40400 2044 40412
rect 2096 40400 2102 40452
rect 26234 40372 26240 40384
rect 26195 40344 26240 40372
rect 26234 40332 26240 40344
rect 26292 40332 26298 40384
rect 26605 40375 26663 40381
rect 26605 40341 26617 40375
rect 26651 40372 26663 40375
rect 26878 40372 26884 40384
rect 26651 40344 26884 40372
rect 26651 40341 26663 40344
rect 26605 40335 26663 40341
rect 26878 40332 26884 40344
rect 26936 40332 26942 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 25869 40171 25927 40177
rect 25869 40137 25881 40171
rect 25915 40168 25927 40171
rect 26418 40168 26424 40180
rect 25915 40140 26424 40168
rect 25915 40137 25927 40140
rect 25869 40131 25927 40137
rect 26418 40128 26424 40140
rect 26476 40128 26482 40180
rect 23474 40060 23480 40112
rect 23532 40100 23538 40112
rect 23532 40072 24886 40100
rect 23532 40060 23538 40072
rect 19242 39992 19248 40044
rect 19300 40032 19306 40044
rect 19889 40035 19947 40041
rect 19889 40032 19901 40035
rect 19300 40004 19901 40032
rect 19300 39992 19306 40004
rect 19889 40001 19901 40004
rect 19935 40001 19947 40035
rect 47578 40032 47584 40044
rect 47539 40004 47584 40032
rect 19889 39995 19947 40001
rect 47578 39992 47584 40004
rect 47636 39992 47642 40044
rect 23842 39924 23848 39976
rect 23900 39964 23906 39976
rect 24121 39967 24179 39973
rect 24121 39964 24133 39967
rect 23900 39936 24133 39964
rect 23900 39924 23906 39936
rect 24121 39933 24133 39936
rect 24167 39933 24179 39967
rect 24121 39927 24179 39933
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39964 24455 39967
rect 25130 39964 25136 39976
rect 24443 39936 25136 39964
rect 24443 39933 24455 39936
rect 24397 39927 24455 39933
rect 25130 39924 25136 39936
rect 25188 39924 25194 39976
rect 19978 39828 19984 39840
rect 19939 39800 19984 39828
rect 19978 39788 19984 39800
rect 20036 39788 20042 39840
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 47673 39831 47731 39837
rect 47673 39828 47685 39831
rect 46532 39800 47685 39828
rect 46532 39788 46538 39800
rect 47673 39797 47685 39800
rect 47719 39797 47731 39831
rect 47673 39791 47731 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 22925 39627 22983 39633
rect 22925 39593 22937 39627
rect 22971 39624 22983 39627
rect 23474 39624 23480 39636
rect 22971 39596 23480 39624
rect 22971 39593 22983 39596
rect 22925 39587 22983 39593
rect 23474 39584 23480 39596
rect 23532 39584 23538 39636
rect 25130 39624 25136 39636
rect 25091 39596 25136 39624
rect 25130 39584 25136 39596
rect 25188 39584 25194 39636
rect 26050 39584 26056 39636
rect 26108 39624 26114 39636
rect 26602 39624 26608 39636
rect 26108 39596 26372 39624
rect 26563 39596 26608 39624
rect 26108 39584 26114 39596
rect 26234 39516 26240 39568
rect 26292 39516 26298 39568
rect 26252 39488 26280 39516
rect 26344 39497 26372 39596
rect 26602 39584 26608 39596
rect 26660 39584 26666 39636
rect 47026 39556 47032 39568
rect 46308 39528 47032 39556
rect 46308 39497 46336 39528
rect 47026 39516 47032 39528
rect 47084 39516 47090 39568
rect 25332 39460 26280 39488
rect 26329 39491 26387 39497
rect 18138 39380 18144 39432
rect 18196 39420 18202 39432
rect 19245 39423 19303 39429
rect 19245 39420 19257 39423
rect 18196 39392 19257 39420
rect 18196 39380 18202 39392
rect 19245 39389 19257 39392
rect 19291 39389 19303 39423
rect 19245 39383 19303 39389
rect 22094 39380 22100 39432
rect 22152 39420 22158 39432
rect 25332 39429 25360 39460
rect 26329 39457 26341 39491
rect 26375 39457 26387 39491
rect 26329 39451 26387 39457
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39457 46351 39491
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46293 39451 46351 39457
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 22833 39423 22891 39429
rect 22833 39420 22845 39423
rect 22152 39392 22845 39420
rect 22152 39380 22158 39392
rect 22833 39389 22845 39392
rect 22879 39389 22891 39423
rect 22833 39383 22891 39389
rect 25317 39423 25375 39429
rect 25317 39389 25329 39423
rect 25363 39389 25375 39423
rect 25317 39383 25375 39389
rect 26237 39423 26295 39429
rect 26237 39389 26249 39423
rect 26283 39420 26295 39423
rect 26418 39420 26424 39432
rect 26283 39392 26424 39420
rect 26283 39389 26295 39392
rect 26237 39383 26295 39389
rect 26418 39380 26424 39392
rect 26476 39380 26482 39432
rect 18966 39312 18972 39364
rect 19024 39352 19030 39364
rect 19521 39355 19579 39361
rect 19521 39352 19533 39355
rect 19024 39324 19533 39352
rect 19024 39312 19030 39324
rect 19521 39321 19533 39324
rect 19567 39321 19579 39355
rect 19521 39315 19579 39321
rect 19978 39312 19984 39364
rect 20036 39312 20042 39364
rect 20990 39284 20996 39296
rect 20951 39256 20996 39284
rect 20990 39244 20996 39256
rect 21048 39244 21054 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 18966 39080 18972 39092
rect 18927 39052 18972 39080
rect 18966 39040 18972 39052
rect 19024 39040 19030 39092
rect 19613 39083 19671 39089
rect 19613 39049 19625 39083
rect 19659 39049 19671 39083
rect 19613 39043 19671 39049
rect 19981 39083 20039 39089
rect 19981 39049 19993 39083
rect 20027 39080 20039 39083
rect 20990 39080 20996 39092
rect 20027 39052 20996 39080
rect 20027 39049 20039 39052
rect 19981 39043 20039 39049
rect 19153 38947 19211 38953
rect 19153 38913 19165 38947
rect 19199 38944 19211 38947
rect 19628 38944 19656 39043
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 25130 38972 25136 39024
rect 25188 38972 25194 39024
rect 26329 39015 26387 39021
rect 26329 38981 26341 39015
rect 26375 39012 26387 39015
rect 26375 38984 27738 39012
rect 26375 38981 26387 38984
rect 26329 38975 26387 38981
rect 19199 38916 19656 38944
rect 19199 38913 19211 38916
rect 19153 38907 19211 38913
rect 21818 38904 21824 38956
rect 21876 38944 21882 38956
rect 21913 38947 21971 38953
rect 21913 38944 21925 38947
rect 21876 38916 21925 38944
rect 21876 38904 21882 38916
rect 21913 38913 21925 38916
rect 21959 38913 21971 38947
rect 21913 38907 21971 38913
rect 23201 38947 23259 38953
rect 23201 38913 23213 38947
rect 23247 38944 23259 38947
rect 23474 38944 23480 38956
rect 23247 38916 23480 38944
rect 23247 38913 23259 38916
rect 23201 38907 23259 38913
rect 23474 38904 23480 38916
rect 23532 38904 23538 38956
rect 26237 38947 26295 38953
rect 26237 38913 26249 38947
rect 26283 38913 26295 38947
rect 29914 38944 29920 38956
rect 29875 38916 29920 38944
rect 26237 38907 26295 38913
rect 20070 38876 20076 38888
rect 20031 38848 20076 38876
rect 20070 38836 20076 38848
rect 20128 38836 20134 38888
rect 20162 38836 20168 38888
rect 20220 38876 20226 38888
rect 20220 38848 20265 38876
rect 20220 38836 20226 38848
rect 22002 38836 22008 38888
rect 22060 38876 22066 38888
rect 23842 38876 23848 38888
rect 22060 38848 23848 38876
rect 22060 38836 22066 38848
rect 23842 38836 23848 38848
rect 23900 38836 23906 38888
rect 24118 38876 24124 38888
rect 24079 38848 24124 38876
rect 24118 38836 24124 38848
rect 24176 38836 24182 38888
rect 24762 38836 24768 38888
rect 24820 38876 24826 38888
rect 26252 38876 26280 38907
rect 29914 38904 29920 38916
rect 29972 38904 29978 38956
rect 45554 38904 45560 38956
rect 45612 38944 45618 38956
rect 46109 38947 46167 38953
rect 46109 38944 46121 38947
rect 45612 38916 46121 38944
rect 45612 38904 45618 38916
rect 46109 38913 46121 38916
rect 46155 38913 46167 38947
rect 47854 38944 47860 38956
rect 47815 38916 47860 38944
rect 46109 38907 46167 38913
rect 47854 38904 47860 38916
rect 47912 38904 47918 38956
rect 24820 38848 26280 38876
rect 26973 38879 27031 38885
rect 24820 38836 24826 38848
rect 26973 38845 26985 38879
rect 27019 38876 27031 38879
rect 27246 38876 27252 38888
rect 27019 38848 27108 38876
rect 27207 38848 27252 38876
rect 27019 38845 27031 38848
rect 26973 38839 27031 38845
rect 19242 38700 19248 38752
rect 19300 38740 19306 38752
rect 22094 38740 22100 38752
rect 19300 38712 22100 38740
rect 19300 38700 19306 38712
rect 22094 38700 22100 38712
rect 22152 38740 22158 38752
rect 23290 38740 23296 38752
rect 22152 38712 22197 38740
rect 23251 38712 23296 38740
rect 22152 38700 22158 38712
rect 23290 38700 23296 38712
rect 23348 38700 23354 38752
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25593 38743 25651 38749
rect 25593 38740 25605 38743
rect 25372 38712 25605 38740
rect 25372 38700 25378 38712
rect 25593 38709 25605 38712
rect 25639 38709 25651 38743
rect 27080 38740 27108 38848
rect 27246 38836 27252 38848
rect 27304 38836 27310 38888
rect 27338 38836 27344 38888
rect 27396 38876 27402 38888
rect 28721 38879 28779 38885
rect 28721 38876 28733 38879
rect 27396 38848 28733 38876
rect 27396 38836 27402 38848
rect 28721 38845 28733 38848
rect 28767 38845 28779 38879
rect 30006 38876 30012 38888
rect 29967 38848 30012 38876
rect 28721 38839 28779 38845
rect 30006 38836 30012 38848
rect 30064 38836 30070 38888
rect 30098 38836 30104 38888
rect 30156 38876 30162 38888
rect 30156 38848 30201 38876
rect 30156 38836 30162 38848
rect 29822 38808 29828 38820
rect 28276 38780 29828 38808
rect 28276 38740 28304 38780
rect 29822 38768 29828 38780
rect 29880 38768 29886 38820
rect 27080 38712 28304 38740
rect 25593 38703 25651 38709
rect 28994 38700 29000 38752
rect 29052 38740 29058 38752
rect 29549 38743 29607 38749
rect 29549 38740 29561 38743
rect 29052 38712 29561 38740
rect 29052 38700 29058 38712
rect 29549 38709 29561 38712
rect 29595 38709 29607 38743
rect 29549 38703 29607 38709
rect 46201 38743 46259 38749
rect 46201 38709 46213 38743
rect 46247 38740 46259 38743
rect 46382 38740 46388 38752
rect 46247 38712 46388 38740
rect 46247 38709 46259 38712
rect 46201 38703 46259 38709
rect 46382 38700 46388 38712
rect 46440 38700 46446 38752
rect 46566 38700 46572 38752
rect 46624 38740 46630 38752
rect 48041 38743 48099 38749
rect 48041 38740 48053 38743
rect 46624 38712 48053 38740
rect 46624 38700 46630 38712
rect 48041 38709 48053 38712
rect 48087 38709 48099 38743
rect 48041 38703 48099 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 20070 38496 20076 38548
rect 20128 38536 20134 38548
rect 20165 38539 20223 38545
rect 20165 38536 20177 38539
rect 20128 38508 20177 38536
rect 20128 38496 20134 38508
rect 20165 38505 20177 38508
rect 20211 38505 20223 38539
rect 20165 38499 20223 38505
rect 24118 38496 24124 38548
rect 24176 38536 24182 38548
rect 24397 38539 24455 38545
rect 24397 38536 24409 38539
rect 24176 38508 24409 38536
rect 24176 38496 24182 38508
rect 24397 38505 24409 38508
rect 24443 38505 24455 38539
rect 25130 38536 25136 38548
rect 25091 38508 25136 38536
rect 24397 38499 24455 38505
rect 25130 38496 25136 38508
rect 25188 38496 25194 38548
rect 25314 38496 25320 38548
rect 25372 38536 25378 38548
rect 25961 38539 26019 38545
rect 25961 38536 25973 38539
rect 25372 38508 25973 38536
rect 25372 38496 25378 38508
rect 25961 38505 25973 38508
rect 26007 38505 26019 38539
rect 25961 38499 26019 38505
rect 29914 38496 29920 38548
rect 29972 38536 29978 38548
rect 31297 38539 31355 38545
rect 31297 38536 31309 38539
rect 29972 38508 31309 38536
rect 29972 38496 29978 38508
rect 31297 38505 31309 38508
rect 31343 38505 31355 38539
rect 31297 38499 31355 38505
rect 20438 38360 20444 38412
rect 20496 38400 20502 38412
rect 20717 38403 20775 38409
rect 20717 38400 20729 38403
rect 20496 38372 20729 38400
rect 20496 38360 20502 38372
rect 20717 38369 20729 38372
rect 20763 38369 20775 38403
rect 20717 38363 20775 38369
rect 23474 38360 23480 38412
rect 23532 38400 23538 38412
rect 24762 38400 24768 38412
rect 23532 38372 24768 38400
rect 23532 38360 23538 38372
rect 24762 38360 24768 38372
rect 24820 38400 24826 38412
rect 26145 38403 26203 38409
rect 24820 38372 25084 38400
rect 24820 38360 24826 38372
rect 18506 38292 18512 38344
rect 18564 38332 18570 38344
rect 19242 38332 19248 38344
rect 18564 38304 19248 38332
rect 18564 38292 18570 38304
rect 19242 38292 19248 38304
rect 19300 38292 19306 38344
rect 20530 38332 20536 38344
rect 20491 38304 20536 38332
rect 20530 38292 20536 38304
rect 20588 38292 20594 38344
rect 21174 38292 21180 38344
rect 21232 38332 21238 38344
rect 22002 38332 22008 38344
rect 21232 38304 22008 38332
rect 21232 38292 21238 38304
rect 22002 38292 22008 38304
rect 22060 38292 22066 38344
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38332 24639 38335
rect 24946 38332 24952 38344
rect 24627 38304 24952 38332
rect 24627 38301 24639 38304
rect 24581 38295 24639 38301
rect 24946 38292 24952 38304
rect 25004 38292 25010 38344
rect 25056 38341 25084 38372
rect 26145 38369 26157 38403
rect 26191 38400 26203 38403
rect 26510 38400 26516 38412
rect 26191 38372 26516 38400
rect 26191 38369 26203 38372
rect 26145 38363 26203 38369
rect 26510 38360 26516 38372
rect 26568 38400 26574 38412
rect 27522 38400 27528 38412
rect 26568 38372 27292 38400
rect 27483 38372 27528 38400
rect 26568 38360 26574 38372
rect 25041 38335 25099 38341
rect 25041 38301 25053 38335
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 26237 38335 26295 38341
rect 26237 38301 26249 38335
rect 26283 38332 26295 38335
rect 26418 38332 26424 38344
rect 26283 38304 26424 38332
rect 26283 38301 26295 38304
rect 26237 38295 26295 38301
rect 26418 38292 26424 38304
rect 26476 38292 26482 38344
rect 27264 38341 27292 38372
rect 27522 38360 27528 38372
rect 27580 38360 27586 38412
rect 29549 38403 29607 38409
rect 29549 38369 29561 38403
rect 29595 38400 29607 38403
rect 29822 38400 29828 38412
rect 29595 38372 29828 38400
rect 29595 38369 29607 38372
rect 29549 38363 29607 38369
rect 29822 38360 29828 38372
rect 29880 38360 29886 38412
rect 46382 38400 46388 38412
rect 46343 38372 46388 38400
rect 46382 38360 46388 38372
rect 46440 38360 46446 38412
rect 48038 38400 48044 38412
rect 47999 38372 48044 38400
rect 48038 38360 48044 38372
rect 48096 38360 48102 38412
rect 27249 38335 27307 38341
rect 27249 38301 27261 38335
rect 27295 38332 27307 38335
rect 27338 38332 27344 38344
rect 27295 38304 27344 38332
rect 27295 38301 27307 38304
rect 27249 38295 27307 38301
rect 27338 38292 27344 38304
rect 27396 38292 27402 38344
rect 28994 38332 29000 38344
rect 28955 38304 29000 38332
rect 28994 38292 29000 38304
rect 29052 38292 29058 38344
rect 46106 38292 46112 38344
rect 46164 38332 46170 38344
rect 46201 38335 46259 38341
rect 46201 38332 46213 38335
rect 46164 38304 46213 38332
rect 46164 38292 46170 38304
rect 46201 38301 46213 38304
rect 46247 38301 46259 38335
rect 46201 38295 46259 38301
rect 22281 38267 22339 38273
rect 22281 38233 22293 38267
rect 22327 38264 22339 38267
rect 22370 38264 22376 38276
rect 22327 38236 22376 38264
rect 22327 38233 22339 38236
rect 22281 38227 22339 38233
rect 22370 38224 22376 38236
rect 22428 38224 22434 38276
rect 23290 38224 23296 38276
rect 23348 38224 23354 38276
rect 25958 38264 25964 38276
rect 25919 38236 25964 38264
rect 25958 38224 25964 38236
rect 26016 38224 26022 38276
rect 29825 38267 29883 38273
rect 29825 38233 29837 38267
rect 29871 38233 29883 38267
rect 31110 38264 31116 38276
rect 31050 38236 31116 38264
rect 29825 38227 29883 38233
rect 19334 38196 19340 38208
rect 19295 38168 19340 38196
rect 19334 38156 19340 38168
rect 19392 38156 19398 38208
rect 20530 38156 20536 38208
rect 20588 38196 20594 38208
rect 20625 38199 20683 38205
rect 20625 38196 20637 38199
rect 20588 38168 20637 38196
rect 20588 38156 20594 38168
rect 20625 38165 20637 38168
rect 20671 38165 20683 38199
rect 23750 38196 23756 38208
rect 23711 38168 23756 38196
rect 20625 38159 20683 38165
rect 23750 38156 23756 38168
rect 23808 38156 23814 38208
rect 26418 38196 26424 38208
rect 26379 38168 26424 38196
rect 26418 38156 26424 38168
rect 26476 38156 26482 38208
rect 26881 38199 26939 38205
rect 26881 38165 26893 38199
rect 26927 38196 26939 38199
rect 27154 38196 27160 38208
rect 26927 38168 27160 38196
rect 26927 38165 26939 38168
rect 26881 38159 26939 38165
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 27338 38156 27344 38208
rect 27396 38196 27402 38208
rect 28813 38199 28871 38205
rect 27396 38168 27441 38196
rect 27396 38156 27402 38168
rect 28813 38165 28825 38199
rect 28859 38196 28871 38199
rect 29840 38196 29868 38227
rect 31110 38224 31116 38236
rect 31168 38224 31174 38276
rect 28859 38168 29868 38196
rect 28859 38165 28871 38168
rect 28813 38159 28871 38165
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 11698 37952 11704 38004
rect 11756 37992 11762 38004
rect 22186 37992 22192 38004
rect 11756 37964 22192 37992
rect 11756 37952 11762 37964
rect 22186 37952 22192 37964
rect 22244 37952 22250 38004
rect 22370 37992 22376 38004
rect 22331 37964 22376 37992
rect 22370 37952 22376 37964
rect 22428 37952 22434 38004
rect 24946 37992 24952 38004
rect 24907 37964 24952 37992
rect 24946 37952 24952 37964
rect 25004 37952 25010 38004
rect 26973 37995 27031 38001
rect 26973 37961 26985 37995
rect 27019 37992 27031 37995
rect 27246 37992 27252 38004
rect 27019 37964 27252 37992
rect 27019 37961 27031 37964
rect 26973 37955 27031 37961
rect 27246 37952 27252 37964
rect 27304 37952 27310 38004
rect 29825 37995 29883 38001
rect 29825 37961 29837 37995
rect 29871 37992 29883 37995
rect 30006 37992 30012 38004
rect 29871 37964 30012 37992
rect 29871 37961 29883 37964
rect 29825 37955 29883 37961
rect 30006 37952 30012 37964
rect 30064 37952 30070 38004
rect 31110 37992 31116 38004
rect 31071 37964 31116 37992
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 18138 37924 18144 37936
rect 17604 37896 18144 37924
rect 17494 37748 17500 37800
rect 17552 37788 17558 37800
rect 17604 37797 17632 37896
rect 18138 37884 18144 37896
rect 18196 37884 18202 37936
rect 19334 37924 19340 37936
rect 19090 37896 19340 37924
rect 19334 37884 19340 37896
rect 19392 37884 19398 37936
rect 21818 37884 21824 37936
rect 21876 37924 21882 37936
rect 21876 37896 23060 37924
rect 21876 37884 21882 37896
rect 20165 37859 20223 37865
rect 20165 37825 20177 37859
rect 20211 37856 20223 37859
rect 20990 37856 20996 37868
rect 20211 37828 20996 37856
rect 20211 37825 20223 37828
rect 20165 37819 20223 37825
rect 20990 37816 20996 37828
rect 21048 37816 21054 37868
rect 22554 37856 22560 37868
rect 22515 37828 22560 37856
rect 22554 37816 22560 37828
rect 22612 37816 22618 37868
rect 23032 37865 23060 37896
rect 25148 37896 25636 37924
rect 23017 37859 23075 37865
rect 23017 37825 23029 37859
rect 23063 37825 23075 37859
rect 23017 37819 23075 37825
rect 17589 37791 17647 37797
rect 17589 37788 17601 37791
rect 17552 37760 17601 37788
rect 17552 37748 17558 37760
rect 17589 37757 17601 37760
rect 17635 37757 17647 37791
rect 17589 37751 17647 37757
rect 17865 37791 17923 37797
rect 17865 37757 17877 37791
rect 17911 37788 17923 37791
rect 18230 37788 18236 37800
rect 17911 37760 18236 37788
rect 17911 37757 17923 37760
rect 17865 37751 17923 37757
rect 18230 37748 18236 37760
rect 18288 37748 18294 37800
rect 19426 37748 19432 37800
rect 19484 37788 19490 37800
rect 20073 37791 20131 37797
rect 20073 37788 20085 37791
rect 19484 37760 20085 37788
rect 19484 37748 19490 37760
rect 20073 37757 20085 37760
rect 20119 37757 20131 37791
rect 25148 37788 25176 37896
rect 25314 37856 25320 37868
rect 25275 37828 25320 37856
rect 25314 37816 25320 37828
rect 25372 37816 25378 37868
rect 25406 37788 25412 37800
rect 20073 37751 20131 37757
rect 20180 37760 25176 37788
rect 25367 37760 25412 37788
rect 20180 37732 20208 37760
rect 25406 37748 25412 37760
rect 25464 37748 25470 37800
rect 25608 37797 25636 37896
rect 25774 37884 25780 37936
rect 25832 37924 25838 37936
rect 25832 37896 35894 37924
rect 25832 37884 25838 37896
rect 27154 37856 27160 37868
rect 27115 37828 27160 37856
rect 27154 37816 27160 37828
rect 27212 37816 27218 37868
rect 30193 37859 30251 37865
rect 30193 37856 30205 37859
rect 29472 37828 30205 37856
rect 25593 37791 25651 37797
rect 25593 37757 25605 37791
rect 25639 37788 25651 37791
rect 27522 37788 27528 37800
rect 25639 37760 27528 37788
rect 25639 37757 25651 37760
rect 25593 37751 25651 37757
rect 27522 37748 27528 37760
rect 27580 37748 27586 37800
rect 20162 37680 20168 37732
rect 20220 37680 20226 37732
rect 20530 37720 20536 37732
rect 20491 37692 20536 37720
rect 20530 37680 20536 37692
rect 20588 37680 20594 37732
rect 22186 37680 22192 37732
rect 22244 37720 22250 37732
rect 29472 37729 29500 37828
rect 30193 37825 30205 37828
rect 30239 37825 30251 37859
rect 30193 37819 30251 37825
rect 30926 37816 30932 37868
rect 30984 37856 30990 37868
rect 31021 37859 31079 37865
rect 31021 37856 31033 37859
rect 30984 37828 31033 37856
rect 30984 37816 30990 37828
rect 31021 37825 31033 37828
rect 31067 37825 31079 37859
rect 31021 37819 31079 37825
rect 33137 37859 33195 37865
rect 33137 37825 33149 37859
rect 33183 37856 33195 37859
rect 33226 37856 33232 37868
rect 33183 37828 33232 37856
rect 33183 37825 33195 37828
rect 33137 37819 33195 37825
rect 33226 37816 33232 37828
rect 33284 37816 33290 37868
rect 35866 37856 35894 37896
rect 46290 37856 46296 37868
rect 35866 37828 46296 37856
rect 46290 37816 46296 37828
rect 46348 37856 46354 37868
rect 46661 37859 46719 37865
rect 46661 37856 46673 37859
rect 46348 37828 46673 37856
rect 46348 37816 46354 37828
rect 46661 37825 46673 37828
rect 46707 37825 46719 37859
rect 46661 37819 46719 37825
rect 30006 37748 30012 37800
rect 30064 37788 30070 37800
rect 30285 37791 30343 37797
rect 30285 37788 30297 37791
rect 30064 37760 30297 37788
rect 30064 37748 30070 37760
rect 30285 37757 30297 37760
rect 30331 37757 30343 37791
rect 30285 37751 30343 37757
rect 30469 37791 30527 37797
rect 30469 37757 30481 37791
rect 30515 37788 30527 37791
rect 34698 37788 34704 37800
rect 30515 37760 34704 37788
rect 30515 37757 30527 37760
rect 30469 37751 30527 37757
rect 34698 37748 34704 37760
rect 34756 37748 34762 37800
rect 29457 37723 29515 37729
rect 29457 37720 29469 37723
rect 22244 37692 29469 37720
rect 22244 37680 22250 37692
rect 29457 37689 29469 37692
rect 29503 37689 29515 37723
rect 29457 37683 29515 37689
rect 19334 37652 19340 37664
rect 19295 37624 19340 37652
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 23201 37655 23259 37661
rect 23201 37621 23213 37655
rect 23247 37652 23259 37655
rect 23474 37652 23480 37664
rect 23247 37624 23480 37652
rect 23247 37621 23259 37624
rect 23201 37615 23259 37621
rect 23474 37612 23480 37624
rect 23532 37612 23538 37664
rect 23658 37612 23664 37664
rect 23716 37652 23722 37664
rect 27890 37652 27896 37664
rect 23716 37624 27896 37652
rect 23716 37612 23722 37624
rect 27890 37612 27896 37624
rect 27948 37652 27954 37664
rect 30098 37652 30104 37664
rect 27948 37624 30104 37652
rect 27948 37612 27954 37624
rect 30098 37612 30104 37624
rect 30156 37612 30162 37664
rect 32674 37612 32680 37664
rect 32732 37652 32738 37664
rect 32953 37655 33011 37661
rect 32953 37652 32965 37655
rect 32732 37624 32965 37652
rect 32732 37612 32738 37624
rect 32953 37621 32965 37624
rect 32999 37621 33011 37655
rect 32953 37615 33011 37621
rect 46474 37612 46480 37664
rect 46532 37652 46538 37664
rect 46753 37655 46811 37661
rect 46753 37652 46765 37655
rect 46532 37624 46765 37652
rect 46532 37612 46538 37624
rect 46753 37621 46765 37624
rect 46799 37621 46811 37655
rect 47762 37652 47768 37664
rect 47723 37624 47768 37652
rect 46753 37615 46811 37621
rect 47762 37612 47768 37624
rect 47820 37612 47826 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 18230 37448 18236 37460
rect 18191 37420 18236 37448
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 22554 37408 22560 37460
rect 22612 37448 22618 37460
rect 23109 37451 23167 37457
rect 23109 37448 23121 37451
rect 22612 37420 23121 37448
rect 22612 37408 22618 37420
rect 23109 37417 23121 37420
rect 23155 37417 23167 37451
rect 27338 37448 27344 37460
rect 27299 37420 27344 37448
rect 23109 37411 23167 37417
rect 27338 37408 27344 37420
rect 27396 37408 27402 37460
rect 30006 37448 30012 37460
rect 29967 37420 30012 37448
rect 30006 37408 30012 37420
rect 30064 37408 30070 37460
rect 26881 37383 26939 37389
rect 26881 37349 26893 37383
rect 26927 37380 26939 37383
rect 26927 37352 27844 37380
rect 26927 37349 26939 37352
rect 26881 37343 26939 37349
rect 19889 37315 19947 37321
rect 19889 37281 19901 37315
rect 19935 37312 19947 37315
rect 20070 37312 20076 37324
rect 19935 37284 20076 37312
rect 19935 37281 19947 37284
rect 19889 37275 19947 37281
rect 20070 37272 20076 37284
rect 20128 37272 20134 37324
rect 23658 37312 23664 37324
rect 23619 37284 23664 37312
rect 23658 37272 23664 37284
rect 23716 37272 23722 37324
rect 26605 37315 26663 37321
rect 26605 37312 26617 37315
rect 26252 37284 26617 37312
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37244 18475 37247
rect 18463 37216 19288 37244
rect 18463 37213 18475 37216
rect 18417 37207 18475 37213
rect 19260 37117 19288 37216
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19392 37216 19625 37244
rect 19392 37204 19398 37216
rect 19613 37213 19625 37216
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 23477 37247 23535 37253
rect 23477 37213 23489 37247
rect 23523 37244 23535 37247
rect 23750 37244 23756 37256
rect 23523 37216 23756 37244
rect 23523 37213 23535 37216
rect 23477 37207 23535 37213
rect 23750 37204 23756 37216
rect 23808 37204 23814 37256
rect 24670 37244 24676 37256
rect 24631 37216 24676 37244
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 24857 37247 24915 37253
rect 24857 37213 24869 37247
rect 24903 37244 24915 37247
rect 25130 37244 25136 37256
rect 24903 37216 25136 37244
rect 24903 37213 24915 37216
rect 24857 37207 24915 37213
rect 25130 37204 25136 37216
rect 25188 37244 25194 37256
rect 26252 37244 26280 37284
rect 26605 37281 26617 37284
rect 26651 37312 26663 37315
rect 27338 37312 27344 37324
rect 26651 37284 27344 37312
rect 26651 37281 26663 37284
rect 26605 37275 26663 37281
rect 27338 37272 27344 37284
rect 27396 37272 27402 37324
rect 26510 37244 26516 37256
rect 25188 37216 26280 37244
rect 26471 37216 26516 37244
rect 25188 37204 25194 37216
rect 26510 37204 26516 37216
rect 26568 37204 26574 37256
rect 27816 37253 27844 37352
rect 27893 37315 27951 37321
rect 27893 37281 27905 37315
rect 27939 37281 27951 37315
rect 29638 37312 29644 37324
rect 29599 37284 29644 37312
rect 27893 37275 27951 37281
rect 27801 37247 27859 37253
rect 27801 37213 27813 37247
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 25590 37136 25596 37188
rect 25648 37176 25654 37188
rect 27908 37176 27936 37275
rect 29638 37272 29644 37284
rect 29696 37272 29702 37324
rect 29914 37312 29920 37324
rect 29748 37284 29920 37312
rect 29748 37253 29776 37284
rect 29914 37272 29920 37284
rect 29972 37272 29978 37324
rect 32674 37312 32680 37324
rect 32635 37284 32680 37312
rect 32674 37272 32680 37284
rect 32732 37272 32738 37324
rect 34698 37272 34704 37324
rect 34756 37312 34762 37324
rect 35250 37312 35256 37324
rect 34756 37284 35256 37312
rect 34756 37272 34762 37284
rect 35250 37272 35256 37284
rect 35308 37272 35314 37324
rect 46474 37312 46480 37324
rect 46435 37284 46480 37312
rect 46474 37272 46480 37284
rect 46532 37272 46538 37324
rect 48130 37312 48136 37324
rect 48091 37284 48136 37312
rect 48130 37272 48136 37284
rect 48188 37272 48194 37324
rect 29733 37247 29791 37253
rect 29733 37213 29745 37247
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 29822 37204 29828 37256
rect 29880 37244 29886 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 29880 37216 32413 37244
rect 29880 37204 29886 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 35069 37247 35127 37253
rect 35069 37213 35081 37247
rect 35115 37244 35127 37247
rect 35342 37244 35348 37256
rect 35115 37216 35348 37244
rect 35115 37213 35127 37216
rect 35069 37207 35127 37213
rect 35342 37204 35348 37216
rect 35400 37204 35406 37256
rect 46293 37247 46351 37253
rect 46293 37213 46305 37247
rect 46339 37213 46351 37247
rect 46293 37207 46351 37213
rect 25648 37148 27936 37176
rect 25648 37136 25654 37148
rect 33686 37136 33692 37188
rect 33744 37136 33750 37188
rect 46308 37176 46336 37207
rect 47762 37176 47768 37188
rect 46308 37148 47768 37176
rect 47762 37136 47768 37148
rect 47820 37136 47826 37188
rect 19245 37111 19303 37117
rect 19245 37077 19257 37111
rect 19291 37077 19303 37111
rect 19245 37071 19303 37077
rect 19705 37111 19763 37117
rect 19705 37077 19717 37111
rect 19751 37108 19763 37111
rect 19978 37108 19984 37120
rect 19751 37080 19984 37108
rect 19751 37077 19763 37080
rect 19705 37071 19763 37077
rect 19978 37068 19984 37080
rect 20036 37068 20042 37120
rect 23566 37068 23572 37120
rect 23624 37108 23630 37120
rect 24762 37108 24768 37120
rect 23624 37080 23669 37108
rect 24723 37080 24768 37108
rect 23624 37068 23630 37080
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 27709 37111 27767 37117
rect 27709 37077 27721 37111
rect 27755 37108 27767 37111
rect 28166 37108 28172 37120
rect 27755 37080 28172 37108
rect 27755 37077 27767 37080
rect 27709 37071 27767 37077
rect 28166 37068 28172 37080
rect 28224 37068 28230 37120
rect 33962 37068 33968 37120
rect 34020 37108 34026 37120
rect 34149 37111 34207 37117
rect 34149 37108 34161 37111
rect 34020 37080 34161 37108
rect 34020 37068 34026 37080
rect 34149 37077 34161 37080
rect 34195 37077 34207 37111
rect 34698 37108 34704 37120
rect 34659 37080 34704 37108
rect 34149 37071 34207 37077
rect 34698 37068 34704 37080
rect 34756 37068 34762 37120
rect 35158 37068 35164 37120
rect 35216 37108 35222 37120
rect 35216 37080 35261 37108
rect 35216 37068 35222 37080
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 19889 36907 19947 36913
rect 19889 36873 19901 36907
rect 19935 36904 19947 36907
rect 19978 36904 19984 36916
rect 19935 36876 19984 36904
rect 19935 36873 19947 36876
rect 19889 36867 19947 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 23477 36907 23535 36913
rect 23477 36873 23489 36907
rect 23523 36904 23535 36907
rect 23566 36904 23572 36916
rect 23523 36876 23572 36904
rect 23523 36873 23535 36876
rect 23477 36867 23535 36873
rect 23566 36864 23572 36876
rect 23624 36864 23630 36916
rect 23937 36907 23995 36913
rect 23937 36873 23949 36907
rect 23983 36904 23995 36907
rect 24762 36904 24768 36916
rect 23983 36876 24768 36904
rect 23983 36873 23995 36876
rect 23937 36867 23995 36873
rect 24762 36864 24768 36876
rect 24820 36864 24826 36916
rect 26510 36904 26516 36916
rect 25884 36876 26516 36904
rect 23750 36796 23756 36848
rect 23808 36836 23814 36848
rect 24854 36836 24860 36848
rect 23808 36808 24860 36836
rect 23808 36796 23814 36808
rect 24854 36796 24860 36808
rect 24912 36836 24918 36848
rect 24949 36839 25007 36845
rect 24949 36836 24961 36839
rect 24912 36808 24961 36836
rect 24912 36796 24918 36808
rect 24949 36805 24961 36808
rect 24995 36805 25007 36839
rect 25130 36836 25136 36848
rect 25091 36808 25136 36836
rect 24949 36799 25007 36805
rect 25130 36796 25136 36808
rect 25188 36796 25194 36848
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 19242 36768 19248 36780
rect 19203 36740 19248 36768
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 20254 36768 20260 36780
rect 20215 36740 20260 36768
rect 20254 36728 20260 36740
rect 20312 36728 20318 36780
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 23845 36771 23903 36777
rect 22152 36740 22197 36768
rect 22152 36728 22158 36740
rect 23845 36737 23857 36771
rect 23891 36768 23903 36771
rect 23934 36768 23940 36780
rect 23891 36740 23940 36768
rect 23891 36737 23903 36740
rect 23845 36731 23903 36737
rect 23934 36728 23940 36740
rect 23992 36728 23998 36780
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36768 24823 36771
rect 25038 36768 25044 36780
rect 24811 36740 25044 36768
rect 24811 36737 24823 36740
rect 24765 36731 24823 36737
rect 25038 36728 25044 36740
rect 25096 36728 25102 36780
rect 25314 36728 25320 36780
rect 25372 36768 25378 36780
rect 25884 36777 25912 36876
rect 26510 36864 26516 36876
rect 26568 36864 26574 36916
rect 30098 36864 30104 36916
rect 30156 36904 30162 36916
rect 33137 36907 33195 36913
rect 30156 36876 31754 36904
rect 30156 36864 30162 36876
rect 30374 36836 30380 36848
rect 29196 36808 30380 36836
rect 25685 36771 25743 36777
rect 25685 36768 25697 36771
rect 25372 36740 25697 36768
rect 25372 36728 25378 36740
rect 25685 36737 25697 36740
rect 25731 36737 25743 36771
rect 25685 36731 25743 36737
rect 25869 36771 25927 36777
rect 25869 36737 25881 36771
rect 25915 36737 25927 36771
rect 25869 36731 25927 36737
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 19337 36703 19395 36709
rect 19337 36669 19349 36703
rect 19383 36700 19395 36703
rect 20349 36703 20407 36709
rect 20349 36700 20361 36703
rect 19383 36672 20361 36700
rect 19383 36669 19395 36672
rect 19337 36663 19395 36669
rect 20349 36669 20361 36672
rect 20395 36669 20407 36703
rect 20349 36663 20407 36669
rect 20438 36660 20444 36712
rect 20496 36700 20502 36712
rect 20533 36703 20591 36709
rect 20533 36700 20545 36703
rect 20496 36672 20545 36700
rect 20496 36660 20502 36672
rect 20533 36669 20545 36672
rect 20579 36700 20591 36703
rect 24029 36703 24087 36709
rect 24029 36700 24041 36703
rect 20579 36672 24041 36700
rect 20579 36669 20591 36672
rect 20533 36663 20591 36669
rect 24029 36669 24041 36672
rect 24075 36700 24087 36703
rect 25590 36700 25596 36712
rect 24075 36672 25596 36700
rect 24075 36669 24087 36672
rect 24029 36663 24087 36669
rect 25590 36660 25596 36672
rect 25648 36660 25654 36712
rect 25700 36700 25728 36731
rect 25958 36728 25964 36780
rect 26016 36768 26022 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 26016 36740 26065 36768
rect 26016 36728 26022 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26234 36768 26240 36780
rect 26195 36740 26240 36768
rect 26053 36731 26111 36737
rect 26234 36728 26240 36740
rect 26292 36728 26298 36780
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 26344 36740 27169 36768
rect 26344 36700 26372 36740
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27338 36768 27344 36780
rect 27299 36740 27344 36768
rect 27157 36731 27215 36737
rect 27338 36728 27344 36740
rect 27396 36728 27402 36780
rect 29196 36777 29224 36808
rect 30374 36796 30380 36808
rect 30432 36796 30438 36848
rect 31110 36796 31116 36848
rect 31168 36796 31174 36848
rect 29181 36771 29239 36777
rect 29181 36737 29193 36771
rect 29227 36737 29239 36771
rect 29181 36731 29239 36737
rect 29365 36771 29423 36777
rect 29365 36737 29377 36771
rect 29411 36768 29423 36771
rect 29638 36768 29644 36780
rect 29411 36740 29644 36768
rect 29411 36737 29423 36740
rect 29365 36731 29423 36737
rect 29638 36728 29644 36740
rect 29696 36728 29702 36780
rect 25700 36672 26372 36700
rect 26421 36703 26479 36709
rect 26421 36669 26433 36703
rect 26467 36700 26479 36703
rect 26510 36700 26516 36712
rect 26467 36672 26516 36700
rect 26467 36669 26479 36672
rect 26421 36663 26479 36669
rect 26510 36660 26516 36672
rect 26568 36660 26574 36712
rect 26602 36660 26608 36712
rect 26660 36700 26666 36712
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 26660 36672 27445 36700
rect 26660 36660 26666 36672
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 29822 36700 29828 36712
rect 29783 36672 29828 36700
rect 27433 36663 27491 36669
rect 29822 36660 29828 36672
rect 29880 36660 29886 36712
rect 30098 36700 30104 36712
rect 30059 36672 30104 36700
rect 30098 36660 30104 36672
rect 30156 36660 30162 36712
rect 30190 36660 30196 36712
rect 30248 36700 30254 36712
rect 31573 36703 31631 36709
rect 31573 36700 31585 36703
rect 30248 36672 31585 36700
rect 30248 36660 30254 36672
rect 31573 36669 31585 36672
rect 31619 36669 31631 36703
rect 31726 36700 31754 36876
rect 33137 36873 33149 36907
rect 33183 36904 33195 36907
rect 33226 36904 33232 36916
rect 33183 36876 33232 36904
rect 33183 36873 33195 36876
rect 33137 36867 33195 36873
rect 33226 36864 33232 36876
rect 33284 36864 33290 36916
rect 33597 36907 33655 36913
rect 33597 36873 33609 36907
rect 33643 36904 33655 36907
rect 34698 36904 34704 36916
rect 33643 36876 34704 36904
rect 33643 36873 33655 36876
rect 33597 36867 33655 36873
rect 34698 36864 34704 36876
rect 34756 36864 34762 36916
rect 34885 36907 34943 36913
rect 34885 36873 34897 36907
rect 34931 36904 34943 36907
rect 35158 36904 35164 36916
rect 34931 36876 35164 36904
rect 34931 36873 34943 36876
rect 34885 36867 34943 36873
rect 35158 36864 35164 36876
rect 35216 36864 35222 36916
rect 33505 36771 33563 36777
rect 33505 36737 33517 36771
rect 33551 36768 33563 36771
rect 33962 36768 33968 36780
rect 33551 36740 33968 36768
rect 33551 36737 33563 36740
rect 33505 36731 33563 36737
rect 33962 36728 33968 36740
rect 34020 36768 34026 36780
rect 34517 36771 34575 36777
rect 34517 36768 34529 36771
rect 34020 36740 34529 36768
rect 34020 36728 34026 36740
rect 34517 36737 34529 36740
rect 34563 36737 34575 36771
rect 34517 36731 34575 36737
rect 33689 36703 33747 36709
rect 33689 36700 33701 36703
rect 31726 36672 33701 36700
rect 31573 36663 31631 36669
rect 33689 36669 33701 36672
rect 33735 36669 33747 36703
rect 34606 36700 34612 36712
rect 34567 36672 34612 36700
rect 33689 36663 33747 36669
rect 34606 36660 34612 36672
rect 34664 36660 34670 36712
rect 12434 36592 12440 36644
rect 12492 36632 12498 36644
rect 26786 36632 26792 36644
rect 12492 36604 26792 36632
rect 12492 36592 12498 36604
rect 26786 36592 26792 36604
rect 26844 36592 26850 36644
rect 22186 36564 22192 36576
rect 22147 36536 22192 36564
rect 22186 36524 22192 36536
rect 22244 36524 22250 36576
rect 24854 36524 24860 36576
rect 24912 36564 24918 36576
rect 25958 36564 25964 36576
rect 24912 36536 25964 36564
rect 24912 36524 24918 36536
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 26142 36524 26148 36576
rect 26200 36564 26206 36576
rect 26973 36567 27031 36573
rect 26973 36564 26985 36567
rect 26200 36536 26985 36564
rect 26200 36524 26206 36536
rect 26973 36533 26985 36536
rect 27019 36533 27031 36567
rect 26973 36527 27031 36533
rect 29181 36567 29239 36573
rect 29181 36533 29193 36567
rect 29227 36564 29239 36567
rect 30834 36564 30840 36576
rect 29227 36536 30840 36564
rect 29227 36533 29239 36536
rect 29181 36527 29239 36533
rect 30834 36524 30840 36536
rect 30892 36524 30898 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 6886 36332 24624 36360
rect 2038 36252 2044 36304
rect 2096 36292 2102 36304
rect 6886 36292 6914 36332
rect 2096 36264 6914 36292
rect 2096 36252 2102 36264
rect 19242 36252 19248 36304
rect 19300 36292 19306 36304
rect 19429 36295 19487 36301
rect 19429 36292 19441 36295
rect 19300 36264 19441 36292
rect 19300 36252 19306 36264
rect 19429 36261 19441 36264
rect 19475 36261 19487 36295
rect 19429 36255 19487 36261
rect 19610 36252 19616 36304
rect 19668 36292 19674 36304
rect 19978 36292 19984 36304
rect 19668 36264 19984 36292
rect 19668 36252 19674 36264
rect 19978 36252 19984 36264
rect 20036 36292 20042 36304
rect 20625 36295 20683 36301
rect 20625 36292 20637 36295
rect 20036 36264 20637 36292
rect 20036 36252 20042 36264
rect 20625 36261 20637 36264
rect 20671 36261 20683 36295
rect 20625 36255 20683 36261
rect 19518 36224 19524 36236
rect 19479 36196 19524 36224
rect 19518 36184 19524 36196
rect 19576 36184 19582 36236
rect 20717 36227 20775 36233
rect 20717 36193 20729 36227
rect 20763 36224 20775 36227
rect 20990 36224 20996 36236
rect 20763 36196 20996 36224
rect 20763 36193 20775 36196
rect 20717 36187 20775 36193
rect 20990 36184 20996 36196
rect 21048 36184 21054 36236
rect 21453 36227 21511 36233
rect 21453 36193 21465 36227
rect 21499 36224 21511 36227
rect 22462 36224 22468 36236
rect 21499 36196 22468 36224
rect 21499 36193 21511 36196
rect 21453 36187 21511 36193
rect 22462 36184 22468 36196
rect 22520 36184 22526 36236
rect 24596 36224 24624 36332
rect 24670 36320 24676 36372
rect 24728 36360 24734 36372
rect 24765 36363 24823 36369
rect 24765 36360 24777 36363
rect 24728 36332 24777 36360
rect 24728 36320 24734 36332
rect 24765 36329 24777 36332
rect 24811 36329 24823 36363
rect 24765 36323 24823 36329
rect 25406 36320 25412 36372
rect 25464 36360 25470 36372
rect 25777 36363 25835 36369
rect 25777 36360 25789 36363
rect 25464 36332 25789 36360
rect 25464 36320 25470 36332
rect 25777 36329 25789 36332
rect 25823 36329 25835 36363
rect 26234 36360 26240 36372
rect 25777 36323 25835 36329
rect 25976 36332 26240 36360
rect 25038 36252 25044 36304
rect 25096 36292 25102 36304
rect 25976 36292 26004 36332
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 28905 36363 28963 36369
rect 28905 36329 28917 36363
rect 28951 36360 28963 36363
rect 29086 36360 29092 36372
rect 28951 36332 29092 36360
rect 28951 36329 28963 36332
rect 28905 36323 28963 36329
rect 29086 36320 29092 36332
rect 29144 36360 29150 36372
rect 29638 36360 29644 36372
rect 29144 36332 29644 36360
rect 29144 36320 29150 36332
rect 29638 36320 29644 36332
rect 29696 36320 29702 36372
rect 30098 36320 30104 36372
rect 30156 36360 30162 36372
rect 30285 36363 30343 36369
rect 30285 36360 30297 36363
rect 30156 36332 30297 36360
rect 30156 36320 30162 36332
rect 30285 36329 30297 36332
rect 30331 36329 30343 36363
rect 30285 36323 30343 36329
rect 31021 36363 31079 36369
rect 31021 36329 31033 36363
rect 31067 36360 31079 36363
rect 31110 36360 31116 36372
rect 31067 36332 31116 36360
rect 31067 36329 31079 36332
rect 31021 36323 31079 36329
rect 31110 36320 31116 36332
rect 31168 36320 31174 36372
rect 33597 36363 33655 36369
rect 33597 36329 33609 36363
rect 33643 36360 33655 36363
rect 33686 36360 33692 36372
rect 33643 36332 33692 36360
rect 33643 36329 33655 36332
rect 33597 36323 33655 36329
rect 33686 36320 33692 36332
rect 33744 36320 33750 36372
rect 26142 36292 26148 36304
rect 25096 36264 26004 36292
rect 26103 36264 26148 36292
rect 25096 36252 25102 36264
rect 26142 36252 26148 36264
rect 26200 36252 26206 36304
rect 28736 36264 30052 36292
rect 24596 36196 28212 36224
rect 2130 36156 2136 36168
rect 2091 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36116 2194 36168
rect 18506 36156 18512 36168
rect 18467 36128 18512 36156
rect 18506 36116 18512 36128
rect 18564 36116 18570 36168
rect 19242 36156 19248 36168
rect 19203 36128 19248 36156
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 20441 36159 20499 36165
rect 19392 36128 19437 36156
rect 19392 36116 19398 36128
rect 20441 36125 20453 36159
rect 20487 36125 20499 36159
rect 21174 36156 21180 36168
rect 21135 36128 21180 36156
rect 20441 36119 20499 36125
rect 20346 36048 20352 36100
rect 20404 36088 20410 36100
rect 20456 36088 20484 36119
rect 21174 36116 21180 36128
rect 21232 36116 21238 36168
rect 24673 36159 24731 36165
rect 24673 36125 24685 36159
rect 24719 36125 24731 36159
rect 24854 36156 24860 36168
rect 24815 36128 24860 36156
rect 24673 36119 24731 36125
rect 20404 36060 21220 36088
rect 20404 36048 20410 36060
rect 18506 35980 18512 36032
rect 18564 36020 18570 36032
rect 18601 36023 18659 36029
rect 18601 36020 18613 36023
rect 18564 35992 18613 36020
rect 18564 35980 18570 35992
rect 18601 35989 18613 35992
rect 18647 35989 18659 36023
rect 18601 35983 18659 35989
rect 20257 36023 20315 36029
rect 20257 35989 20269 36023
rect 20303 36020 20315 36023
rect 21082 36020 21088 36032
rect 20303 35992 21088 36020
rect 20303 35989 20315 35992
rect 20257 35983 20315 35989
rect 21082 35980 21088 35992
rect 21140 35980 21146 36032
rect 21192 36020 21220 36060
rect 22186 36048 22192 36100
rect 22244 36048 22250 36100
rect 24688 36088 24716 36119
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 25961 36159 26019 36165
rect 25961 36125 25973 36159
rect 26007 36125 26019 36159
rect 25961 36119 26019 36125
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36125 26111 36159
rect 26053 36119 26111 36125
rect 26237 36159 26295 36165
rect 26237 36125 26249 36159
rect 26283 36156 26295 36159
rect 27157 36159 27215 36165
rect 27157 36156 27169 36159
rect 26283 36128 27169 36156
rect 26283 36125 26295 36128
rect 26237 36119 26295 36125
rect 27157 36125 27169 36128
rect 27203 36125 27215 36159
rect 27157 36119 27215 36125
rect 25038 36088 25044 36100
rect 24688 36060 25044 36088
rect 25038 36048 25044 36060
rect 25096 36048 25102 36100
rect 22370 36020 22376 36032
rect 21192 35992 22376 36020
rect 22370 35980 22376 35992
rect 22428 36020 22434 36032
rect 22925 36023 22983 36029
rect 22925 36020 22937 36023
rect 22428 35992 22937 36020
rect 22428 35980 22434 35992
rect 22925 35989 22937 35992
rect 22971 35989 22983 36023
rect 25976 36020 26004 36119
rect 26068 36088 26096 36119
rect 26510 36088 26516 36100
rect 26068 36060 26516 36088
rect 26510 36048 26516 36060
rect 26568 36048 26574 36100
rect 26786 36088 26792 36100
rect 26747 36060 26792 36088
rect 26786 36048 26792 36060
rect 26844 36048 26850 36100
rect 26973 36091 27031 36097
rect 26973 36057 26985 36091
rect 27019 36088 27031 36091
rect 28074 36088 28080 36100
rect 27019 36060 28080 36088
rect 27019 36057 27031 36060
rect 26973 36051 27031 36057
rect 28074 36048 28080 36060
rect 28132 36048 28138 36100
rect 28184 36088 28212 36196
rect 28736 36165 28764 36264
rect 29917 36227 29975 36233
rect 29917 36224 29929 36227
rect 28828 36196 29929 36224
rect 28721 36159 28779 36165
rect 28721 36125 28733 36159
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 28828 36088 28856 36196
rect 29917 36193 29929 36196
rect 29963 36193 29975 36227
rect 29917 36187 29975 36193
rect 30024 36224 30052 36264
rect 30190 36224 30196 36236
rect 30024 36196 30196 36224
rect 28994 36156 29000 36168
rect 28955 36128 29000 36156
rect 28994 36116 29000 36128
rect 29052 36116 29058 36168
rect 29549 36159 29607 36165
rect 29549 36125 29561 36159
rect 29595 36125 29607 36159
rect 29730 36156 29736 36168
rect 29691 36128 29736 36156
rect 29549 36119 29607 36125
rect 28184 36060 28856 36088
rect 29564 36088 29592 36119
rect 29730 36116 29736 36128
rect 29788 36116 29794 36168
rect 29825 36159 29883 36165
rect 29825 36125 29837 36159
rect 29871 36156 29883 36159
rect 30024 36156 30052 36196
rect 30190 36184 30196 36196
rect 30248 36184 30254 36236
rect 29871 36128 30052 36156
rect 30101 36159 30159 36165
rect 29871 36125 29883 36128
rect 29825 36119 29883 36125
rect 30101 36125 30113 36159
rect 30147 36156 30159 36159
rect 30466 36156 30472 36168
rect 30147 36128 30472 36156
rect 30147 36125 30159 36128
rect 30101 36119 30159 36125
rect 30466 36116 30472 36128
rect 30524 36116 30530 36168
rect 30926 36156 30932 36168
rect 30887 36128 30932 36156
rect 30926 36116 30932 36128
rect 30984 36116 30990 36168
rect 32306 36116 32312 36168
rect 32364 36156 32370 36168
rect 33505 36159 33563 36165
rect 33505 36156 33517 36159
rect 32364 36128 33517 36156
rect 32364 36116 32370 36128
rect 33505 36125 33517 36128
rect 33551 36125 33563 36159
rect 33505 36119 33563 36125
rect 31294 36088 31300 36100
rect 29564 36060 31300 36088
rect 31294 36048 31300 36060
rect 31352 36048 31358 36100
rect 27062 36020 27068 36032
rect 25976 35992 27068 36020
rect 22925 35983 22983 35989
rect 27062 35980 27068 35992
rect 27120 35980 27126 36032
rect 28537 36023 28595 36029
rect 28537 35989 28549 36023
rect 28583 36020 28595 36023
rect 30190 36020 30196 36032
rect 28583 35992 30196 36020
rect 28583 35989 28595 35992
rect 28537 35983 28595 35989
rect 30190 35980 30196 35992
rect 30248 35980 30254 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 17494 35776 17500 35828
rect 17552 35816 17558 35828
rect 21174 35816 21180 35828
rect 17552 35788 21180 35816
rect 17552 35776 17558 35788
rect 21174 35776 21180 35788
rect 21232 35776 21238 35828
rect 21358 35776 21364 35828
rect 21416 35816 21422 35828
rect 21416 35788 22048 35816
rect 21416 35776 21422 35788
rect 17773 35751 17831 35757
rect 17773 35717 17785 35751
rect 17819 35748 17831 35751
rect 17819 35720 19380 35748
rect 17819 35717 17831 35720
rect 17773 35711 17831 35717
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 17954 35680 17960 35692
rect 17915 35652 17960 35680
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18616 35689 18644 35720
rect 19352 35692 19380 35720
rect 21082 35708 21088 35760
rect 21140 35748 21146 35760
rect 21140 35720 21956 35748
rect 21140 35708 21146 35720
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35649 18659 35683
rect 18601 35643 18659 35649
rect 18785 35683 18843 35689
rect 18785 35649 18797 35683
rect 18831 35649 18843 35683
rect 19334 35680 19340 35692
rect 19247 35652 19340 35680
rect 18785 35643 18843 35649
rect 17972 35612 18000 35640
rect 18800 35612 18828 35643
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 19426 35640 19432 35692
rect 19484 35680 19490 35692
rect 20165 35683 20223 35689
rect 20165 35680 20177 35683
rect 19484 35652 20177 35680
rect 19484 35640 19490 35652
rect 20165 35649 20177 35652
rect 20211 35649 20223 35683
rect 20346 35680 20352 35692
rect 20307 35652 20352 35680
rect 20165 35643 20223 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21744 35652 21833 35680
rect 17972 35584 18828 35612
rect 19352 35612 19380 35640
rect 20438 35612 20444 35624
rect 19352 35584 20444 35612
rect 16666 35504 16672 35556
rect 16724 35544 16730 35556
rect 18693 35547 18751 35553
rect 18693 35544 18705 35547
rect 16724 35516 18705 35544
rect 16724 35504 16730 35516
rect 18693 35513 18705 35516
rect 18739 35513 18751 35547
rect 18693 35507 18751 35513
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 1854 35476 1860 35488
rect 1443 35448 1860 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 1854 35436 1860 35448
rect 1912 35436 1918 35488
rect 16942 35436 16948 35488
rect 17000 35476 17006 35488
rect 18141 35479 18199 35485
rect 18141 35476 18153 35479
rect 17000 35448 18153 35476
rect 17000 35436 17006 35448
rect 18141 35445 18153 35448
rect 18187 35445 18199 35479
rect 18800 35476 18828 35584
rect 20438 35572 20444 35584
rect 20496 35572 20502 35624
rect 19705 35547 19763 35553
rect 19705 35513 19717 35547
rect 19751 35544 19763 35547
rect 19978 35544 19984 35556
rect 19751 35516 19984 35544
rect 19751 35513 19763 35516
rect 19705 35507 19763 35513
rect 19978 35504 19984 35516
rect 20036 35504 20042 35556
rect 20990 35544 20996 35556
rect 20364 35516 20996 35544
rect 19242 35476 19248 35488
rect 18800 35448 19248 35476
rect 18141 35439 18199 35445
rect 19242 35436 19248 35448
rect 19300 35476 19306 35488
rect 20364 35485 20392 35516
rect 20990 35504 20996 35516
rect 21048 35504 21054 35556
rect 21744 35544 21772 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 21928 35612 21956 35720
rect 22020 35689 22048 35788
rect 22462 35776 22468 35828
rect 22520 35816 22526 35828
rect 22557 35819 22615 35825
rect 22557 35816 22569 35819
rect 22520 35788 22569 35816
rect 22520 35776 22526 35788
rect 22557 35785 22569 35788
rect 22603 35785 22615 35819
rect 22557 35779 22615 35785
rect 30374 35776 30380 35828
rect 30432 35816 30438 35828
rect 30469 35819 30527 35825
rect 30469 35816 30481 35819
rect 30432 35788 30481 35816
rect 30432 35776 30438 35788
rect 30469 35785 30481 35788
rect 30515 35785 30527 35819
rect 31294 35816 31300 35828
rect 31255 35788 31300 35816
rect 30469 35779 30527 35785
rect 31294 35776 31300 35788
rect 31352 35776 31358 35828
rect 28994 35708 29000 35760
rect 29052 35748 29058 35760
rect 29914 35748 29920 35760
rect 29052 35720 29920 35748
rect 29052 35708 29058 35720
rect 29914 35708 29920 35720
rect 29972 35748 29978 35760
rect 30101 35751 30159 35757
rect 30101 35748 30113 35751
rect 29972 35720 30113 35748
rect 29972 35708 29978 35720
rect 30101 35717 30113 35720
rect 30147 35717 30159 35751
rect 30101 35711 30159 35717
rect 30190 35708 30196 35760
rect 30248 35748 30254 35760
rect 30248 35720 30972 35748
rect 30248 35708 30254 35720
rect 22005 35683 22063 35689
rect 22005 35649 22017 35683
rect 22051 35649 22063 35683
rect 22370 35680 22376 35692
rect 22331 35652 22376 35680
rect 22005 35643 22063 35649
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 30282 35680 30288 35692
rect 30243 35652 30288 35680
rect 30282 35640 30288 35652
rect 30340 35640 30346 35692
rect 30944 35689 30972 35720
rect 30929 35683 30987 35689
rect 30929 35649 30941 35683
rect 30975 35649 30987 35683
rect 48130 35680 48136 35692
rect 48091 35652 48136 35680
rect 30929 35643 30987 35649
rect 48130 35640 48136 35652
rect 48188 35640 48194 35692
rect 22097 35615 22155 35621
rect 22097 35612 22109 35615
rect 21928 35584 22109 35612
rect 22097 35581 22109 35584
rect 22143 35581 22155 35615
rect 22097 35575 22155 35581
rect 22186 35572 22192 35624
rect 22244 35612 22250 35624
rect 22244 35584 22289 35612
rect 22244 35572 22250 35584
rect 28074 35572 28080 35624
rect 28132 35612 28138 35624
rect 28813 35615 28871 35621
rect 28813 35612 28825 35615
rect 28132 35584 28825 35612
rect 28132 35572 28138 35584
rect 28813 35581 28825 35584
rect 28859 35581 28871 35615
rect 28813 35575 28871 35581
rect 29089 35615 29147 35621
rect 29089 35581 29101 35615
rect 29135 35612 29147 35615
rect 29178 35612 29184 35624
rect 29135 35584 29184 35612
rect 29135 35581 29147 35584
rect 29089 35575 29147 35581
rect 29178 35572 29184 35584
rect 29236 35612 29242 35624
rect 30466 35612 30472 35624
rect 29236 35584 30472 35612
rect 29236 35572 29242 35584
rect 30466 35572 30472 35584
rect 30524 35572 30530 35624
rect 31021 35615 31079 35621
rect 31021 35581 31033 35615
rect 31067 35581 31079 35615
rect 31021 35575 31079 35581
rect 28994 35544 29000 35556
rect 21744 35516 29000 35544
rect 28994 35504 29000 35516
rect 29052 35504 29058 35556
rect 29914 35504 29920 35556
rect 29972 35544 29978 35556
rect 31036 35544 31064 35575
rect 29972 35516 31064 35544
rect 29972 35504 29978 35516
rect 19337 35479 19395 35485
rect 19337 35476 19349 35479
rect 19300 35448 19349 35476
rect 19300 35436 19306 35448
rect 19337 35445 19349 35448
rect 19383 35445 19395 35479
rect 19337 35439 19395 35445
rect 20349 35479 20407 35485
rect 20349 35445 20361 35479
rect 20395 35445 20407 35479
rect 20530 35476 20536 35488
rect 20491 35448 20536 35476
rect 20349 35439 20407 35445
rect 20530 35436 20536 35448
rect 20588 35436 20594 35488
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 30929 35479 30987 35485
rect 30929 35476 30941 35479
rect 30892 35448 30941 35476
rect 30892 35436 30898 35448
rect 30929 35445 30941 35448
rect 30975 35445 30987 35479
rect 30929 35439 30987 35445
rect 47118 35436 47124 35488
rect 47176 35476 47182 35488
rect 47949 35479 48007 35485
rect 47949 35476 47961 35479
rect 47176 35448 47961 35476
rect 47176 35436 47182 35448
rect 47949 35445 47961 35448
rect 47995 35445 48007 35479
rect 47949 35439 48007 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 20438 35232 20444 35284
rect 20496 35272 20502 35284
rect 20625 35275 20683 35281
rect 20625 35272 20637 35275
rect 20496 35244 20637 35272
rect 20496 35232 20502 35244
rect 20625 35241 20637 35244
rect 20671 35241 20683 35275
rect 20625 35235 20683 35241
rect 21174 35232 21180 35284
rect 21232 35272 21238 35284
rect 22002 35272 22008 35284
rect 21232 35244 22008 35272
rect 21232 35232 21238 35244
rect 22002 35232 22008 35244
rect 22060 35272 22066 35284
rect 22557 35275 22615 35281
rect 22557 35272 22569 35275
rect 22060 35244 22569 35272
rect 22060 35232 22066 35244
rect 22557 35241 22569 35244
rect 22603 35241 22615 35275
rect 28994 35272 29000 35284
rect 28955 35244 29000 35272
rect 22557 35235 22615 35241
rect 28994 35232 29000 35244
rect 29052 35232 29058 35284
rect 33873 35275 33931 35281
rect 33873 35241 33885 35275
rect 33919 35272 33931 35275
rect 34606 35272 34612 35284
rect 33919 35244 34612 35272
rect 33919 35241 33931 35244
rect 33873 35235 33931 35241
rect 34606 35232 34612 35244
rect 34664 35232 34670 35284
rect 17954 35204 17960 35216
rect 17696 35176 17960 35204
rect 17696 35145 17724 35176
rect 17954 35164 17960 35176
rect 18012 35164 18018 35216
rect 17681 35139 17739 35145
rect 16776 35108 17540 35136
rect 16666 35068 16672 35080
rect 16627 35040 16672 35068
rect 16666 35028 16672 35040
rect 16724 35028 16730 35080
rect 16776 35000 16804 35108
rect 16942 35068 16948 35080
rect 16903 35040 16948 35068
rect 16942 35028 16948 35040
rect 17000 35028 17006 35080
rect 17405 35071 17463 35077
rect 17405 35037 17417 35071
rect 17451 35037 17463 35071
rect 17405 35031 17463 35037
rect 16853 35003 16911 35009
rect 16853 35000 16865 35003
rect 16776 34972 16865 35000
rect 16853 34969 16865 34972
rect 16899 34969 16911 35003
rect 17420 35000 17448 35031
rect 16853 34963 16911 34969
rect 16960 34972 17448 35000
rect 17512 35000 17540 35108
rect 17681 35105 17693 35139
rect 17727 35105 17739 35139
rect 19334 35136 19340 35148
rect 19247 35108 19340 35136
rect 17681 35099 17739 35105
rect 19334 35096 19340 35108
rect 19392 35136 19398 35148
rect 20346 35136 20352 35148
rect 19392 35108 20352 35136
rect 19392 35096 19398 35108
rect 20346 35096 20352 35108
rect 20404 35136 20410 35148
rect 20717 35139 20775 35145
rect 20717 35136 20729 35139
rect 20404 35108 20729 35136
rect 20404 35096 20410 35108
rect 20717 35105 20729 35108
rect 20763 35105 20775 35139
rect 20717 35099 20775 35105
rect 22186 35096 22192 35148
rect 22244 35136 22250 35148
rect 28169 35139 28227 35145
rect 28169 35136 28181 35139
rect 22244 35108 28181 35136
rect 22244 35096 22250 35108
rect 28169 35105 28181 35108
rect 28215 35136 28227 35139
rect 28215 35108 28764 35136
rect 28215 35105 28227 35108
rect 28169 35099 28227 35105
rect 17586 35028 17592 35080
rect 17644 35068 17650 35080
rect 17644 35040 17689 35068
rect 17644 35028 17650 35040
rect 17770 35028 17776 35080
rect 17828 35068 17834 35080
rect 17957 35071 18015 35077
rect 17828 35040 17873 35068
rect 17828 35028 17834 35040
rect 17957 35037 17969 35071
rect 18003 35068 18015 35071
rect 18230 35068 18236 35080
rect 18003 35040 18236 35068
rect 18003 35037 18015 35040
rect 17957 35031 18015 35037
rect 18230 35028 18236 35040
rect 18288 35028 18294 35080
rect 19242 35028 19248 35080
rect 19300 35068 19306 35080
rect 19613 35071 19671 35077
rect 19613 35068 19625 35071
rect 19300 35040 19625 35068
rect 19300 35028 19306 35040
rect 19613 35037 19625 35040
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 20530 35028 20536 35080
rect 20588 35068 20594 35080
rect 20625 35071 20683 35077
rect 20625 35068 20637 35071
rect 20588 35040 20637 35068
rect 20588 35028 20594 35040
rect 20625 35037 20637 35040
rect 20671 35037 20683 35071
rect 20625 35031 20683 35037
rect 23474 35028 23480 35080
rect 23532 35068 23538 35080
rect 23569 35071 23627 35077
rect 23569 35068 23581 35071
rect 23532 35040 23581 35068
rect 23532 35028 23538 35040
rect 23569 35037 23581 35040
rect 23615 35068 23627 35071
rect 24118 35068 24124 35080
rect 23615 35040 24124 35068
rect 23615 35037 23627 35040
rect 23569 35031 23627 35037
rect 24118 35028 24124 35040
rect 24176 35028 24182 35080
rect 19150 35000 19156 35012
rect 17512 34972 19156 35000
rect 16960 34941 16988 34972
rect 19150 34960 19156 34972
rect 19208 34960 19214 35012
rect 22465 35003 22523 35009
rect 22465 34969 22477 35003
rect 22511 35000 22523 35003
rect 22922 35000 22928 35012
rect 22511 34972 22928 35000
rect 22511 34969 22523 34972
rect 22465 34963 22523 34969
rect 22922 34960 22928 34972
rect 22980 34960 22986 35012
rect 27982 35000 27988 35012
rect 27943 34972 27988 35000
rect 27982 34960 27988 34972
rect 28040 34960 28046 35012
rect 28626 35000 28632 35012
rect 28587 34972 28632 35000
rect 28626 34960 28632 34972
rect 28684 34960 28690 35012
rect 28736 35000 28764 35108
rect 29270 35096 29276 35148
rect 29328 35136 29334 35148
rect 29822 35136 29828 35148
rect 29328 35108 29828 35136
rect 29328 35096 29334 35108
rect 29822 35096 29828 35108
rect 29880 35136 29886 35148
rect 31297 35139 31355 35145
rect 31297 35136 31309 35139
rect 29880 35108 31309 35136
rect 29880 35096 29886 35108
rect 31297 35105 31309 35108
rect 31343 35105 31355 35139
rect 33962 35136 33968 35148
rect 33923 35108 33968 35136
rect 31297 35099 31355 35105
rect 33962 35096 33968 35108
rect 34020 35096 34026 35148
rect 35342 35136 35348 35148
rect 35255 35108 35348 35136
rect 35342 35096 35348 35108
rect 35400 35136 35406 35148
rect 35802 35136 35808 35148
rect 35400 35108 35808 35136
rect 35400 35096 35406 35108
rect 35802 35096 35808 35108
rect 35860 35096 35866 35148
rect 28813 35071 28871 35077
rect 28813 35037 28825 35071
rect 28859 35068 28871 35071
rect 29178 35068 29184 35080
rect 28859 35040 29184 35068
rect 28859 35037 28871 35040
rect 28813 35031 28871 35037
rect 29178 35028 29184 35040
rect 29236 35028 29242 35080
rect 30006 35068 30012 35080
rect 29967 35040 30012 35068
rect 30006 35028 30012 35040
rect 30064 35028 30070 35080
rect 30193 35071 30251 35077
rect 30193 35037 30205 35071
rect 30239 35037 30251 35071
rect 30193 35031 30251 35037
rect 30285 35071 30343 35077
rect 30285 35037 30297 35071
rect 30331 35037 30343 35071
rect 30285 35031 30343 35037
rect 30377 35071 30435 35077
rect 30377 35037 30389 35071
rect 30423 35037 30435 35071
rect 30377 35031 30435 35037
rect 29730 35000 29736 35012
rect 28736 34972 29736 35000
rect 29730 34960 29736 34972
rect 29788 35000 29794 35012
rect 30098 35000 30104 35012
rect 29788 34972 30104 35000
rect 29788 34960 29794 34972
rect 30098 34960 30104 34972
rect 30156 35000 30162 35012
rect 30208 35000 30236 35031
rect 30156 34972 30236 35000
rect 30156 34960 30162 34972
rect 16945 34935 17003 34941
rect 16945 34901 16957 34935
rect 16991 34901 17003 34935
rect 16945 34895 17003 34901
rect 18046 34892 18052 34944
rect 18104 34932 18110 34944
rect 18141 34935 18199 34941
rect 18141 34932 18153 34935
rect 18104 34904 18153 34932
rect 18104 34892 18110 34904
rect 18141 34901 18153 34904
rect 18187 34901 18199 34935
rect 18141 34895 18199 34901
rect 20993 34935 21051 34941
rect 20993 34901 21005 34935
rect 21039 34932 21051 34935
rect 21450 34932 21456 34944
rect 21039 34904 21456 34932
rect 21039 34901 21051 34904
rect 20993 34895 21051 34901
rect 21450 34892 21456 34904
rect 21508 34892 21514 34944
rect 23566 34892 23572 34944
rect 23624 34932 23630 34944
rect 23661 34935 23719 34941
rect 23661 34932 23673 34935
rect 23624 34904 23673 34932
rect 23624 34892 23630 34904
rect 23661 34901 23673 34904
rect 23707 34901 23719 34935
rect 30300 34932 30328 35031
rect 30392 35000 30420 35031
rect 30466 35028 30472 35080
rect 30524 35068 30530 35080
rect 30561 35071 30619 35077
rect 30561 35068 30573 35071
rect 30524 35040 30573 35068
rect 30524 35028 30530 35040
rect 30561 35037 30573 35040
rect 30607 35037 30619 35071
rect 31202 35068 31208 35080
rect 30561 35031 30619 35037
rect 30668 35040 31208 35068
rect 30668 35000 30696 35040
rect 31202 35028 31208 35040
rect 31260 35028 31266 35080
rect 33689 35071 33747 35077
rect 33689 35068 33701 35071
rect 33060 35040 33701 35068
rect 30392 34972 30696 35000
rect 30745 35003 30803 35009
rect 30745 34969 30757 35003
rect 30791 35000 30803 35003
rect 31573 35003 31631 35009
rect 31573 35000 31585 35003
rect 30791 34972 31585 35000
rect 30791 34969 30803 34972
rect 30745 34963 30803 34969
rect 31573 34969 31585 34972
rect 31619 34969 31631 35003
rect 31573 34963 31631 34969
rect 32582 34960 32588 35012
rect 32640 34960 32646 35012
rect 33060 34941 33088 35040
rect 33689 35037 33701 35040
rect 33735 35037 33747 35071
rect 33689 35031 33747 35037
rect 33704 35000 33732 35031
rect 34790 35028 34796 35080
rect 34848 35068 34854 35080
rect 35069 35071 35127 35077
rect 35069 35068 35081 35071
rect 34848 35040 35081 35068
rect 34848 35028 34854 35040
rect 35069 35037 35081 35040
rect 35115 35037 35127 35071
rect 35069 35031 35127 35037
rect 47026 35028 47032 35080
rect 47084 35068 47090 35080
rect 47854 35068 47860 35080
rect 47084 35040 47860 35068
rect 47084 35028 47090 35040
rect 47854 35028 47860 35040
rect 47912 35028 47918 35080
rect 48038 35028 48044 35080
rect 48096 35068 48102 35080
rect 48133 35071 48191 35077
rect 48133 35068 48145 35071
rect 48096 35040 48145 35068
rect 48096 35028 48102 35040
rect 48133 35037 48145 35040
rect 48179 35037 48191 35071
rect 48133 35031 48191 35037
rect 34054 35000 34060 35012
rect 33704 34972 34060 35000
rect 34054 34960 34060 34972
rect 34112 34960 34118 35012
rect 33045 34935 33103 34941
rect 33045 34932 33057 34935
rect 30300 34904 33057 34932
rect 23661 34895 23719 34901
rect 33045 34901 33057 34904
rect 33091 34901 33103 34935
rect 33502 34932 33508 34944
rect 33463 34904 33508 34932
rect 33045 34895 33103 34901
rect 33502 34892 33508 34904
rect 33560 34892 33566 34944
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 34701 34935 34759 34941
rect 34701 34932 34713 34935
rect 34572 34904 34713 34932
rect 34572 34892 34578 34904
rect 34701 34901 34713 34904
rect 34747 34901 34759 34935
rect 34701 34895 34759 34901
rect 35161 34935 35219 34941
rect 35161 34901 35173 34935
rect 35207 34932 35219 34935
rect 35618 34932 35624 34944
rect 35207 34904 35624 34932
rect 35207 34901 35219 34904
rect 35161 34895 35219 34901
rect 35618 34892 35624 34904
rect 35676 34892 35682 34944
rect 47854 34892 47860 34944
rect 47912 34932 47918 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47912 34904 47961 34932
rect 47912 34892 47918 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 17586 34688 17592 34740
rect 17644 34728 17650 34740
rect 19245 34731 19303 34737
rect 17644 34700 19196 34728
rect 17644 34688 17650 34700
rect 17773 34663 17831 34669
rect 17773 34629 17785 34663
rect 17819 34660 17831 34663
rect 18046 34660 18052 34672
rect 17819 34632 18052 34660
rect 17819 34629 17831 34632
rect 17773 34623 17831 34629
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 18506 34620 18512 34672
rect 18564 34620 18570 34672
rect 19168 34660 19196 34700
rect 19245 34697 19257 34731
rect 19291 34728 19303 34731
rect 19334 34728 19340 34740
rect 19291 34700 19340 34728
rect 19291 34697 19303 34700
rect 19245 34691 19303 34697
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 25498 34688 25504 34740
rect 25556 34728 25562 34740
rect 28445 34731 28503 34737
rect 28445 34728 28457 34731
rect 25556 34700 28457 34728
rect 25556 34688 25562 34700
rect 28445 34697 28457 34700
rect 28491 34697 28503 34731
rect 28445 34691 28503 34697
rect 30006 34688 30012 34740
rect 30064 34728 30070 34740
rect 30285 34731 30343 34737
rect 30285 34728 30297 34731
rect 30064 34700 30297 34728
rect 30064 34688 30070 34700
rect 30285 34697 30297 34700
rect 30331 34697 30343 34731
rect 30285 34691 30343 34697
rect 31389 34731 31447 34737
rect 31389 34697 31401 34731
rect 31435 34697 31447 34731
rect 32582 34728 32588 34740
rect 32543 34700 32588 34728
rect 31389 34691 31447 34697
rect 21913 34663 21971 34669
rect 19168 34632 20300 34660
rect 17494 34592 17500 34604
rect 17455 34564 17500 34592
rect 17494 34552 17500 34564
rect 17552 34552 17558 34604
rect 20162 34524 20168 34536
rect 20123 34496 20168 34524
rect 20162 34484 20168 34496
rect 20220 34484 20226 34536
rect 20272 34524 20300 34632
rect 21913 34629 21925 34663
rect 21959 34660 21971 34663
rect 22186 34660 22192 34672
rect 21959 34632 22192 34660
rect 21959 34629 21971 34632
rect 21913 34623 21971 34629
rect 22186 34620 22192 34632
rect 22244 34620 22250 34672
rect 23566 34620 23572 34672
rect 23624 34620 23630 34672
rect 24118 34620 24124 34672
rect 24176 34660 24182 34672
rect 24176 34632 26188 34660
rect 24176 34620 24182 34632
rect 20438 34592 20444 34604
rect 20399 34564 20444 34592
rect 20438 34552 20444 34564
rect 20496 34552 20502 34604
rect 22002 34552 22008 34604
rect 22060 34592 22066 34604
rect 22557 34595 22615 34601
rect 22557 34592 22569 34595
rect 22060 34564 22569 34592
rect 22060 34552 22066 34564
rect 22557 34561 22569 34564
rect 22603 34561 22615 34595
rect 24762 34592 24768 34604
rect 24723 34564 24768 34592
rect 22557 34555 22615 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25038 34592 25044 34604
rect 24951 34564 25044 34592
rect 25038 34552 25044 34564
rect 25096 34592 25102 34604
rect 26160 34601 26188 34632
rect 26418 34620 26424 34672
rect 26476 34660 26482 34672
rect 26973 34663 27031 34669
rect 26973 34660 26985 34663
rect 26476 34632 26985 34660
rect 26476 34620 26482 34632
rect 26973 34629 26985 34632
rect 27019 34629 27031 34663
rect 29178 34660 29184 34672
rect 26973 34623 27031 34629
rect 28276 34632 29184 34660
rect 26145 34595 26203 34601
rect 25096 34564 25728 34592
rect 25096 34552 25102 34564
rect 22830 34524 22836 34536
rect 20272 34496 22140 34524
rect 22791 34496 22836 34524
rect 22112 34465 22140 34496
rect 22830 34484 22836 34496
rect 22888 34484 22894 34536
rect 25133 34527 25191 34533
rect 25133 34524 25145 34527
rect 24136 34496 25145 34524
rect 22097 34459 22155 34465
rect 22097 34425 22109 34459
rect 22143 34456 22155 34459
rect 22554 34456 22560 34468
rect 22143 34428 22560 34456
rect 22143 34425 22155 34428
rect 22097 34419 22155 34425
rect 22554 34416 22560 34428
rect 22612 34416 22618 34468
rect 19150 34348 19156 34400
rect 19208 34388 19214 34400
rect 21266 34388 21272 34400
rect 19208 34360 21272 34388
rect 19208 34348 19214 34360
rect 21266 34348 21272 34360
rect 21324 34388 21330 34400
rect 24136 34388 24164 34496
rect 25133 34493 25145 34496
rect 25179 34524 25191 34527
rect 25222 34524 25228 34536
rect 25179 34496 25228 34524
rect 25179 34493 25191 34496
rect 25133 34487 25191 34493
rect 25222 34484 25228 34496
rect 25280 34484 25286 34536
rect 25700 34524 25728 34564
rect 26145 34561 26157 34595
rect 26191 34561 26203 34595
rect 26145 34555 26203 34561
rect 27157 34595 27215 34601
rect 27157 34561 27169 34595
rect 27203 34592 27215 34595
rect 27246 34592 27252 34604
rect 27203 34564 27252 34592
rect 27203 34561 27215 34564
rect 27157 34555 27215 34561
rect 27246 34552 27252 34564
rect 27304 34552 27310 34604
rect 28276 34601 28304 34632
rect 29178 34620 29184 34632
rect 29236 34620 29242 34672
rect 31404 34660 31432 34691
rect 32582 34688 32588 34700
rect 32640 34688 32646 34740
rect 34241 34731 34299 34737
rect 34241 34728 34253 34731
rect 32692 34700 34253 34728
rect 32692 34660 32720 34700
rect 34241 34697 34253 34700
rect 34287 34697 34299 34731
rect 34241 34691 34299 34697
rect 34606 34688 34612 34740
rect 34664 34728 34670 34740
rect 35069 34731 35127 34737
rect 35069 34728 35081 34731
rect 34664 34700 35081 34728
rect 34664 34688 34670 34700
rect 35069 34697 35081 34700
rect 35115 34697 35127 34731
rect 35618 34728 35624 34740
rect 35579 34700 35624 34728
rect 35069 34691 35127 34697
rect 29748 34632 31432 34660
rect 31726 34632 32720 34660
rect 33781 34663 33839 34669
rect 29748 34604 29776 34632
rect 28261 34595 28319 34601
rect 28261 34561 28273 34595
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 28350 34552 28356 34604
rect 28408 34592 28414 34604
rect 29089 34595 29147 34601
rect 29089 34592 29101 34595
rect 28408 34564 29101 34592
rect 28408 34552 28414 34564
rect 29089 34561 29101 34564
rect 29135 34561 29147 34595
rect 29730 34592 29736 34604
rect 29643 34564 29736 34592
rect 29089 34555 29147 34561
rect 29730 34552 29736 34564
rect 29788 34552 29794 34604
rect 30929 34595 30987 34601
rect 30929 34561 30941 34595
rect 30975 34592 30987 34595
rect 31110 34592 31116 34604
rect 30975 34564 31116 34592
rect 30975 34561 30987 34564
rect 30929 34555 30987 34561
rect 31110 34552 31116 34564
rect 31168 34552 31174 34604
rect 31570 34592 31576 34604
rect 31531 34564 31576 34592
rect 31570 34552 31576 34564
rect 31628 34592 31634 34604
rect 31726 34592 31754 34632
rect 33781 34629 33793 34663
rect 33827 34660 33839 34663
rect 35084 34660 35112 34691
rect 35618 34688 35624 34700
rect 35676 34688 35682 34740
rect 33827 34632 34652 34660
rect 35084 34632 35756 34660
rect 33827 34629 33839 34632
rect 33781 34623 33839 34629
rect 34624 34604 34652 34632
rect 32490 34592 32496 34604
rect 31628 34564 31754 34592
rect 32451 34564 32496 34592
rect 31628 34552 31634 34564
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 34054 34592 34060 34604
rect 34015 34564 34060 34592
rect 34054 34552 34060 34564
rect 34112 34552 34118 34604
rect 34606 34552 34612 34604
rect 34664 34592 34670 34604
rect 34701 34595 34759 34601
rect 34701 34592 34713 34595
rect 34664 34564 34713 34592
rect 34664 34552 34670 34564
rect 34701 34561 34713 34564
rect 34747 34561 34759 34595
rect 34701 34555 34759 34561
rect 34790 34552 34796 34604
rect 34848 34592 34854 34604
rect 34885 34595 34943 34601
rect 34885 34592 34897 34595
rect 34848 34564 34897 34592
rect 34848 34552 34854 34564
rect 34885 34561 34897 34564
rect 34931 34561 34943 34595
rect 35526 34592 35532 34604
rect 35487 34564 35532 34592
rect 34885 34555 34943 34561
rect 35526 34552 35532 34564
rect 35584 34552 35590 34604
rect 35728 34601 35756 34632
rect 35713 34595 35771 34601
rect 35713 34561 35725 34595
rect 35759 34561 35771 34595
rect 47762 34592 47768 34604
rect 47723 34564 47768 34592
rect 35713 34555 35771 34561
rect 47762 34552 47768 34564
rect 47820 34552 47826 34604
rect 26237 34527 26295 34533
rect 25700 34496 26188 34524
rect 24210 34416 24216 34468
rect 24268 34456 24274 34468
rect 24857 34459 24915 34465
rect 24857 34456 24869 34459
rect 24268 34428 24869 34456
rect 24268 34416 24274 34428
rect 24857 34425 24869 34428
rect 24903 34425 24915 34459
rect 26160 34456 26188 34496
rect 26237 34493 26249 34527
rect 26283 34524 26295 34527
rect 26418 34524 26424 34536
rect 26283 34496 26424 34524
rect 26283 34493 26295 34496
rect 26237 34487 26295 34493
rect 26418 34484 26424 34496
rect 26476 34484 26482 34536
rect 29270 34524 29276 34536
rect 29231 34496 29276 34524
rect 29270 34484 29276 34496
rect 29328 34484 29334 34536
rect 29914 34484 29920 34536
rect 29972 34524 29978 34536
rect 30009 34527 30067 34533
rect 30009 34524 30021 34527
rect 29972 34496 30021 34524
rect 29972 34484 29978 34496
rect 30009 34493 30021 34496
rect 30055 34493 30067 34527
rect 30009 34487 30067 34493
rect 33965 34527 34023 34533
rect 33965 34493 33977 34527
rect 34011 34524 34023 34527
rect 34808 34524 34836 34552
rect 34011 34496 34836 34524
rect 34011 34493 34023 34496
rect 33965 34487 34023 34493
rect 27430 34456 27436 34468
rect 26160 34428 27436 34456
rect 24857 34419 24915 34425
rect 27430 34416 27436 34428
rect 27488 34416 27494 34468
rect 33502 34456 33508 34468
rect 30116 34428 33508 34456
rect 24302 34388 24308 34400
rect 21324 34360 24164 34388
rect 24263 34360 24308 34388
rect 21324 34348 21330 34360
rect 24302 34348 24308 34360
rect 24360 34348 24366 34400
rect 24946 34348 24952 34400
rect 25004 34388 25010 34400
rect 27338 34388 27344 34400
rect 25004 34360 25049 34388
rect 27299 34360 27344 34388
rect 25004 34348 25010 34360
rect 27338 34348 27344 34360
rect 27396 34348 27402 34400
rect 30116 34397 30144 34428
rect 33502 34416 33508 34428
rect 33560 34416 33566 34468
rect 30101 34391 30159 34397
rect 30101 34357 30113 34391
rect 30147 34357 30159 34391
rect 30742 34388 30748 34400
rect 30703 34360 30748 34388
rect 30101 34351 30159 34357
rect 30742 34348 30748 34360
rect 30800 34348 30806 34400
rect 33962 34388 33968 34400
rect 33923 34360 33968 34388
rect 33962 34348 33968 34360
rect 34020 34348 34026 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47581 34391 47639 34397
rect 47581 34388 47593 34391
rect 47268 34360 47593 34388
rect 47268 34348 47274 34360
rect 47581 34357 47593 34360
rect 47627 34357 47639 34391
rect 47581 34351 47639 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 20162 34144 20168 34196
rect 20220 34184 20226 34196
rect 20533 34187 20591 34193
rect 20533 34184 20545 34187
rect 20220 34156 20545 34184
rect 20220 34144 20226 34156
rect 20533 34153 20545 34156
rect 20579 34184 20591 34187
rect 20806 34184 20812 34196
rect 20579 34156 20812 34184
rect 20579 34153 20591 34156
rect 20533 34147 20591 34153
rect 20806 34144 20812 34156
rect 20864 34144 20870 34196
rect 21358 34184 21364 34196
rect 21319 34156 21364 34184
rect 21358 34144 21364 34156
rect 21416 34144 21422 34196
rect 22830 34144 22836 34196
rect 22888 34184 22894 34196
rect 23477 34187 23535 34193
rect 23477 34184 23489 34187
rect 22888 34156 23489 34184
rect 22888 34144 22894 34156
rect 23477 34153 23489 34156
rect 23523 34153 23535 34187
rect 23477 34147 23535 34153
rect 24581 34187 24639 34193
rect 24581 34153 24593 34187
rect 24627 34184 24639 34187
rect 24762 34184 24768 34196
rect 24627 34156 24768 34184
rect 24627 34153 24639 34156
rect 24581 34147 24639 34153
rect 24762 34144 24768 34156
rect 24820 34144 24826 34196
rect 27154 34144 27160 34196
rect 27212 34184 27218 34196
rect 27341 34187 27399 34193
rect 27341 34184 27353 34187
rect 27212 34156 27353 34184
rect 27212 34144 27218 34156
rect 27341 34153 27353 34156
rect 27387 34153 27399 34187
rect 27341 34147 27399 34153
rect 27430 34144 27436 34196
rect 27488 34184 27494 34196
rect 27801 34187 27859 34193
rect 27801 34184 27813 34187
rect 27488 34156 27813 34184
rect 27488 34144 27494 34156
rect 27801 34153 27813 34156
rect 27847 34153 27859 34187
rect 27801 34147 27859 34153
rect 34793 34187 34851 34193
rect 34793 34153 34805 34187
rect 34839 34184 34851 34187
rect 35526 34184 35532 34196
rect 34839 34156 35532 34184
rect 34839 34153 34851 34156
rect 34793 34147 34851 34153
rect 35526 34144 35532 34156
rect 35584 34144 35590 34196
rect 9490 34076 9496 34128
rect 9548 34116 9554 34128
rect 29270 34116 29276 34128
rect 9548 34088 22094 34116
rect 9548 34076 9554 34088
rect 20438 34048 20444 34060
rect 20399 34020 20444 34048
rect 20438 34008 20444 34020
rect 20496 34008 20502 34060
rect 22066 34048 22094 34088
rect 27356 34088 29276 34116
rect 23109 34051 23167 34057
rect 23109 34048 23121 34051
rect 22066 34020 23121 34048
rect 23109 34017 23121 34020
rect 23155 34017 23167 34051
rect 23109 34011 23167 34017
rect 25133 34051 25191 34057
rect 25133 34017 25145 34051
rect 25179 34048 25191 34051
rect 27356 34048 27384 34088
rect 29270 34076 29276 34088
rect 29328 34076 29334 34128
rect 25179 34020 27384 34048
rect 27525 34051 27583 34057
rect 25179 34017 25191 34020
rect 25133 34011 25191 34017
rect 27525 34017 27537 34051
rect 27571 34048 27583 34051
rect 27706 34048 27712 34060
rect 27571 34020 27712 34048
rect 27571 34017 27583 34020
rect 27525 34011 27583 34017
rect 27706 34008 27712 34020
rect 27764 34008 27770 34060
rect 28629 34051 28687 34057
rect 28629 34017 28641 34051
rect 28675 34048 28687 34051
rect 28902 34048 28908 34060
rect 28675 34020 28908 34048
rect 28675 34017 28687 34020
rect 28629 34011 28687 34017
rect 28902 34008 28908 34020
rect 28960 34048 28966 34060
rect 30193 34051 30251 34057
rect 30193 34048 30205 34051
rect 28960 34020 30205 34048
rect 28960 34008 28966 34020
rect 30193 34017 30205 34020
rect 30239 34048 30251 34051
rect 30742 34048 30748 34060
rect 30239 34020 30748 34048
rect 30239 34017 30251 34020
rect 30193 34011 30251 34017
rect 30742 34008 30748 34020
rect 30800 34008 30806 34060
rect 32858 34008 32864 34060
rect 32916 34048 32922 34060
rect 33965 34051 34023 34057
rect 33965 34048 33977 34051
rect 32916 34020 33977 34048
rect 32916 34008 32922 34020
rect 33965 34017 33977 34020
rect 34011 34017 34023 34051
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 33965 34011 34023 34017
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47578 34048 47584 34060
rect 47539 34020 47584 34048
rect 47578 34008 47584 34020
rect 47636 34008 47642 34060
rect 1578 33980 1584 33992
rect 1539 33952 1584 33980
rect 1578 33940 1584 33952
rect 1636 33940 1642 33992
rect 20346 33940 20352 33992
rect 20404 33980 20410 33992
rect 20533 33983 20591 33989
rect 20533 33980 20545 33983
rect 20404 33952 20545 33980
rect 20404 33940 20410 33952
rect 20533 33949 20545 33952
rect 20579 33949 20591 33983
rect 21266 33980 21272 33992
rect 21227 33952 21272 33980
rect 20533 33943 20591 33949
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 21450 33980 21456 33992
rect 21411 33952 21456 33980
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 22738 33980 22744 33992
rect 22699 33952 22744 33980
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 22830 33940 22836 33992
rect 22888 33980 22894 33992
rect 22925 33983 22983 33989
rect 22925 33980 22937 33983
rect 22888 33952 22937 33980
rect 22888 33940 22894 33952
rect 22925 33949 22937 33952
rect 22971 33949 22983 33983
rect 22925 33943 22983 33949
rect 23017 33983 23075 33989
rect 23017 33949 23029 33983
rect 23063 33949 23075 33983
rect 23290 33980 23296 33992
rect 23251 33952 23296 33980
rect 23017 33943 23075 33949
rect 20257 33915 20315 33921
rect 20257 33881 20269 33915
rect 20303 33912 20315 33915
rect 20898 33912 20904 33924
rect 20303 33884 20904 33912
rect 20303 33881 20315 33884
rect 20257 33875 20315 33881
rect 20898 33872 20904 33884
rect 20956 33872 20962 33924
rect 23032 33912 23060 33943
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 24489 33983 24547 33989
rect 24489 33949 24501 33983
rect 24535 33949 24547 33983
rect 24489 33943 24547 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33949 27675 33983
rect 27617 33943 27675 33949
rect 28813 33983 28871 33989
rect 28813 33949 28825 33983
rect 28859 33980 28871 33983
rect 29178 33980 29184 33992
rect 28859 33952 29184 33980
rect 28859 33949 28871 33952
rect 28813 33943 28871 33949
rect 23750 33912 23756 33924
rect 23032 33884 23756 33912
rect 23750 33872 23756 33884
rect 23808 33912 23814 33924
rect 24302 33912 24308 33924
rect 23808 33884 24308 33912
rect 23808 33872 23814 33884
rect 24302 33872 24308 33884
rect 24360 33872 24366 33924
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1946 33844 1952 33856
rect 1443 33816 1952 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1946 33804 1952 33816
rect 2004 33804 2010 33856
rect 20714 33804 20720 33856
rect 20772 33844 20778 33856
rect 24504 33844 24532 33943
rect 25406 33912 25412 33924
rect 25367 33884 25412 33912
rect 25406 33872 25412 33884
rect 25464 33872 25470 33924
rect 26418 33872 26424 33924
rect 26476 33872 26482 33924
rect 27246 33872 27252 33924
rect 27304 33912 27310 33924
rect 27341 33915 27399 33921
rect 27341 33912 27353 33915
rect 27304 33884 27353 33912
rect 27304 33872 27310 33884
rect 27341 33881 27353 33884
rect 27387 33881 27399 33915
rect 27341 33875 27399 33881
rect 27430 33872 27436 33924
rect 27488 33912 27494 33924
rect 27632 33912 27660 33943
rect 29178 33940 29184 33952
rect 29236 33980 29242 33992
rect 29730 33980 29736 33992
rect 29236 33952 29736 33980
rect 29236 33940 29242 33952
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 29917 33983 29975 33989
rect 29917 33949 29929 33983
rect 29963 33980 29975 33983
rect 30006 33980 30012 33992
rect 29963 33952 30012 33980
rect 29963 33949 29975 33952
rect 29917 33943 29975 33949
rect 30006 33940 30012 33952
rect 30064 33940 30070 33992
rect 30098 33940 30104 33992
rect 30156 33980 30162 33992
rect 30156 33952 30201 33980
rect 30156 33940 30162 33952
rect 30282 33940 30288 33992
rect 30340 33980 30346 33992
rect 30340 33952 30385 33980
rect 30340 33940 30346 33952
rect 30466 33940 30472 33992
rect 30524 33980 30530 33992
rect 32953 33983 33011 33989
rect 30524 33952 30569 33980
rect 30524 33940 30530 33952
rect 32953 33949 32965 33983
rect 32999 33980 33011 33983
rect 33873 33983 33931 33989
rect 32999 33952 33456 33980
rect 32999 33949 33011 33952
rect 32953 33943 33011 33949
rect 31110 33912 31116 33924
rect 27488 33884 31116 33912
rect 27488 33872 27494 33884
rect 31110 33872 31116 33884
rect 31168 33872 31174 33924
rect 26326 33844 26332 33856
rect 20772 33816 20817 33844
rect 24504 33816 26332 33844
rect 20772 33804 20778 33816
rect 26326 33804 26332 33816
rect 26384 33844 26390 33856
rect 26881 33847 26939 33853
rect 26881 33844 26893 33847
rect 26384 33816 26893 33844
rect 26384 33804 26390 33816
rect 26881 33813 26893 33816
rect 26927 33813 26939 33847
rect 26881 33807 26939 33813
rect 28997 33847 29055 33853
rect 28997 33813 29009 33847
rect 29043 33844 29055 33847
rect 29546 33844 29552 33856
rect 29043 33816 29552 33844
rect 29043 33813 29055 33816
rect 28997 33807 29055 33813
rect 29546 33804 29552 33816
rect 29604 33804 29610 33856
rect 30653 33847 30711 33853
rect 30653 33813 30665 33847
rect 30699 33844 30711 33847
rect 31294 33844 31300 33856
rect 30699 33816 31300 33844
rect 30699 33813 30711 33816
rect 30653 33807 30711 33813
rect 31294 33804 31300 33816
rect 31352 33804 31358 33856
rect 32766 33844 32772 33856
rect 32727 33816 32772 33844
rect 32766 33804 32772 33816
rect 32824 33804 32830 33856
rect 33428 33853 33456 33952
rect 33873 33949 33885 33983
rect 33919 33980 33931 33983
rect 34514 33980 34520 33992
rect 33919 33952 34520 33980
rect 33919 33949 33931 33952
rect 33873 33943 33931 33949
rect 34514 33940 34520 33952
rect 34572 33940 34578 33992
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34664 33952 34713 33980
rect 34664 33940 34670 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 34885 33983 34943 33989
rect 34885 33980 34897 33983
rect 34848 33952 34897 33980
rect 34848 33940 34854 33952
rect 34885 33949 34897 33952
rect 34931 33980 34943 33983
rect 35158 33980 35164 33992
rect 34931 33952 35164 33980
rect 34931 33949 34943 33952
rect 34885 33943 34943 33949
rect 35158 33940 35164 33952
rect 35216 33940 35222 33992
rect 33781 33915 33839 33921
rect 33781 33881 33793 33915
rect 33827 33912 33839 33915
rect 34808 33912 34836 33940
rect 33827 33884 34836 33912
rect 33827 33881 33839 33884
rect 33781 33875 33839 33881
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 33413 33847 33471 33853
rect 33413 33813 33425 33847
rect 33459 33813 33471 33847
rect 33413 33807 33471 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 19058 33600 19064 33652
rect 19116 33640 19122 33652
rect 20714 33640 20720 33652
rect 19116 33612 20720 33640
rect 19116 33600 19122 33612
rect 20714 33600 20720 33612
rect 20772 33600 20778 33652
rect 22738 33600 22744 33652
rect 22796 33640 22802 33652
rect 23477 33643 23535 33649
rect 23477 33640 23489 33643
rect 22796 33612 23489 33640
rect 22796 33600 22802 33612
rect 23477 33609 23489 33612
rect 23523 33609 23535 33643
rect 23477 33603 23535 33609
rect 23750 33600 23756 33652
rect 23808 33600 23814 33652
rect 23842 33600 23848 33652
rect 23900 33640 23906 33652
rect 24210 33640 24216 33652
rect 23900 33612 24216 33640
rect 23900 33600 23906 33612
rect 24210 33600 24216 33612
rect 24268 33600 24274 33652
rect 29178 33640 29184 33652
rect 28644 33612 29184 33640
rect 22833 33575 22891 33581
rect 22833 33541 22845 33575
rect 22879 33572 22891 33575
rect 23566 33572 23572 33584
rect 22879 33544 23572 33572
rect 22879 33541 22891 33544
rect 22833 33535 22891 33541
rect 23566 33532 23572 33544
rect 23624 33532 23630 33584
rect 14366 33464 14372 33516
rect 14424 33504 14430 33516
rect 20441 33507 20499 33513
rect 20441 33504 20453 33507
rect 14424 33476 20453 33504
rect 14424 33464 14430 33476
rect 20441 33473 20453 33476
rect 20487 33473 20499 33507
rect 20441 33467 20499 33473
rect 20533 33507 20591 33513
rect 20533 33473 20545 33507
rect 20579 33504 20591 33507
rect 20990 33504 20996 33516
rect 20579 33476 20996 33504
rect 20579 33473 20591 33476
rect 20533 33467 20591 33473
rect 20990 33464 20996 33476
rect 21048 33464 21054 33516
rect 23658 33504 23664 33516
rect 23619 33476 23664 33504
rect 23658 33464 23664 33476
rect 23716 33464 23722 33516
rect 23768 33513 23796 33600
rect 27157 33575 27215 33581
rect 27157 33541 27169 33575
rect 27203 33572 27215 33575
rect 27338 33572 27344 33584
rect 27203 33544 27344 33572
rect 27203 33541 27215 33544
rect 27157 33535 27215 33541
rect 27338 33532 27344 33544
rect 27396 33532 27402 33584
rect 28644 33581 28672 33612
rect 29178 33600 29184 33612
rect 29236 33600 29242 33652
rect 30006 33640 30012 33652
rect 29967 33612 30012 33640
rect 30006 33600 30012 33612
rect 30064 33600 30070 33652
rect 35158 33640 35164 33652
rect 35119 33612 35164 33640
rect 35158 33600 35164 33612
rect 35216 33600 35222 33652
rect 47762 33600 47768 33652
rect 47820 33640 47826 33652
rect 48041 33643 48099 33649
rect 48041 33640 48053 33643
rect 47820 33612 48053 33640
rect 47820 33600 47826 33612
rect 48041 33609 48053 33612
rect 48087 33609 48099 33643
rect 48041 33603 48099 33609
rect 28629 33575 28687 33581
rect 28629 33541 28641 33575
rect 28675 33541 28687 33575
rect 28629 33535 28687 33541
rect 28813 33575 28871 33581
rect 28813 33541 28825 33575
rect 28859 33572 28871 33575
rect 28902 33572 28908 33584
rect 28859 33544 28908 33572
rect 28859 33541 28871 33544
rect 28813 33535 28871 33541
rect 28902 33532 28908 33544
rect 28960 33532 28966 33584
rect 28997 33575 29055 33581
rect 28997 33541 29009 33575
rect 29043 33572 29055 33575
rect 29086 33572 29092 33584
rect 29043 33544 29092 33572
rect 29043 33541 29055 33544
rect 28997 33535 29055 33541
rect 29086 33532 29092 33544
rect 29144 33532 29150 33584
rect 29270 33532 29276 33584
rect 29328 33572 29334 33584
rect 31018 33572 31024 33584
rect 29328 33544 31024 33572
rect 29328 33532 29334 33544
rect 31018 33532 31024 33544
rect 31076 33572 31082 33584
rect 31076 33544 31800 33572
rect 31076 33532 31082 33544
rect 23753 33507 23811 33513
rect 23753 33473 23765 33507
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 23937 33507 23995 33513
rect 23937 33504 23949 33507
rect 23900 33476 23949 33504
rect 23900 33464 23906 33476
rect 23937 33473 23949 33476
rect 23983 33473 23995 33507
rect 23937 33467 23995 33473
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33504 24087 33507
rect 24118 33504 24124 33516
rect 24075 33476 24124 33504
rect 24075 33473 24087 33476
rect 24029 33467 24087 33473
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24670 33504 24676 33516
rect 24631 33476 24676 33504
rect 24670 33464 24676 33476
rect 24728 33464 24734 33516
rect 27430 33504 27436 33516
rect 27391 33476 27436 33504
rect 27430 33464 27436 33476
rect 27488 33464 27494 33516
rect 29104 33504 29132 33532
rect 29454 33504 29460 33516
rect 29104 33476 29460 33504
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1670 33436 1676 33448
rect 1631 33408 1676 33436
rect 1670 33396 1676 33408
rect 1728 33396 1734 33448
rect 20717 33439 20775 33445
rect 20717 33405 20729 33439
rect 20763 33436 20775 33439
rect 21082 33436 21088 33448
rect 20763 33408 21088 33436
rect 20763 33405 20775 33408
rect 20717 33399 20775 33405
rect 21082 33396 21088 33408
rect 21140 33436 21146 33448
rect 26970 33436 26976 33448
rect 21140 33408 26976 33436
rect 21140 33396 21146 33408
rect 26970 33396 26976 33408
rect 27028 33396 27034 33448
rect 27341 33439 27399 33445
rect 27341 33405 27353 33439
rect 27387 33436 27399 33439
rect 27706 33436 27712 33448
rect 27387 33408 27712 33436
rect 27387 33405 27399 33408
rect 27341 33399 27399 33405
rect 27706 33396 27712 33408
rect 27764 33436 27770 33448
rect 28442 33436 28448 33448
rect 27764 33408 28448 33436
rect 27764 33396 27770 33408
rect 28442 33396 28448 33408
rect 28500 33396 28506 33448
rect 28718 33396 28724 33448
rect 28776 33436 28782 33448
rect 29733 33439 29791 33445
rect 29733 33436 29745 33439
rect 28776 33408 29745 33436
rect 28776 33396 28782 33408
rect 29733 33405 29745 33408
rect 29779 33436 29791 33439
rect 29914 33436 29920 33448
rect 29779 33408 29920 33436
rect 29779 33405 29791 33408
rect 29733 33399 29791 33405
rect 29914 33396 29920 33408
rect 29972 33396 29978 33448
rect 31772 33436 31800 33544
rect 32766 33532 32772 33584
rect 32824 33572 32830 33584
rect 33689 33575 33747 33581
rect 33689 33572 33701 33575
rect 32824 33544 33701 33572
rect 32824 33532 32830 33544
rect 33689 33541 33701 33544
rect 33735 33541 33747 33575
rect 33689 33535 33747 33541
rect 32309 33507 32367 33513
rect 32309 33473 32321 33507
rect 32355 33504 32367 33507
rect 32490 33504 32496 33516
rect 32355 33476 32496 33504
rect 32355 33473 32367 33476
rect 32309 33467 32367 33473
rect 32490 33464 32496 33476
rect 32548 33504 32554 33516
rect 33042 33504 33048 33516
rect 32548 33476 33048 33504
rect 32548 33464 32554 33476
rect 33042 33464 33048 33476
rect 33100 33464 33106 33516
rect 34790 33464 34796 33516
rect 34848 33464 34854 33516
rect 46750 33504 46756 33516
rect 46711 33476 46756 33504
rect 46750 33464 46756 33476
rect 46808 33464 46814 33516
rect 47486 33464 47492 33516
rect 47544 33504 47550 33516
rect 47581 33507 47639 33513
rect 47581 33504 47593 33507
rect 47544 33476 47593 33504
rect 47544 33464 47550 33476
rect 47581 33473 47593 33476
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 33413 33439 33471 33445
rect 33413 33436 33425 33439
rect 31772 33408 33425 33436
rect 33413 33405 33425 33408
rect 33459 33405 33471 33439
rect 33413 33399 33471 33405
rect 20806 33328 20812 33380
rect 20864 33368 20870 33380
rect 27617 33371 27675 33377
rect 27617 33368 27629 33371
rect 20864 33340 27629 33368
rect 20864 33328 20870 33340
rect 27617 33337 27629 33340
rect 27663 33337 27675 33371
rect 31570 33368 31576 33380
rect 27617 33331 27675 33337
rect 29380 33340 31576 33368
rect 19794 33260 19800 33312
rect 19852 33300 19858 33312
rect 20073 33303 20131 33309
rect 20073 33300 20085 33303
rect 19852 33272 20085 33300
rect 19852 33260 19858 33272
rect 20073 33269 20085 33272
rect 20119 33269 20131 33303
rect 22922 33300 22928 33312
rect 22883 33272 22928 33300
rect 20073 33263 20131 33269
rect 22922 33260 22928 33272
rect 22980 33260 22986 33312
rect 23566 33260 23572 33312
rect 23624 33300 23630 33312
rect 25961 33303 26019 33309
rect 25961 33300 25973 33303
rect 23624 33272 25973 33300
rect 23624 33260 23630 33272
rect 25961 33269 25973 33272
rect 26007 33300 26019 33303
rect 26234 33300 26240 33312
rect 26007 33272 26240 33300
rect 26007 33269 26019 33272
rect 25961 33263 26019 33269
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 27154 33300 27160 33312
rect 27115 33272 27160 33300
rect 27154 33260 27160 33272
rect 27212 33300 27218 33312
rect 29380 33300 29408 33340
rect 31570 33328 31576 33340
rect 31628 33328 31634 33380
rect 31726 33340 32536 33368
rect 29546 33300 29552 33312
rect 27212 33272 29408 33300
rect 29507 33272 29552 33300
rect 27212 33260 27218 33272
rect 29546 33260 29552 33272
rect 29604 33260 29610 33312
rect 29638 33260 29644 33312
rect 29696 33300 29702 33312
rect 31726 33300 31754 33340
rect 32398 33300 32404 33312
rect 29696 33272 31754 33300
rect 32359 33272 32404 33300
rect 29696 33260 29702 33272
rect 32398 33260 32404 33272
rect 32456 33260 32462 33312
rect 32508 33300 32536 33340
rect 46937 33303 46995 33309
rect 46937 33300 46949 33303
rect 32508 33272 46949 33300
rect 46937 33269 46949 33272
rect 46983 33269 46995 33303
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 46937 33263 46995 33269
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1946 33096 1952 33108
rect 1907 33068 1952 33096
rect 1946 33056 1952 33068
rect 2004 33056 2010 33108
rect 20990 33096 20996 33108
rect 20951 33068 20996 33096
rect 20990 33056 20996 33068
rect 21048 33056 21054 33108
rect 23661 33099 23719 33105
rect 23661 33065 23673 33099
rect 23707 33096 23719 33099
rect 23842 33096 23848 33108
rect 23707 33068 23848 33096
rect 23707 33065 23719 33068
rect 23661 33059 23719 33065
rect 23842 33056 23848 33068
rect 23900 33056 23906 33108
rect 25406 33056 25412 33108
rect 25464 33096 25470 33108
rect 25593 33099 25651 33105
rect 25593 33096 25605 33099
rect 25464 33068 25605 33096
rect 25464 33056 25470 33068
rect 25593 33065 25605 33068
rect 25639 33065 25651 33099
rect 25593 33059 25651 33065
rect 26053 33099 26111 33105
rect 26053 33065 26065 33099
rect 26099 33065 26111 33099
rect 26053 33059 26111 33065
rect 26513 33099 26571 33105
rect 26513 33065 26525 33099
rect 26559 33096 26571 33099
rect 27246 33096 27252 33108
rect 26559 33068 27252 33096
rect 26559 33065 26571 33068
rect 26513 33059 26571 33065
rect 20898 32988 20904 33040
rect 20956 33028 20962 33040
rect 21913 33031 21971 33037
rect 21913 33028 21925 33031
rect 20956 33000 21925 33028
rect 20956 32988 20962 33000
rect 21913 32997 21925 33000
rect 21959 32997 21971 33031
rect 24302 33028 24308 33040
rect 21913 32991 21971 32997
rect 23860 33000 24308 33028
rect 2317 32963 2375 32969
rect 2317 32929 2329 32963
rect 2363 32929 2375 32963
rect 2317 32923 2375 32929
rect 1670 32852 1676 32904
rect 1728 32892 1734 32904
rect 1857 32895 1915 32901
rect 1857 32892 1869 32895
rect 1728 32864 1869 32892
rect 1728 32852 1734 32864
rect 1857 32861 1869 32864
rect 1903 32892 1915 32895
rect 1946 32892 1952 32904
rect 1903 32864 1952 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 1946 32852 1952 32864
rect 2004 32852 2010 32904
rect 2332 32892 2360 32923
rect 18230 32920 18236 32972
rect 18288 32960 18294 32972
rect 19794 32960 19800 32972
rect 18288 32932 19472 32960
rect 19755 32932 19800 32960
rect 18288 32920 18294 32932
rect 2961 32895 3019 32901
rect 2961 32892 2973 32895
rect 2332 32864 2973 32892
rect 2961 32861 2973 32864
rect 3007 32861 3019 32895
rect 2961 32855 3019 32861
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32892 18751 32895
rect 18739 32864 19380 32892
rect 18739 32861 18751 32864
rect 18693 32855 18751 32861
rect 2222 32716 2228 32768
rect 2280 32756 2286 32768
rect 2777 32759 2835 32765
rect 2777 32756 2789 32759
rect 2280 32728 2789 32756
rect 2280 32716 2286 32728
rect 2777 32725 2789 32728
rect 2823 32725 2835 32759
rect 2777 32719 2835 32725
rect 18138 32716 18144 32768
rect 18196 32756 18202 32768
rect 19352 32765 19380 32864
rect 18509 32759 18567 32765
rect 18509 32756 18521 32759
rect 18196 32728 18521 32756
rect 18196 32716 18202 32728
rect 18509 32725 18521 32728
rect 18555 32725 18567 32759
rect 18509 32719 18567 32725
rect 19337 32759 19395 32765
rect 19337 32725 19349 32759
rect 19383 32725 19395 32759
rect 19444 32756 19472 32932
rect 19794 32920 19800 32932
rect 19852 32920 19858 32972
rect 19981 32963 20039 32969
rect 19981 32929 19993 32963
rect 20027 32960 20039 32963
rect 20070 32960 20076 32972
rect 20027 32932 20076 32960
rect 20027 32929 20039 32932
rect 19981 32923 20039 32929
rect 20070 32920 20076 32932
rect 20128 32920 20134 32972
rect 20809 32963 20867 32969
rect 20809 32929 20821 32963
rect 20855 32960 20867 32963
rect 21450 32960 21456 32972
rect 20855 32932 21456 32960
rect 20855 32929 20867 32932
rect 20809 32923 20867 32929
rect 21450 32920 21456 32932
rect 21508 32920 21514 32972
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32892 19763 32895
rect 20530 32892 20536 32904
rect 19751 32864 20536 32892
rect 19751 32861 19763 32864
rect 19705 32855 19763 32861
rect 20530 32852 20536 32864
rect 20588 32892 20594 32904
rect 20717 32895 20775 32901
rect 20717 32892 20729 32895
rect 20588 32864 20729 32892
rect 20588 32852 20594 32864
rect 20717 32861 20729 32864
rect 20763 32892 20775 32895
rect 21545 32895 21603 32901
rect 21545 32892 21557 32895
rect 20763 32864 21557 32892
rect 20763 32861 20775 32864
rect 20717 32855 20775 32861
rect 21545 32861 21557 32864
rect 21591 32861 21603 32895
rect 23658 32892 23664 32904
rect 23619 32864 23664 32892
rect 21545 32855 21603 32861
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 23860 32901 23888 33000
rect 24302 32988 24308 33000
rect 24360 33028 24366 33040
rect 26068 33028 26096 33059
rect 27246 33056 27252 33068
rect 27304 33056 27310 33108
rect 27522 33056 27528 33108
rect 27580 33096 27586 33108
rect 27617 33099 27675 33105
rect 27617 33096 27629 33099
rect 27580 33068 27629 33096
rect 27580 33056 27586 33068
rect 27617 33065 27629 33068
rect 27663 33065 27675 33099
rect 27617 33059 27675 33065
rect 28629 33099 28687 33105
rect 28629 33065 28641 33099
rect 28675 33096 28687 33099
rect 29178 33096 29184 33108
rect 28675 33068 29184 33096
rect 28675 33065 28687 33068
rect 28629 33059 28687 33065
rect 29178 33056 29184 33068
rect 29236 33056 29242 33108
rect 31110 33056 31116 33108
rect 31168 33096 31174 33108
rect 32769 33099 32827 33105
rect 32769 33096 32781 33099
rect 31168 33068 32781 33096
rect 31168 33056 31174 33068
rect 32769 33065 32781 33068
rect 32815 33065 32827 33099
rect 34790 33096 34796 33108
rect 34751 33068 34796 33096
rect 32769 33059 32827 33065
rect 34790 33056 34796 33068
rect 34848 33056 34854 33108
rect 24360 33000 26096 33028
rect 24360 32988 24366 33000
rect 27338 32988 27344 33040
rect 27396 33028 27402 33040
rect 29638 33028 29644 33040
rect 27396 33000 29644 33028
rect 27396 32988 27402 33000
rect 29638 32988 29644 33000
rect 29696 32988 29702 33040
rect 25225 32963 25283 32969
rect 25225 32929 25237 32963
rect 25271 32960 25283 32963
rect 25314 32960 25320 32972
rect 25271 32932 25320 32960
rect 25271 32929 25283 32932
rect 25225 32923 25283 32929
rect 25314 32920 25320 32932
rect 25372 32960 25378 32972
rect 25869 32963 25927 32969
rect 25869 32960 25881 32963
rect 25372 32932 25881 32960
rect 25372 32920 25378 32932
rect 25869 32929 25881 32932
rect 25915 32929 25927 32963
rect 25869 32923 25927 32929
rect 25958 32920 25964 32972
rect 26016 32960 26022 32972
rect 26145 32963 26203 32969
rect 26145 32960 26157 32963
rect 26016 32932 26157 32960
rect 26016 32920 26022 32932
rect 26145 32929 26157 32932
rect 26191 32929 26203 32963
rect 26145 32923 26203 32929
rect 28258 32920 28264 32972
rect 28316 32960 28322 32972
rect 28316 32932 29684 32960
rect 28316 32920 28322 32932
rect 23845 32895 23903 32901
rect 23845 32861 23857 32895
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 24946 32892 24952 32904
rect 24903 32864 24952 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 24946 32852 24952 32864
rect 25004 32852 25010 32904
rect 25041 32895 25099 32901
rect 25041 32861 25053 32895
rect 25087 32861 25099 32895
rect 25041 32855 25099 32861
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25406 32892 25412 32904
rect 25367 32864 25412 32892
rect 25133 32855 25191 32861
rect 20346 32784 20352 32836
rect 20404 32824 20410 32836
rect 21729 32827 21787 32833
rect 21729 32824 21741 32827
rect 20404 32796 21741 32824
rect 20404 32784 20410 32796
rect 21729 32793 21741 32796
rect 21775 32793 21787 32827
rect 21729 32787 21787 32793
rect 22830 32784 22836 32836
rect 22888 32824 22894 32836
rect 23014 32824 23020 32836
rect 22888 32796 23020 32824
rect 22888 32784 22894 32796
rect 23014 32784 23020 32796
rect 23072 32824 23078 32836
rect 25056 32824 25084 32855
rect 23072 32796 25084 32824
rect 25148 32824 25176 32855
rect 25406 32852 25412 32864
rect 25464 32852 25470 32904
rect 26326 32892 26332 32904
rect 25516 32864 26332 32892
rect 25516 32824 25544 32864
rect 26326 32852 26332 32864
rect 26384 32852 26390 32904
rect 27433 32895 27491 32901
rect 27433 32861 27445 32895
rect 27479 32892 27491 32895
rect 27982 32892 27988 32904
rect 27479 32864 27988 32892
rect 27479 32861 27491 32864
rect 27433 32855 27491 32861
rect 27982 32852 27988 32864
rect 28040 32852 28046 32904
rect 28442 32892 28448 32904
rect 28403 32864 28448 32892
rect 28442 32852 28448 32864
rect 28500 32852 28506 32904
rect 28534 32852 28540 32904
rect 28592 32892 28598 32904
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28592 32864 28641 32892
rect 28592 32852 28598 32864
rect 28629 32861 28641 32864
rect 28675 32892 28687 32895
rect 28902 32892 28908 32904
rect 28675 32864 28908 32892
rect 28675 32861 28687 32864
rect 28629 32855 28687 32861
rect 28902 32852 28908 32864
rect 28960 32852 28966 32904
rect 29454 32852 29460 32904
rect 29512 32892 29518 32904
rect 29656 32901 29684 32932
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 29825 32963 29883 32969
rect 29825 32960 29837 32963
rect 29788 32932 29837 32960
rect 29788 32920 29794 32932
rect 29825 32929 29837 32932
rect 29871 32929 29883 32963
rect 31018 32960 31024 32972
rect 30979 32932 31024 32960
rect 29825 32923 29883 32929
rect 31018 32920 31024 32932
rect 31076 32920 31082 32972
rect 31294 32960 31300 32972
rect 31255 32932 31300 32960
rect 31294 32920 31300 32932
rect 31352 32920 31358 32972
rect 29549 32895 29607 32901
rect 29549 32892 29561 32895
rect 29512 32864 29561 32892
rect 29512 32852 29518 32864
rect 29549 32861 29561 32864
rect 29595 32861 29607 32895
rect 29549 32855 29607 32861
rect 29641 32895 29699 32901
rect 29641 32861 29653 32895
rect 29687 32892 29699 32895
rect 30374 32892 30380 32904
rect 29687 32864 30380 32892
rect 29687 32861 29699 32864
rect 29641 32855 29699 32861
rect 30374 32852 30380 32864
rect 30432 32852 30438 32904
rect 32398 32852 32404 32904
rect 32456 32852 32462 32904
rect 33042 32852 33048 32904
rect 33100 32892 33106 32904
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 33100 32864 34713 32892
rect 33100 32852 33106 32864
rect 34701 32861 34713 32864
rect 34747 32892 34759 32895
rect 35710 32892 35716 32904
rect 34747 32864 35716 32892
rect 34747 32861 34759 32864
rect 34701 32855 34759 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 45833 32895 45891 32901
rect 45833 32861 45845 32895
rect 45879 32892 45891 32895
rect 46293 32895 46351 32901
rect 46293 32892 46305 32895
rect 45879 32864 46305 32892
rect 45879 32861 45891 32864
rect 45833 32855 45891 32861
rect 46293 32861 46305 32864
rect 46339 32861 46351 32895
rect 46293 32855 46351 32861
rect 25148 32796 25544 32824
rect 26053 32827 26111 32833
rect 23072 32784 23078 32796
rect 26053 32793 26065 32827
rect 26099 32824 26111 32827
rect 26142 32824 26148 32836
rect 26099 32796 26148 32824
rect 26099 32793 26111 32796
rect 26053 32787 26111 32793
rect 26142 32784 26148 32796
rect 26200 32784 26206 32836
rect 27522 32784 27528 32836
rect 27580 32824 27586 32836
rect 31386 32824 31392 32836
rect 27580 32796 31392 32824
rect 27580 32784 27586 32796
rect 31386 32784 31392 32796
rect 31444 32784 31450 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 46934 32824 46940 32836
rect 46523 32796 46940 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 46934 32784 46940 32796
rect 46992 32784 46998 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 23290 32756 23296 32768
rect 19444 32728 23296 32756
rect 19337 32719 19395 32725
rect 23290 32716 23296 32728
rect 23348 32756 23354 32768
rect 25406 32756 25412 32768
rect 23348 32728 25412 32756
rect 23348 32716 23354 32728
rect 25406 32716 25412 32728
rect 25464 32716 25470 32768
rect 25498 32716 25504 32768
rect 25556 32756 25562 32768
rect 28813 32759 28871 32765
rect 28813 32756 28825 32759
rect 25556 32728 28825 32756
rect 25556 32716 25562 32728
rect 28813 32725 28825 32728
rect 28859 32725 28871 32759
rect 28813 32719 28871 32725
rect 29546 32716 29552 32768
rect 29604 32756 29610 32768
rect 29825 32759 29883 32765
rect 29825 32756 29837 32759
rect 29604 32728 29837 32756
rect 29604 32716 29610 32728
rect 29825 32725 29837 32728
rect 29871 32725 29883 32759
rect 29825 32719 29883 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 3786 32512 3792 32564
rect 3844 32552 3850 32564
rect 3844 32524 22094 32552
rect 3844 32512 3850 32524
rect 2222 32484 2228 32496
rect 2183 32456 2228 32484
rect 2222 32444 2228 32456
rect 2280 32444 2286 32496
rect 18138 32484 18144 32496
rect 18099 32456 18144 32484
rect 18138 32444 18144 32456
rect 18196 32444 18202 32496
rect 22066 32484 22094 32524
rect 23658 32512 23664 32564
rect 23716 32552 23722 32564
rect 25041 32555 25099 32561
rect 25041 32552 25053 32555
rect 23716 32524 25053 32552
rect 23716 32512 23722 32524
rect 25041 32521 25053 32524
rect 25087 32521 25099 32555
rect 26329 32555 26387 32561
rect 25041 32515 25099 32521
rect 25148 32524 26280 32552
rect 25148 32484 25176 32524
rect 25958 32484 25964 32496
rect 22066 32456 25176 32484
rect 25608 32456 25964 32484
rect 1854 32376 1860 32428
rect 1912 32416 1918 32428
rect 2041 32419 2099 32425
rect 2041 32416 2053 32419
rect 1912 32388 2053 32416
rect 1912 32376 1918 32388
rect 2041 32385 2053 32388
rect 2087 32385 2099 32419
rect 2041 32379 2099 32385
rect 19242 32376 19248 32428
rect 19300 32376 19306 32428
rect 20257 32419 20315 32425
rect 20257 32416 20269 32419
rect 19352 32388 20269 32416
rect 3881 32351 3939 32357
rect 3881 32317 3893 32351
rect 3927 32348 3939 32351
rect 4614 32348 4620 32360
rect 3927 32320 4620 32348
rect 3927 32317 3939 32320
rect 3881 32311 3939 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32317 17923 32351
rect 17865 32311 17923 32317
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 1452 32184 1593 32212
rect 1452 32172 1458 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 1581 32175 1639 32181
rect 7466 32172 7472 32224
rect 7524 32212 7530 32224
rect 17678 32212 17684 32224
rect 7524 32184 17684 32212
rect 7524 32172 7530 32184
rect 17678 32172 17684 32184
rect 17736 32172 17742 32224
rect 17880 32212 17908 32311
rect 19150 32308 19156 32360
rect 19208 32348 19214 32360
rect 19352 32348 19380 32388
rect 20257 32385 20269 32388
rect 20303 32416 20315 32419
rect 20346 32416 20352 32428
rect 20303 32388 20352 32416
rect 20303 32385 20315 32388
rect 20257 32379 20315 32385
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 20530 32416 20536 32428
rect 20491 32388 20536 32416
rect 20530 32376 20536 32388
rect 20588 32376 20594 32428
rect 20898 32376 20904 32428
rect 20956 32416 20962 32428
rect 20993 32419 21051 32425
rect 20993 32416 21005 32419
rect 20956 32388 21005 32416
rect 20956 32376 20962 32388
rect 20993 32385 21005 32388
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32416 21235 32419
rect 21450 32416 21456 32428
rect 21223 32388 21456 32416
rect 21223 32385 21235 32388
rect 21177 32379 21235 32385
rect 19208 32320 19380 32348
rect 19613 32351 19671 32357
rect 19208 32308 19214 32320
rect 19613 32317 19625 32351
rect 19659 32348 19671 32351
rect 20548 32348 20576 32376
rect 19659 32320 20576 32348
rect 19659 32317 19671 32320
rect 19613 32311 19671 32317
rect 20441 32283 20499 32289
rect 20441 32249 20453 32283
rect 20487 32280 20499 32283
rect 21192 32280 21220 32379
rect 21450 32376 21456 32388
rect 21508 32376 21514 32428
rect 24026 32376 24032 32428
rect 24084 32416 24090 32428
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 24084 32388 24685 32416
rect 24084 32376 24090 32388
rect 24673 32385 24685 32388
rect 24719 32416 24731 32419
rect 25498 32416 25504 32428
rect 24719 32388 25504 32416
rect 24719 32385 24731 32388
rect 24673 32379 24731 32385
rect 25498 32376 25504 32388
rect 25556 32376 25562 32428
rect 24578 32308 24584 32360
rect 24636 32348 24642 32360
rect 24765 32351 24823 32357
rect 24765 32348 24777 32351
rect 24636 32320 24777 32348
rect 24636 32308 24642 32320
rect 24765 32317 24777 32320
rect 24811 32348 24823 32351
rect 25608 32348 25636 32456
rect 25958 32444 25964 32456
rect 26016 32444 26022 32496
rect 26252 32484 26280 32524
rect 26329 32521 26341 32555
rect 26375 32552 26387 32555
rect 28350 32552 28356 32564
rect 26375 32524 28356 32552
rect 26375 32521 26387 32524
rect 26329 32515 26387 32521
rect 28350 32512 28356 32524
rect 28408 32512 28414 32564
rect 28442 32512 28448 32564
rect 28500 32552 28506 32564
rect 28902 32552 28908 32564
rect 28500 32524 28908 32552
rect 28500 32512 28506 32524
rect 28902 32512 28908 32524
rect 28960 32512 28966 32564
rect 28994 32512 29000 32564
rect 29052 32552 29058 32564
rect 32858 32552 32864 32564
rect 29052 32524 32864 32552
rect 29052 32512 29058 32524
rect 32858 32512 32864 32524
rect 32916 32512 32922 32564
rect 46934 32552 46940 32564
rect 46895 32524 46940 32552
rect 46934 32512 46940 32524
rect 46992 32512 46998 32564
rect 29454 32484 29460 32496
rect 26252 32456 29460 32484
rect 29454 32444 29460 32456
rect 29512 32444 29518 32496
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32416 25743 32419
rect 26142 32416 26148 32428
rect 25731 32388 26148 32416
rect 25731 32385 25743 32388
rect 25685 32379 25743 32385
rect 24811 32320 25636 32348
rect 24811 32317 24823 32320
rect 24765 32311 24823 32317
rect 25700 32280 25728 32379
rect 26142 32376 26148 32388
rect 26200 32376 26206 32428
rect 26234 32376 26240 32428
rect 26292 32416 26298 32428
rect 27430 32416 27436 32428
rect 26292 32388 26337 32416
rect 27391 32388 27436 32416
rect 26292 32376 26298 32388
rect 27430 32376 27436 32388
rect 27488 32376 27494 32428
rect 28258 32376 28264 32428
rect 28316 32416 28322 32428
rect 28353 32419 28411 32425
rect 28353 32416 28365 32419
rect 28316 32388 28365 32416
rect 28316 32376 28322 32388
rect 28353 32385 28365 32388
rect 28399 32385 28411 32419
rect 28353 32379 28411 32385
rect 28629 32419 28687 32425
rect 28629 32385 28641 32419
rect 28675 32416 28687 32419
rect 29730 32416 29736 32428
rect 28675 32388 29736 32416
rect 28675 32385 28687 32388
rect 28629 32379 28687 32385
rect 29730 32376 29736 32388
rect 29788 32376 29794 32428
rect 30926 32376 30932 32428
rect 30984 32416 30990 32428
rect 31021 32419 31079 32425
rect 31021 32416 31033 32419
rect 30984 32388 31033 32416
rect 30984 32376 30990 32388
rect 31021 32385 31033 32388
rect 31067 32385 31079 32419
rect 31021 32379 31079 32385
rect 31386 32376 31392 32428
rect 31444 32416 31450 32428
rect 32125 32419 32183 32425
rect 32125 32416 32137 32419
rect 31444 32388 32137 32416
rect 31444 32376 31450 32388
rect 32125 32385 32137 32388
rect 32171 32385 32183 32419
rect 32125 32379 32183 32385
rect 46474 32376 46480 32428
rect 46532 32416 46538 32428
rect 46845 32419 46903 32425
rect 46845 32416 46857 32419
rect 46532 32388 46857 32416
rect 46532 32376 46538 32388
rect 46845 32385 46857 32388
rect 46891 32416 46903 32419
rect 47394 32416 47400 32428
rect 46891 32388 47400 32416
rect 46891 32385 46903 32388
rect 46845 32379 46903 32385
rect 47394 32376 47400 32388
rect 47452 32376 47458 32428
rect 47946 32416 47952 32428
rect 47907 32388 47952 32416
rect 47946 32376 47952 32388
rect 48004 32376 48010 32428
rect 28537 32351 28595 32357
rect 28537 32317 28549 32351
rect 28583 32348 28595 32351
rect 29178 32348 29184 32360
rect 28583 32320 29184 32348
rect 28583 32317 28595 32320
rect 28537 32311 28595 32317
rect 29178 32308 29184 32320
rect 29236 32308 29242 32360
rect 29822 32348 29828 32360
rect 29783 32320 29828 32348
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 29914 32308 29920 32360
rect 29972 32348 29978 32360
rect 29972 32320 30017 32348
rect 29972 32308 29978 32320
rect 20487 32252 21220 32280
rect 24872 32252 25728 32280
rect 20487 32249 20499 32252
rect 20441 32243 20499 32249
rect 18874 32212 18880 32224
rect 17880 32184 18880 32212
rect 18874 32172 18880 32184
rect 18932 32172 18938 32224
rect 20070 32212 20076 32224
rect 20031 32184 20076 32212
rect 20070 32172 20076 32184
rect 20128 32172 20134 32224
rect 20990 32212 20996 32224
rect 20951 32184 20996 32212
rect 20990 32172 20996 32184
rect 21048 32172 21054 32224
rect 24210 32172 24216 32224
rect 24268 32212 24274 32224
rect 24872 32221 24900 32252
rect 25774 32240 25780 32292
rect 25832 32280 25838 32292
rect 48133 32283 48191 32289
rect 48133 32280 48145 32283
rect 25832 32252 48145 32280
rect 25832 32240 25838 32252
rect 48133 32249 48145 32252
rect 48179 32249 48191 32283
rect 48133 32243 48191 32249
rect 24857 32215 24915 32221
rect 24857 32212 24869 32215
rect 24268 32184 24869 32212
rect 24268 32172 24274 32184
rect 24857 32181 24869 32184
rect 24903 32181 24915 32215
rect 25498 32212 25504 32224
rect 25459 32184 25504 32212
rect 24857 32175 24915 32181
rect 25498 32172 25504 32184
rect 25556 32172 25562 32224
rect 25590 32172 25596 32224
rect 25648 32212 25654 32224
rect 27617 32215 27675 32221
rect 27617 32212 27629 32215
rect 25648 32184 27629 32212
rect 25648 32172 25654 32184
rect 27617 32181 27629 32184
rect 27663 32181 27675 32215
rect 28534 32212 28540 32224
rect 28495 32184 28540 32212
rect 27617 32175 27675 32181
rect 28534 32172 28540 32184
rect 28592 32172 28598 32224
rect 28813 32215 28871 32221
rect 28813 32181 28825 32215
rect 28859 32212 28871 32215
rect 29178 32212 29184 32224
rect 28859 32184 29184 32212
rect 28859 32181 28871 32184
rect 28813 32175 28871 32181
rect 29178 32172 29184 32184
rect 29236 32172 29242 32224
rect 29365 32215 29423 32221
rect 29365 32181 29377 32215
rect 29411 32212 29423 32215
rect 30742 32212 30748 32224
rect 29411 32184 30748 32212
rect 29411 32181 29423 32184
rect 29365 32175 29423 32181
rect 30742 32172 30748 32184
rect 30800 32172 30806 32224
rect 31113 32215 31171 32221
rect 31113 32181 31125 32215
rect 31159 32212 31171 32215
rect 31478 32212 31484 32224
rect 31159 32184 31484 32212
rect 31159 32181 31171 32184
rect 31113 32175 31171 32181
rect 31478 32172 31484 32184
rect 31536 32172 31542 32224
rect 32030 32172 32036 32224
rect 32088 32212 32094 32224
rect 32309 32215 32367 32221
rect 32309 32212 32321 32215
rect 32088 32184 32321 32212
rect 32088 32172 32094 32184
rect 32309 32181 32321 32184
rect 32355 32181 32367 32215
rect 32309 32175 32367 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 3878 31968 3884 32020
rect 3936 32008 3942 32020
rect 3936 31980 15332 32008
rect 3936 31968 3942 31980
rect 1946 31900 1952 31952
rect 2004 31940 2010 31952
rect 2004 31912 3924 31940
rect 2004 31900 2010 31912
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 3786 31872 3792 31884
rect 3747 31844 3792 31872
rect 3786 31832 3792 31844
rect 3844 31832 3850 31884
rect 3896 31872 3924 31912
rect 8294 31900 8300 31952
rect 8352 31940 8358 31952
rect 8352 31912 12480 31940
rect 8352 31900 8358 31912
rect 3973 31875 4031 31881
rect 3973 31872 3985 31875
rect 3896 31844 3985 31872
rect 3973 31841 3985 31844
rect 4019 31841 4031 31875
rect 4614 31872 4620 31884
rect 4575 31844 4620 31872
rect 3973 31835 4031 31841
rect 4614 31832 4620 31844
rect 4672 31872 4678 31884
rect 5442 31872 5448 31884
rect 4672 31844 5448 31872
rect 4672 31832 4678 31844
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 12452 31881 12480 31912
rect 12437 31875 12495 31881
rect 12437 31841 12449 31875
rect 12483 31841 12495 31875
rect 12437 31835 12495 31841
rect 14829 31875 14887 31881
rect 14829 31841 14841 31875
rect 14875 31872 14887 31875
rect 15194 31872 15200 31884
rect 14875 31844 15200 31872
rect 14875 31841 14887 31844
rect 14829 31835 14887 31841
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 15304 31881 15332 31980
rect 19242 31968 19248 32020
rect 19300 32008 19306 32020
rect 19337 32011 19395 32017
rect 19337 32008 19349 32011
rect 19300 31980 19349 32008
rect 19300 31968 19306 31980
rect 19337 31977 19349 31980
rect 19383 31977 19395 32011
rect 19337 31971 19395 31977
rect 20070 31968 20076 32020
rect 20128 32008 20134 32020
rect 20441 32011 20499 32017
rect 20441 32008 20453 32011
rect 20128 31980 20453 32008
rect 20128 31968 20134 31980
rect 20441 31977 20453 31980
rect 20487 31977 20499 32011
rect 24118 32008 24124 32020
rect 20441 31971 20499 31977
rect 21284 31980 24124 32008
rect 20809 31943 20867 31949
rect 20809 31940 20821 31943
rect 17604 31912 20821 31940
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31841 15347 31875
rect 15289 31835 15347 31841
rect 11698 31804 11704 31816
rect 11659 31776 11704 31804
rect 11698 31764 11704 31776
rect 11756 31764 11762 31816
rect 17604 31813 17632 31912
rect 20809 31909 20821 31912
rect 20855 31909 20867 31943
rect 20809 31903 20867 31909
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 17957 31875 18015 31881
rect 17957 31872 17969 31875
rect 17736 31844 17969 31872
rect 17736 31832 17742 31844
rect 17957 31841 17969 31844
rect 18003 31841 18015 31875
rect 19150 31872 19156 31884
rect 17957 31835 18015 31841
rect 18064 31844 19156 31872
rect 17589 31807 17647 31813
rect 17589 31773 17601 31807
rect 17635 31773 17647 31807
rect 17770 31804 17776 31816
rect 17731 31776 17776 31804
rect 17589 31767 17647 31773
rect 17770 31764 17776 31776
rect 17828 31764 17834 31816
rect 17865 31807 17923 31813
rect 17865 31773 17877 31807
rect 17911 31804 17923 31807
rect 18064 31804 18092 31844
rect 19150 31832 19156 31844
rect 19208 31832 19214 31884
rect 19426 31872 19432 31884
rect 19260 31844 19432 31872
rect 17911 31776 18092 31804
rect 18141 31807 18199 31813
rect 17911 31773 17923 31776
rect 17865 31767 17923 31773
rect 18141 31773 18153 31807
rect 18187 31804 18199 31807
rect 18230 31804 18236 31816
rect 18187 31776 18236 31804
rect 18187 31773 18199 31776
rect 18141 31767 18199 31773
rect 18230 31764 18236 31776
rect 18288 31764 18294 31816
rect 19260 31813 19288 31844
rect 19426 31832 19432 31844
rect 19484 31832 19490 31884
rect 21284 31872 21312 31980
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 26970 31968 26976 32020
rect 27028 32008 27034 32020
rect 27249 32011 27307 32017
rect 27249 32008 27261 32011
rect 27028 31980 27261 32008
rect 27028 31968 27034 31980
rect 27249 31977 27261 31980
rect 27295 31977 27307 32011
rect 27249 31971 27307 31977
rect 28813 32011 28871 32017
rect 28813 31977 28825 32011
rect 28859 32008 28871 32011
rect 29730 32008 29736 32020
rect 28859 31980 29736 32008
rect 28859 31977 28871 31980
rect 28813 31971 28871 31977
rect 29730 31968 29736 31980
rect 29788 32008 29794 32020
rect 31849 32011 31907 32017
rect 31849 32008 31861 32011
rect 29788 31980 31861 32008
rect 29788 31968 29794 31980
rect 31849 31977 31861 31980
rect 31895 31977 31907 32011
rect 31849 31971 31907 31977
rect 41690 31968 41696 32020
rect 41748 32008 41754 32020
rect 47578 32008 47584 32020
rect 41748 31980 47584 32008
rect 41748 31968 41754 31980
rect 47578 31968 47584 31980
rect 47636 31968 47642 32020
rect 23753 31943 23811 31949
rect 23753 31909 23765 31943
rect 23799 31940 23811 31943
rect 24578 31940 24584 31952
rect 23799 31912 24584 31940
rect 23799 31909 23811 31912
rect 23753 31903 23811 31909
rect 24578 31900 24584 31912
rect 24636 31900 24642 31952
rect 24762 31900 24768 31952
rect 24820 31940 24826 31952
rect 26513 31943 26571 31949
rect 26513 31940 26525 31943
rect 24820 31912 26525 31940
rect 24820 31900 24826 31912
rect 26513 31909 26525 31912
rect 26559 31940 26571 31943
rect 27890 31940 27896 31952
rect 26559 31912 27896 31940
rect 26559 31909 26571 31912
rect 26513 31903 26571 31909
rect 27890 31900 27896 31912
rect 27948 31940 27954 31952
rect 29914 31940 29920 31952
rect 27948 31912 29920 31940
rect 27948 31900 27954 31912
rect 29914 31900 29920 31912
rect 29972 31900 29978 31952
rect 32490 31940 32496 31952
rect 32451 31912 32496 31940
rect 32490 31900 32496 31912
rect 32548 31900 32554 31952
rect 47486 31940 47492 31952
rect 46584 31912 47492 31940
rect 22922 31872 22928 31884
rect 20456 31844 21312 31872
rect 21376 31844 22928 31872
rect 20456 31813 20484 31844
rect 19245 31807 19303 31813
rect 19245 31773 19257 31807
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31773 20499 31807
rect 20441 31767 20499 31773
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31804 20683 31807
rect 20714 31804 20720 31816
rect 20671 31776 20720 31804
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 20714 31764 20720 31776
rect 20772 31804 20778 31816
rect 20990 31804 20996 31816
rect 20772 31776 20996 31804
rect 20772 31764 20778 31776
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 21376 31813 21404 31844
rect 22922 31832 22928 31844
rect 22980 31832 22986 31884
rect 24121 31875 24179 31881
rect 24121 31841 24133 31875
rect 24167 31872 24179 31875
rect 25406 31872 25412 31884
rect 24167 31844 25412 31872
rect 24167 31841 24179 31844
rect 24121 31835 24179 31841
rect 25406 31832 25412 31844
rect 25464 31832 25470 31884
rect 25590 31832 25596 31884
rect 25648 31872 25654 31884
rect 25685 31875 25743 31881
rect 25685 31872 25697 31875
rect 25648 31844 25697 31872
rect 25648 31832 25654 31844
rect 25685 31841 25697 31844
rect 25731 31841 25743 31875
rect 25685 31835 25743 31841
rect 28258 31832 28264 31884
rect 28316 31872 28322 31884
rect 28316 31844 28764 31872
rect 28316 31832 28322 31844
rect 21361 31807 21419 31813
rect 21361 31773 21373 31807
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 21545 31807 21603 31813
rect 21545 31773 21557 31807
rect 21591 31804 21603 31807
rect 22002 31804 22008 31816
rect 21591 31776 22008 31804
rect 21591 31773 21603 31776
rect 21545 31767 21603 31773
rect 22002 31764 22008 31776
rect 22060 31764 22066 31816
rect 24026 31804 24032 31816
rect 23987 31776 24032 31804
rect 24026 31764 24032 31776
rect 24084 31764 24090 31816
rect 24210 31804 24216 31816
rect 24171 31776 24216 31804
rect 24210 31764 24216 31776
rect 24268 31764 24274 31816
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25501 31807 25559 31813
rect 25501 31804 25513 31807
rect 24903 31776 25513 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25501 31773 25513 31776
rect 25547 31804 25559 31807
rect 25774 31804 25780 31816
rect 25547 31776 25780 31804
rect 25547 31773 25559 31776
rect 25501 31767 25559 31773
rect 25774 31764 25780 31776
rect 25832 31764 25838 31816
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 26970 31804 26976 31816
rect 26375 31776 26976 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 27157 31807 27215 31813
rect 27157 31773 27169 31807
rect 27203 31804 27215 31807
rect 27430 31804 27436 31816
rect 27203 31776 27436 31804
rect 27203 31773 27215 31776
rect 27157 31767 27215 31773
rect 27430 31764 27436 31776
rect 27488 31764 27494 31816
rect 27706 31764 27712 31816
rect 27764 31804 27770 31816
rect 28736 31813 28764 31844
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 31444 31844 32352 31872
rect 31444 31832 31450 31844
rect 28537 31807 28595 31813
rect 28537 31804 28549 31807
rect 27764 31776 28549 31804
rect 27764 31764 27770 31776
rect 28537 31773 28549 31776
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 28721 31807 28779 31813
rect 28721 31773 28733 31807
rect 28767 31773 28779 31807
rect 28721 31767 28779 31773
rect 28813 31807 28871 31813
rect 28813 31773 28825 31807
rect 28859 31804 28871 31807
rect 29086 31804 29092 31816
rect 28859 31776 29092 31804
rect 28859 31773 28871 31776
rect 28813 31767 28871 31773
rect 29086 31764 29092 31776
rect 29144 31764 29150 31816
rect 30098 31804 30104 31816
rect 30059 31776 30104 31804
rect 30098 31764 30104 31776
rect 30156 31764 30162 31816
rect 31478 31764 31484 31816
rect 31536 31764 31542 31816
rect 32324 31813 32352 31844
rect 32858 31832 32864 31884
rect 32916 31872 32922 31884
rect 35253 31875 35311 31881
rect 35253 31872 35265 31875
rect 32916 31844 35265 31872
rect 32916 31832 32922 31844
rect 35253 31841 35265 31844
rect 35299 31841 35311 31875
rect 35253 31835 35311 31841
rect 32309 31807 32367 31813
rect 32309 31773 32321 31807
rect 32355 31773 32367 31807
rect 32309 31767 32367 31773
rect 45830 31764 45836 31816
rect 45888 31804 45894 31816
rect 46584 31804 46612 31912
rect 47486 31900 47492 31912
rect 47544 31900 47550 31952
rect 46750 31872 46756 31884
rect 46711 31844 46756 31872
rect 46750 31832 46756 31844
rect 46808 31832 46814 31884
rect 47578 31872 47584 31884
rect 47539 31844 47584 31872
rect 47578 31832 47584 31844
rect 47636 31832 47642 31884
rect 45888 31776 46612 31804
rect 45888 31764 45894 31776
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 11885 31739 11943 31745
rect 11885 31705 11897 31739
rect 11931 31736 11943 31739
rect 12894 31736 12900 31748
rect 11931 31708 12900 31736
rect 11931 31705 11943 31708
rect 11885 31699 11943 31705
rect 12894 31696 12900 31708
rect 12952 31696 12958 31748
rect 15010 31736 15016 31748
rect 14971 31708 15016 31736
rect 15010 31696 15016 31708
rect 15068 31696 15074 31748
rect 22278 31736 22284 31748
rect 22239 31708 22284 31736
rect 22278 31696 22284 31708
rect 22336 31696 22342 31748
rect 23566 31736 23572 31748
rect 23506 31708 23572 31736
rect 23566 31696 23572 31708
rect 23624 31696 23630 31748
rect 30374 31736 30380 31748
rect 30335 31708 30380 31736
rect 30374 31696 30380 31708
rect 30432 31696 30438 31748
rect 34790 31696 34796 31748
rect 34848 31736 34854 31748
rect 35161 31739 35219 31745
rect 35161 31736 35173 31739
rect 34848 31708 35173 31736
rect 34848 31696 34854 31708
rect 35161 31705 35173 31708
rect 35207 31705 35219 31739
rect 46584 31736 46612 31776
rect 46845 31739 46903 31745
rect 46845 31736 46857 31739
rect 46584 31708 46857 31736
rect 35161 31699 35219 31705
rect 46845 31705 46857 31708
rect 46891 31705 46903 31739
rect 46845 31699 46903 31705
rect 18322 31668 18328 31680
rect 18283 31640 18328 31668
rect 18322 31628 18328 31640
rect 18380 31628 18386 31680
rect 25130 31668 25136 31680
rect 25091 31640 25136 31668
rect 25130 31628 25136 31640
rect 25188 31628 25194 31680
rect 25590 31668 25596 31680
rect 25551 31640 25596 31668
rect 25590 31628 25596 31640
rect 25648 31628 25654 31680
rect 28902 31628 28908 31680
rect 28960 31668 28966 31680
rect 28997 31671 29055 31677
rect 28997 31668 29009 31671
rect 28960 31640 29009 31668
rect 28960 31628 28966 31640
rect 28997 31637 29009 31640
rect 29043 31637 29055 31671
rect 34698 31668 34704 31680
rect 34659 31640 34704 31668
rect 28997 31631 29055 31637
rect 34698 31628 34704 31640
rect 34756 31628 34762 31680
rect 35069 31671 35127 31677
rect 35069 31637 35081 31671
rect 35115 31668 35127 31671
rect 35342 31668 35348 31680
rect 35115 31640 35348 31668
rect 35115 31637 35127 31640
rect 35069 31631 35127 31637
rect 35342 31628 35348 31640
rect 35400 31628 35406 31680
rect 36814 31628 36820 31680
rect 36872 31668 36878 31680
rect 43070 31668 43076 31680
rect 36872 31640 43076 31668
rect 36872 31628 36878 31640
rect 43070 31628 43076 31640
rect 43128 31628 43134 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 1636 31436 2237 31464
rect 1636 31424 1642 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 12894 31464 12900 31476
rect 12855 31436 12900 31464
rect 2225 31427 2283 31433
rect 12894 31424 12900 31436
rect 12952 31424 12958 31476
rect 14829 31467 14887 31473
rect 14829 31433 14841 31467
rect 14875 31464 14887 31467
rect 15010 31464 15016 31476
rect 14875 31436 15016 31464
rect 14875 31433 14887 31436
rect 14829 31427 14887 31433
rect 15010 31424 15016 31436
rect 15068 31424 15074 31476
rect 19061 31467 19119 31473
rect 19061 31433 19073 31467
rect 19107 31464 19119 31467
rect 19150 31464 19156 31476
rect 19107 31436 19156 31464
rect 19107 31433 19119 31436
rect 19061 31427 19119 31433
rect 19150 31424 19156 31436
rect 19208 31424 19214 31476
rect 22278 31424 22284 31476
rect 22336 31464 22342 31476
rect 22649 31467 22707 31473
rect 22649 31464 22661 31467
rect 22336 31436 22661 31464
rect 22336 31424 22342 31436
rect 22649 31433 22661 31436
rect 22695 31433 22707 31467
rect 22649 31427 22707 31433
rect 23293 31467 23351 31473
rect 23293 31433 23305 31467
rect 23339 31433 23351 31467
rect 23293 31427 23351 31433
rect 23753 31467 23811 31473
rect 23753 31433 23765 31467
rect 23799 31464 23811 31467
rect 25130 31464 25136 31476
rect 23799 31436 25136 31464
rect 23799 31433 23811 31436
rect 23753 31427 23811 31433
rect 19613 31399 19671 31405
rect 19613 31396 19625 31399
rect 18814 31368 19625 31396
rect 19613 31365 19625 31368
rect 19659 31365 19671 31399
rect 19613 31359 19671 31365
rect 2038 31288 2044 31340
rect 2096 31328 2102 31340
rect 2133 31331 2191 31337
rect 2133 31328 2145 31331
rect 2096 31300 2145 31328
rect 2096 31288 2102 31300
rect 2133 31297 2145 31300
rect 2179 31297 2191 31331
rect 2133 31291 2191 31297
rect 12805 31331 12863 31337
rect 12805 31297 12817 31331
rect 12851 31328 12863 31331
rect 14734 31328 14740 31340
rect 12851 31300 14740 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 14734 31288 14740 31300
rect 14792 31288 14798 31340
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19521 31331 19579 31337
rect 19521 31328 19533 31331
rect 19484 31300 19533 31328
rect 19484 31288 19490 31300
rect 19521 31297 19533 31300
rect 19567 31297 19579 31331
rect 19521 31291 19579 31297
rect 22833 31331 22891 31337
rect 22833 31297 22845 31331
rect 22879 31328 22891 31331
rect 23308 31328 23336 31427
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 27617 31467 27675 31473
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 27982 31464 27988 31476
rect 27663 31436 27988 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 27982 31424 27988 31436
rect 28040 31424 28046 31476
rect 28813 31467 28871 31473
rect 28813 31433 28825 31467
rect 28859 31433 28871 31467
rect 28813 31427 28871 31433
rect 29365 31467 29423 31473
rect 29365 31433 29377 31467
rect 29411 31464 29423 31467
rect 29822 31464 29828 31476
rect 29411 31436 29828 31464
rect 29411 31433 29423 31436
rect 29365 31427 29423 31433
rect 24118 31356 24124 31408
rect 24176 31396 24182 31408
rect 28828 31396 28856 31427
rect 29822 31424 29828 31436
rect 29880 31424 29886 31476
rect 30374 31424 30380 31476
rect 30432 31464 30438 31476
rect 30561 31467 30619 31473
rect 30561 31464 30573 31467
rect 30432 31436 30573 31464
rect 30432 31424 30438 31436
rect 30561 31433 30573 31436
rect 30607 31433 30619 31467
rect 30561 31427 30619 31433
rect 31386 31424 31392 31476
rect 31444 31464 31450 31476
rect 31481 31467 31539 31473
rect 31481 31464 31493 31467
rect 31444 31436 31493 31464
rect 31444 31424 31450 31436
rect 31481 31433 31493 31436
rect 31527 31433 31539 31467
rect 36814 31464 36820 31476
rect 31481 31427 31539 31433
rect 32324 31436 36820 31464
rect 24176 31368 28856 31396
rect 24176 31356 24182 31368
rect 27632 31340 27660 31368
rect 22879 31300 23336 31328
rect 23661 31331 23719 31337
rect 22879 31297 22891 31300
rect 22833 31291 22891 31297
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 24578 31328 24584 31340
rect 23707 31300 24584 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 24578 31288 24584 31300
rect 24636 31328 24642 31340
rect 24949 31331 25007 31337
rect 24949 31328 24961 31331
rect 24636 31300 24961 31328
rect 24636 31288 24642 31300
rect 24949 31297 24961 31300
rect 24995 31297 25007 31331
rect 24949 31291 25007 31297
rect 25406 31288 25412 31340
rect 25464 31328 25470 31340
rect 25777 31331 25835 31337
rect 25777 31328 25789 31331
rect 25464 31300 25789 31328
rect 25464 31288 25470 31300
rect 25777 31297 25789 31300
rect 25823 31297 25835 31331
rect 25777 31291 25835 31297
rect 26970 31288 26976 31340
rect 27028 31328 27034 31340
rect 27433 31331 27491 31337
rect 27433 31328 27445 31331
rect 27028 31300 27445 31328
rect 27028 31288 27034 31300
rect 27433 31297 27445 31300
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 27614 31288 27620 31340
rect 27672 31288 27678 31340
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31328 28687 31331
rect 28718 31328 28724 31340
rect 28675 31300 28724 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 28718 31288 28724 31300
rect 28776 31288 28782 31340
rect 29730 31328 29736 31340
rect 29691 31300 29736 31328
rect 29730 31288 29736 31300
rect 29788 31288 29794 31340
rect 30742 31328 30748 31340
rect 30703 31300 30748 31328
rect 30742 31288 30748 31300
rect 30800 31288 30806 31340
rect 31389 31331 31447 31337
rect 31389 31297 31401 31331
rect 31435 31328 31447 31331
rect 32214 31328 32220 31340
rect 31435 31300 32220 31328
rect 31435 31297 31447 31300
rect 31389 31291 31447 31297
rect 32214 31288 32220 31300
rect 32272 31288 32278 31340
rect 32324 31337 32352 31436
rect 36814 31424 36820 31436
rect 36872 31424 36878 31476
rect 35805 31399 35863 31405
rect 35805 31396 35817 31399
rect 35006 31368 35817 31396
rect 35805 31365 35817 31368
rect 35851 31365 35863 31399
rect 35805 31359 35863 31365
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31297 32367 31331
rect 35710 31328 35716 31340
rect 35671 31300 35716 31328
rect 32309 31291 32367 31297
rect 35710 31288 35716 31300
rect 35768 31288 35774 31340
rect 17313 31263 17371 31269
rect 17313 31229 17325 31263
rect 17359 31260 17371 31263
rect 17589 31263 17647 31269
rect 17359 31232 17448 31260
rect 17359 31229 17371 31232
rect 17313 31223 17371 31229
rect 17420 31124 17448 31232
rect 17589 31229 17601 31263
rect 17635 31260 17647 31263
rect 18322 31260 18328 31272
rect 17635 31232 18328 31260
rect 17635 31229 17647 31232
rect 17589 31223 17647 31229
rect 18322 31220 18328 31232
rect 18380 31220 18386 31272
rect 23937 31263 23995 31269
rect 23937 31229 23949 31263
rect 23983 31260 23995 31263
rect 24762 31260 24768 31272
rect 23983 31232 24768 31260
rect 23983 31229 23995 31232
rect 23937 31223 23995 31229
rect 24762 31220 24768 31232
rect 24820 31220 24826 31272
rect 25041 31263 25099 31269
rect 25041 31229 25053 31263
rect 25087 31229 25099 31263
rect 25041 31223 25099 31229
rect 25317 31263 25375 31269
rect 25317 31229 25329 31263
rect 25363 31260 25375 31263
rect 25590 31260 25596 31272
rect 25363 31232 25596 31260
rect 25363 31229 25375 31232
rect 25317 31223 25375 31229
rect 25056 31192 25084 31223
rect 25590 31220 25596 31232
rect 25648 31220 25654 31272
rect 29638 31220 29644 31272
rect 29696 31260 29702 31272
rect 29825 31263 29883 31269
rect 29825 31260 29837 31263
rect 29696 31232 29837 31260
rect 29696 31220 29702 31232
rect 29825 31229 29837 31232
rect 29871 31229 29883 31263
rect 29825 31223 29883 31229
rect 30009 31263 30067 31269
rect 30009 31229 30021 31263
rect 30055 31260 30067 31263
rect 32030 31260 32036 31272
rect 30055 31232 32036 31260
rect 30055 31229 30067 31232
rect 30009 31223 30067 31229
rect 32030 31220 32036 31232
rect 32088 31220 32094 31272
rect 32125 31263 32183 31269
rect 32125 31229 32137 31263
rect 32171 31229 32183 31263
rect 32125 31223 32183 31229
rect 25498 31192 25504 31204
rect 25056 31164 25504 31192
rect 25498 31152 25504 31164
rect 25556 31192 25562 31204
rect 25556 31164 25912 31192
rect 25556 31152 25562 31164
rect 18966 31124 18972 31136
rect 17420 31096 18972 31124
rect 18966 31084 18972 31096
rect 19024 31084 19030 31136
rect 25884 31133 25912 31164
rect 28074 31152 28080 31204
rect 28132 31192 28138 31204
rect 31754 31192 31760 31204
rect 28132 31164 31760 31192
rect 28132 31152 28138 31164
rect 31754 31152 31760 31164
rect 31812 31192 31818 31204
rect 32140 31192 32168 31223
rect 32398 31220 32404 31272
rect 32456 31260 32462 31272
rect 33505 31263 33563 31269
rect 33505 31260 33517 31263
rect 32456 31232 33517 31260
rect 32456 31220 32462 31232
rect 33505 31229 33517 31232
rect 33551 31229 33563 31263
rect 33505 31223 33563 31229
rect 33781 31263 33839 31269
rect 33781 31229 33793 31263
rect 33827 31260 33839 31263
rect 33870 31260 33876 31272
rect 33827 31232 33876 31260
rect 33827 31229 33839 31232
rect 33781 31223 33839 31229
rect 33870 31220 33876 31232
rect 33928 31220 33934 31272
rect 31812 31164 32168 31192
rect 31812 31152 31818 31164
rect 25869 31127 25927 31133
rect 25869 31093 25881 31127
rect 25915 31093 25927 31127
rect 25869 31087 25927 31093
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 26237 31127 26295 31133
rect 26237 31124 26249 31127
rect 26016 31096 26249 31124
rect 26016 31084 26022 31096
rect 26237 31093 26249 31096
rect 26283 31093 26295 31127
rect 26237 31087 26295 31093
rect 30650 31084 30656 31136
rect 30708 31124 30714 31136
rect 32493 31127 32551 31133
rect 32493 31124 32505 31127
rect 30708 31096 32505 31124
rect 30708 31084 30714 31096
rect 32493 31093 32505 31096
rect 32539 31093 32551 31127
rect 32493 31087 32551 31093
rect 35253 31127 35311 31133
rect 35253 31093 35265 31127
rect 35299 31124 35311 31127
rect 35342 31124 35348 31136
rect 35299 31096 35348 31124
rect 35299 31093 35311 31096
rect 35253 31087 35311 31093
rect 35342 31084 35348 31096
rect 35400 31084 35406 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 23477 30923 23535 30929
rect 23477 30889 23489 30923
rect 23523 30920 23535 30923
rect 23566 30920 23572 30932
rect 23523 30892 23572 30920
rect 23523 30889 23535 30892
rect 23477 30883 23535 30889
rect 23566 30880 23572 30892
rect 23624 30880 23630 30932
rect 26970 30920 26976 30932
rect 26931 30892 26976 30920
rect 26970 30880 26976 30892
rect 27028 30880 27034 30932
rect 29638 30920 29644 30932
rect 29599 30892 29644 30920
rect 29638 30880 29644 30892
rect 29696 30880 29702 30932
rect 31665 30923 31723 30929
rect 31665 30889 31677 30923
rect 31711 30920 31723 30923
rect 33042 30920 33048 30932
rect 31711 30892 33048 30920
rect 31711 30889 31723 30892
rect 31665 30883 31723 30889
rect 33042 30880 33048 30892
rect 33100 30880 33106 30932
rect 33870 30920 33876 30932
rect 33831 30892 33876 30920
rect 33870 30880 33876 30892
rect 33928 30880 33934 30932
rect 34701 30923 34759 30929
rect 34701 30889 34713 30923
rect 34747 30920 34759 30923
rect 34790 30920 34796 30932
rect 34747 30892 34796 30920
rect 34747 30889 34759 30892
rect 34701 30883 34759 30889
rect 34790 30880 34796 30892
rect 34848 30880 34854 30932
rect 17862 30784 17868 30796
rect 17823 30756 17868 30784
rect 17862 30744 17868 30756
rect 17920 30744 17926 30796
rect 26786 30784 26792 30796
rect 25792 30756 26792 30784
rect 12526 30716 12532 30728
rect 12487 30688 12532 30716
rect 12526 30676 12532 30688
rect 12584 30676 12590 30728
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30716 13047 30719
rect 13446 30716 13452 30728
rect 13035 30688 13452 30716
rect 13035 30685 13047 30688
rect 12989 30679 13047 30685
rect 13446 30676 13452 30688
rect 13504 30676 13510 30728
rect 14182 30676 14188 30728
rect 14240 30716 14246 30728
rect 14737 30719 14795 30725
rect 14737 30716 14749 30719
rect 14240 30688 14749 30716
rect 14240 30676 14246 30688
rect 14737 30685 14749 30688
rect 14783 30685 14795 30719
rect 16298 30716 16304 30728
rect 16259 30688 16304 30716
rect 14737 30679 14795 30685
rect 16298 30676 16304 30688
rect 16356 30676 16362 30728
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 20162 30716 20168 30728
rect 19843 30688 20168 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20162 30676 20168 30688
rect 20220 30676 20226 30728
rect 20257 30719 20315 30725
rect 20257 30685 20269 30719
rect 20303 30685 20315 30719
rect 20257 30679 20315 30685
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 24302 30716 24308 30728
rect 23431 30688 24308 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 15010 30648 15016 30660
rect 14971 30620 15016 30648
rect 15010 30608 15016 30620
rect 15068 30608 15074 30660
rect 16485 30651 16543 30657
rect 16485 30617 16497 30651
rect 16531 30648 16543 30651
rect 16574 30648 16580 30660
rect 16531 30620 16580 30648
rect 16531 30617 16543 30620
rect 16485 30611 16543 30617
rect 16574 30608 16580 30620
rect 16632 30608 16638 30660
rect 19426 30608 19432 30660
rect 19484 30648 19490 30660
rect 20272 30648 20300 30679
rect 24302 30676 24308 30688
rect 24360 30676 24366 30728
rect 25792 30725 25820 30756
rect 26786 30744 26792 30756
rect 26844 30744 26850 30796
rect 27062 30744 27068 30796
rect 27120 30784 27126 30796
rect 28074 30784 28080 30796
rect 27120 30756 28080 30784
rect 27120 30744 27126 30756
rect 25958 30725 25964 30728
rect 25777 30719 25835 30725
rect 25777 30685 25789 30719
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 25925 30719 25964 30725
rect 25925 30685 25937 30719
rect 25925 30679 25964 30685
rect 25958 30676 25964 30679
rect 26016 30676 26022 30728
rect 26142 30716 26148 30728
rect 26103 30688 26148 30716
rect 26142 30676 26148 30688
rect 26200 30676 26206 30728
rect 27172 30725 27200 30756
rect 28074 30744 28080 30756
rect 28132 30744 28138 30796
rect 29178 30744 29184 30796
rect 29236 30784 29242 30796
rect 29236 30756 29776 30784
rect 29236 30744 29242 30756
rect 26283 30719 26341 30725
rect 26283 30685 26295 30719
rect 26329 30716 26341 30719
rect 27157 30719 27215 30725
rect 26329 30688 27108 30716
rect 26329 30685 26341 30688
rect 26283 30679 26341 30685
rect 19484 30620 20300 30648
rect 19484 30608 19490 30620
rect 25222 30608 25228 30660
rect 25280 30648 25286 30660
rect 25682 30648 25688 30660
rect 25280 30620 25688 30648
rect 25280 30608 25286 30620
rect 25682 30608 25688 30620
rect 25740 30648 25746 30660
rect 26053 30651 26111 30657
rect 26053 30648 26065 30651
rect 25740 30620 26065 30648
rect 25740 30608 25746 30620
rect 26053 30617 26065 30620
rect 26099 30617 26111 30651
rect 27080 30648 27108 30688
rect 27157 30685 27169 30719
rect 27203 30685 27215 30719
rect 27157 30679 27215 30685
rect 27433 30719 27491 30725
rect 27433 30685 27445 30719
rect 27479 30716 27491 30719
rect 27522 30716 27528 30728
rect 27479 30688 27528 30716
rect 27479 30685 27491 30688
rect 27433 30679 27491 30685
rect 27522 30676 27528 30688
rect 27580 30676 27586 30728
rect 28350 30716 28356 30728
rect 28311 30688 28356 30716
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 29546 30716 29552 30728
rect 29507 30688 29552 30716
rect 29546 30676 29552 30688
rect 29604 30676 29610 30728
rect 29748 30725 29776 30756
rect 32030 30744 32036 30796
rect 32088 30784 32094 30796
rect 35345 30787 35403 30793
rect 35345 30784 35357 30787
rect 32088 30756 35357 30784
rect 32088 30744 32094 30756
rect 35345 30753 35357 30756
rect 35391 30784 35403 30787
rect 35802 30784 35808 30796
rect 35391 30756 35808 30784
rect 35391 30753 35403 30756
rect 35345 30747 35403 30753
rect 35802 30744 35808 30756
rect 35860 30744 35866 30796
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 31478 30716 31484 30728
rect 31439 30688 31484 30716
rect 29733 30679 29791 30685
rect 31478 30676 31484 30688
rect 31536 30676 31542 30728
rect 34057 30719 34115 30725
rect 34057 30685 34069 30719
rect 34103 30716 34115 30719
rect 34698 30716 34704 30728
rect 34103 30688 34704 30716
rect 34103 30685 34115 30688
rect 34057 30679 34115 30685
rect 34698 30676 34704 30688
rect 34756 30676 34762 30728
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30716 35127 30719
rect 39298 30716 39304 30728
rect 35115 30688 39304 30716
rect 35115 30685 35127 30688
rect 35069 30679 35127 30685
rect 39298 30676 39304 30688
rect 39356 30676 39362 30728
rect 27890 30648 27896 30660
rect 27080 30620 27896 30648
rect 26053 30611 26111 30617
rect 27890 30608 27896 30620
rect 27948 30648 27954 30660
rect 28442 30648 28448 30660
rect 27948 30620 28448 30648
rect 27948 30608 27954 30620
rect 28442 30608 28448 30620
rect 28500 30608 28506 30660
rect 28537 30651 28595 30657
rect 28537 30617 28549 30651
rect 28583 30648 28595 30651
rect 28994 30648 29000 30660
rect 28583 30620 29000 30648
rect 28583 30617 28595 30620
rect 28537 30611 28595 30617
rect 28994 30608 29000 30620
rect 29052 30648 29058 30660
rect 30098 30648 30104 30660
rect 29052 30620 30104 30648
rect 29052 30608 29058 30620
rect 30098 30608 30104 30620
rect 30156 30608 30162 30660
rect 32214 30608 32220 30660
rect 32272 30648 32278 30660
rect 32309 30651 32367 30657
rect 32309 30648 32321 30651
rect 32272 30620 32321 30648
rect 32272 30608 32278 30620
rect 32309 30617 32321 30620
rect 32355 30617 32367 30651
rect 32309 30611 32367 30617
rect 12345 30583 12403 30589
rect 12345 30549 12357 30583
rect 12391 30580 12403 30583
rect 12434 30580 12440 30592
rect 12391 30552 12440 30580
rect 12391 30549 12403 30552
rect 12345 30543 12403 30549
rect 12434 30540 12440 30552
rect 12492 30540 12498 30592
rect 13078 30580 13084 30592
rect 13039 30552 13084 30580
rect 13078 30540 13084 30552
rect 13136 30540 13142 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 19392 30552 19625 30580
rect 19392 30540 19398 30552
rect 19613 30549 19625 30552
rect 19659 30549 19671 30583
rect 20346 30580 20352 30592
rect 20307 30552 20352 30580
rect 19613 30543 19671 30549
rect 20346 30540 20352 30552
rect 20404 30540 20410 30592
rect 24854 30540 24860 30592
rect 24912 30580 24918 30592
rect 26421 30583 26479 30589
rect 26421 30580 26433 30583
rect 24912 30552 26433 30580
rect 24912 30540 24918 30552
rect 26421 30549 26433 30552
rect 26467 30549 26479 30583
rect 27338 30580 27344 30592
rect 27299 30552 27344 30580
rect 26421 30543 26479 30549
rect 27338 30540 27344 30552
rect 27396 30540 27402 30592
rect 31754 30540 31760 30592
rect 31812 30580 31818 30592
rect 32401 30583 32459 30589
rect 32401 30580 32413 30583
rect 31812 30552 32413 30580
rect 31812 30540 31818 30552
rect 32401 30549 32413 30552
rect 32447 30549 32459 30583
rect 32401 30543 32459 30549
rect 35158 30540 35164 30592
rect 35216 30580 35222 30592
rect 35216 30552 35261 30580
rect 35216 30540 35222 30552
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 13909 30379 13967 30385
rect 13909 30345 13921 30379
rect 13955 30376 13967 30379
rect 14366 30376 14372 30388
rect 13955 30348 14372 30376
rect 13955 30345 13967 30348
rect 13909 30339 13967 30345
rect 14366 30336 14372 30348
rect 14424 30376 14430 30388
rect 16298 30376 16304 30388
rect 14424 30348 16304 30376
rect 14424 30336 14430 30348
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 25133 30379 25191 30385
rect 24044 30348 24992 30376
rect 12434 30308 12440 30320
rect 12395 30280 12440 30308
rect 12434 30268 12440 30280
rect 12492 30268 12498 30320
rect 13078 30268 13084 30320
rect 13136 30268 13142 30320
rect 14090 30268 14096 30320
rect 14148 30308 14154 30320
rect 14734 30308 14740 30320
rect 14148 30280 14740 30308
rect 14148 30268 14154 30280
rect 14734 30268 14740 30280
rect 14792 30308 14798 30320
rect 19245 30311 19303 30317
rect 14792 30280 15700 30308
rect 14792 30268 14798 30280
rect 9766 30240 9772 30252
rect 9727 30212 9772 30240
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30209 10287 30243
rect 10229 30203 10287 30209
rect 9214 30132 9220 30184
rect 9272 30172 9278 30184
rect 10244 30172 10272 30203
rect 14274 30200 14280 30252
rect 14332 30240 14338 30252
rect 15672 30249 15700 30280
rect 19245 30277 19257 30311
rect 19291 30308 19303 30311
rect 19334 30308 19340 30320
rect 19291 30280 19340 30308
rect 19291 30277 19303 30280
rect 19245 30271 19303 30277
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 24044 30308 24072 30348
rect 22296 30280 24072 30308
rect 14829 30243 14887 30249
rect 14829 30240 14841 30243
rect 14332 30212 14841 30240
rect 14332 30200 14338 30212
rect 14829 30209 14841 30212
rect 14875 30240 14887 30243
rect 15657 30243 15715 30249
rect 14875 30212 15056 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 9272 30144 10272 30172
rect 12161 30175 12219 30181
rect 9272 30132 9278 30144
rect 12161 30141 12173 30175
rect 12207 30141 12219 30175
rect 12161 30135 12219 30141
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30141 14979 30175
rect 15028 30172 15056 30212
rect 15657 30209 15669 30243
rect 15703 30209 15715 30243
rect 15657 30203 15715 30209
rect 20346 30200 20352 30252
rect 20404 30200 20410 30252
rect 22296 30249 22324 30280
rect 24394 30268 24400 30320
rect 24452 30268 24458 30320
rect 24964 30308 24992 30348
rect 25133 30345 25145 30379
rect 25179 30376 25191 30379
rect 26142 30376 26148 30388
rect 25179 30348 26148 30376
rect 25179 30345 25191 30348
rect 25133 30339 25191 30345
rect 26142 30336 26148 30348
rect 26200 30336 26206 30388
rect 26970 30336 26976 30388
rect 27028 30376 27034 30388
rect 27522 30376 27528 30388
rect 27028 30348 27528 30376
rect 27028 30336 27034 30348
rect 27522 30336 27528 30348
rect 27580 30376 27586 30388
rect 34701 30379 34759 30385
rect 27580 30348 28396 30376
rect 27580 30336 27586 30348
rect 27338 30308 27344 30320
rect 24964 30280 27344 30308
rect 27338 30268 27344 30280
rect 27396 30308 27402 30320
rect 27433 30311 27491 30317
rect 27433 30308 27445 30311
rect 27396 30280 27445 30308
rect 27396 30268 27402 30280
rect 27433 30277 27445 30280
rect 27479 30277 27491 30311
rect 27433 30271 27491 30277
rect 27617 30311 27675 30317
rect 27617 30277 27629 30311
rect 27663 30308 27675 30311
rect 27798 30308 27804 30320
rect 27663 30280 27804 30308
rect 27663 30277 27675 30280
rect 27617 30271 27675 30277
rect 27798 30268 27804 30280
rect 27856 30308 27862 30320
rect 28261 30311 28319 30317
rect 28261 30308 28273 30311
rect 27856 30280 28273 30308
rect 27856 30268 27862 30280
rect 28261 30277 28273 30280
rect 28307 30277 28319 30311
rect 28261 30271 28319 30277
rect 22281 30243 22339 30249
rect 22281 30209 22293 30243
rect 22327 30209 22339 30243
rect 28074 30240 28080 30252
rect 28035 30212 28080 30240
rect 22281 30203 22339 30209
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 28368 30249 28396 30348
rect 34701 30345 34713 30379
rect 34747 30376 34759 30379
rect 35158 30376 35164 30388
rect 34747 30348 35164 30376
rect 34747 30345 34759 30348
rect 34701 30339 34759 30345
rect 35158 30336 35164 30348
rect 35216 30336 35222 30388
rect 28442 30268 28448 30320
rect 28500 30308 28506 30320
rect 29365 30311 29423 30317
rect 29365 30308 29377 30311
rect 28500 30280 29377 30308
rect 28500 30268 28506 30280
rect 29365 30277 29377 30280
rect 29411 30277 29423 30311
rect 29365 30271 29423 30277
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28353 30203 28411 30209
rect 29181 30243 29239 30249
rect 29181 30209 29193 30243
rect 29227 30209 29239 30243
rect 34514 30240 34520 30252
rect 34475 30212 34520 30240
rect 29181 30203 29239 30209
rect 16666 30172 16672 30184
rect 15028 30144 16672 30172
rect 14921 30135 14979 30141
rect 9585 30039 9643 30045
rect 9585 30005 9597 30039
rect 9631 30036 9643 30039
rect 9674 30036 9680 30048
rect 9631 30008 9680 30036
rect 9631 30005 9643 30008
rect 9585 29999 9643 30005
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 10318 30036 10324 30048
rect 10279 30008 10324 30036
rect 10318 29996 10324 30008
rect 10376 29996 10382 30048
rect 12176 30036 12204 30135
rect 14936 30104 14964 30135
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 16853 30175 16911 30181
rect 16853 30141 16865 30175
rect 16899 30172 16911 30175
rect 17494 30172 17500 30184
rect 16899 30144 17500 30172
rect 16899 30141 16911 30144
rect 16853 30135 16911 30141
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 17589 30175 17647 30181
rect 17589 30141 17601 30175
rect 17635 30141 17647 30175
rect 18966 30172 18972 30184
rect 18927 30144 18972 30172
rect 17589 30135 17647 30141
rect 15470 30104 15476 30116
rect 14936 30076 15476 30104
rect 15470 30064 15476 30076
rect 15528 30064 15534 30116
rect 12618 30036 12624 30048
rect 12176 30008 12624 30036
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 15197 30039 15255 30045
rect 15197 30005 15209 30039
rect 15243 30036 15255 30039
rect 15378 30036 15384 30048
rect 15243 30008 15384 30036
rect 15243 30005 15255 30008
rect 15197 29999 15255 30005
rect 15378 29996 15384 30008
rect 15436 29996 15442 30048
rect 15746 30036 15752 30048
rect 15707 30008 15752 30036
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 15838 29996 15844 30048
rect 15896 30036 15902 30048
rect 17604 30036 17632 30135
rect 18966 30132 18972 30144
rect 19024 30132 19030 30184
rect 22094 30132 22100 30184
rect 22152 30172 22158 30184
rect 22646 30172 22652 30184
rect 22152 30144 22652 30172
rect 22152 30132 22158 30144
rect 22646 30132 22652 30144
rect 22704 30172 22710 30184
rect 23385 30175 23443 30181
rect 23385 30172 23397 30175
rect 22704 30144 23397 30172
rect 22704 30132 22710 30144
rect 23385 30141 23397 30144
rect 23431 30141 23443 30175
rect 23385 30135 23443 30141
rect 23661 30175 23719 30181
rect 23661 30141 23673 30175
rect 23707 30172 23719 30175
rect 24854 30172 24860 30184
rect 23707 30144 24860 30172
rect 23707 30141 23719 30144
rect 23661 30135 23719 30141
rect 24854 30132 24860 30144
rect 24912 30132 24918 30184
rect 29196 30172 29224 30203
rect 34514 30200 34520 30212
rect 34572 30200 34578 30252
rect 34606 30200 34612 30252
rect 34664 30240 34670 30252
rect 34701 30243 34759 30249
rect 34701 30240 34713 30243
rect 34664 30212 34713 30240
rect 34664 30200 34670 30212
rect 34701 30209 34713 30212
rect 34747 30240 34759 30243
rect 34790 30240 34796 30252
rect 34747 30212 34796 30240
rect 34747 30209 34759 30212
rect 34701 30203 34759 30209
rect 34790 30200 34796 30212
rect 34848 30200 34854 30252
rect 30006 30172 30012 30184
rect 28092 30144 30012 30172
rect 28092 30113 28120 30144
rect 30006 30132 30012 30144
rect 30064 30132 30070 30184
rect 28077 30107 28135 30113
rect 28077 30073 28089 30107
rect 28123 30073 28135 30107
rect 28077 30067 28135 30073
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 32490 30104 32496 30116
rect 28408 30076 32496 30104
rect 28408 30064 28414 30076
rect 32490 30064 32496 30076
rect 32548 30064 32554 30116
rect 15896 30008 17632 30036
rect 20717 30039 20775 30045
rect 15896 29996 15902 30008
rect 20717 30005 20729 30039
rect 20763 30036 20775 30039
rect 20898 30036 20904 30048
rect 20763 30008 20904 30036
rect 20763 30005 20775 30008
rect 20717 29999 20775 30005
rect 20898 29996 20904 30008
rect 20956 29996 20962 30048
rect 22278 29996 22284 30048
rect 22336 30036 22342 30048
rect 22373 30039 22431 30045
rect 22373 30036 22385 30039
rect 22336 30008 22385 30036
rect 22336 29996 22342 30008
rect 22373 30005 22385 30008
rect 22419 30005 22431 30039
rect 22373 29999 22431 30005
rect 25682 29996 25688 30048
rect 25740 30036 25746 30048
rect 28534 30036 28540 30048
rect 25740 30008 28540 30036
rect 25740 29996 25746 30008
rect 28534 29996 28540 30008
rect 28592 29996 28598 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 12989 29835 13047 29841
rect 12989 29832 13001 29835
rect 12124 29804 13001 29832
rect 12124 29792 12130 29804
rect 12989 29801 13001 29804
rect 13035 29801 13047 29835
rect 12989 29795 13047 29801
rect 16666 29792 16672 29844
rect 16724 29832 16730 29844
rect 16853 29835 16911 29841
rect 16853 29832 16865 29835
rect 16724 29804 16865 29832
rect 16724 29792 16730 29804
rect 16853 29801 16865 29804
rect 16899 29801 16911 29835
rect 17494 29832 17500 29844
rect 17455 29804 17500 29832
rect 16853 29795 16911 29801
rect 17494 29792 17500 29804
rect 17552 29792 17558 29844
rect 20162 29792 20168 29844
rect 20220 29832 20226 29844
rect 20441 29835 20499 29841
rect 20441 29832 20453 29835
rect 20220 29804 20453 29832
rect 20220 29792 20226 29804
rect 20441 29801 20453 29804
rect 20487 29801 20499 29835
rect 20441 29795 20499 29801
rect 20806 29792 20812 29844
rect 20864 29832 20870 29844
rect 21818 29832 21824 29844
rect 20864 29804 21824 29832
rect 20864 29792 20870 29804
rect 21818 29792 21824 29804
rect 21876 29832 21882 29844
rect 21876 29804 23428 29832
rect 21876 29792 21882 29804
rect 11882 29724 11888 29776
rect 11940 29764 11946 29776
rect 14185 29767 14243 29773
rect 14185 29764 14197 29767
rect 11940 29736 14197 29764
rect 11940 29724 11946 29736
rect 14185 29733 14197 29736
rect 14231 29733 14243 29767
rect 14185 29727 14243 29733
rect 9674 29696 9680 29708
rect 9635 29668 9680 29696
rect 9674 29656 9680 29668
rect 9732 29656 9738 29708
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11698 29696 11704 29708
rect 11195 29668 11704 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11698 29656 11704 29668
rect 11756 29696 11762 29708
rect 12069 29699 12127 29705
rect 12069 29696 12081 29699
rect 11756 29668 12081 29696
rect 11756 29656 11762 29668
rect 12069 29665 12081 29668
rect 12115 29665 12127 29699
rect 12069 29659 12127 29665
rect 12544 29668 13492 29696
rect 9306 29588 9312 29640
rect 9364 29628 9370 29640
rect 9401 29631 9459 29637
rect 9401 29628 9413 29631
rect 9364 29600 9413 29628
rect 9364 29588 9370 29600
rect 9401 29597 9413 29600
rect 9447 29597 9459 29631
rect 12158 29628 12164 29640
rect 12119 29600 12164 29628
rect 9401 29591 9459 29597
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 12544 29637 12572 29668
rect 13464 29637 13492 29668
rect 15010 29656 15016 29708
rect 15068 29696 15074 29708
rect 15105 29699 15163 29705
rect 15105 29696 15117 29699
rect 15068 29668 15117 29696
rect 15068 29656 15074 29668
rect 15105 29665 15117 29668
rect 15151 29665 15163 29699
rect 15378 29696 15384 29708
rect 15339 29668 15384 29696
rect 15105 29659 15163 29665
rect 15378 29656 15384 29668
rect 15436 29656 15442 29708
rect 20806 29696 20812 29708
rect 19260 29668 20812 29696
rect 19260 29640 19288 29668
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 21082 29696 21088 29708
rect 21043 29668 21088 29696
rect 21082 29656 21088 29668
rect 21140 29696 21146 29708
rect 21726 29696 21732 29708
rect 21140 29668 21732 29696
rect 21140 29656 21146 29668
rect 21726 29656 21732 29668
rect 21784 29656 21790 29708
rect 21821 29699 21879 29705
rect 21821 29665 21833 29699
rect 21867 29696 21879 29699
rect 22741 29699 22799 29705
rect 22741 29696 22753 29699
rect 21867 29668 22753 29696
rect 21867 29665 21879 29668
rect 21821 29659 21879 29665
rect 22741 29665 22753 29668
rect 22787 29665 22799 29699
rect 22741 29659 22799 29665
rect 12529 29631 12587 29637
rect 12529 29597 12541 29631
rect 12575 29597 12587 29631
rect 13219 29631 13277 29637
rect 13219 29628 13231 29631
rect 12529 29591 12587 29597
rect 13207 29597 13231 29628
rect 13265 29597 13277 29631
rect 13207 29591 13277 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29628 13507 29631
rect 14274 29628 14280 29640
rect 13495 29600 14136 29628
rect 14235 29600 14280 29628
rect 13495 29597 13507 29600
rect 13449 29591 13507 29597
rect 10318 29520 10324 29572
rect 10376 29520 10382 29572
rect 12986 29560 12992 29572
rect 12360 29532 12992 29560
rect 11238 29452 11244 29504
rect 11296 29492 11302 29504
rect 12360 29501 12388 29532
rect 12986 29520 12992 29532
rect 13044 29560 13050 29572
rect 13207 29560 13235 29591
rect 14108 29569 14136 29600
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14366 29588 14372 29640
rect 14424 29628 14430 29640
rect 17405 29631 17463 29637
rect 14424 29600 14469 29628
rect 14424 29588 14430 29600
rect 17405 29597 17417 29631
rect 17451 29628 17463 29631
rect 18414 29628 18420 29640
rect 17451 29600 18420 29628
rect 17451 29597 17463 29600
rect 17405 29591 17463 29597
rect 18414 29588 18420 29600
rect 18472 29588 18478 29640
rect 19242 29628 19248 29640
rect 19155 29600 19248 29628
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 20714 29588 20720 29640
rect 20772 29628 20778 29640
rect 21913 29631 21971 29637
rect 21913 29628 21925 29631
rect 20772 29600 21925 29628
rect 20772 29588 20778 29600
rect 21913 29597 21925 29600
rect 21959 29597 21971 29631
rect 21913 29591 21971 29597
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29597 22063 29631
rect 22005 29591 22063 29597
rect 13357 29563 13415 29569
rect 13357 29560 13369 29563
rect 13044 29532 13235 29560
rect 13280 29532 13369 29560
rect 13044 29520 13050 29532
rect 11885 29495 11943 29501
rect 11885 29492 11897 29495
rect 11296 29464 11897 29492
rect 11296 29452 11302 29464
rect 11885 29461 11897 29464
rect 11931 29461 11943 29495
rect 11885 29455 11943 29461
rect 12345 29495 12403 29501
rect 12345 29461 12357 29495
rect 12391 29461 12403 29495
rect 12345 29455 12403 29461
rect 12437 29495 12495 29501
rect 12437 29461 12449 29495
rect 12483 29492 12495 29495
rect 13078 29492 13084 29504
rect 12483 29464 13084 29492
rect 12483 29461 12495 29464
rect 12437 29455 12495 29461
rect 13078 29452 13084 29464
rect 13136 29492 13142 29504
rect 13280 29492 13308 29532
rect 13357 29529 13369 29532
rect 13403 29529 13415 29563
rect 13357 29523 13415 29529
rect 14093 29563 14151 29569
rect 14093 29529 14105 29563
rect 14139 29560 14151 29563
rect 15470 29560 15476 29572
rect 14139 29532 15476 29560
rect 14139 29529 14151 29532
rect 14093 29523 14151 29529
rect 15470 29520 15476 29532
rect 15528 29520 15534 29572
rect 16758 29560 16764 29572
rect 16606 29532 16764 29560
rect 16758 29520 16764 29532
rect 16816 29520 16822 29572
rect 21082 29520 21088 29572
rect 21140 29560 21146 29572
rect 22020 29560 22048 29591
rect 22094 29588 22100 29640
rect 22152 29628 22158 29640
rect 22152 29600 22197 29628
rect 22152 29588 22158 29600
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 23400 29637 23428 29804
rect 24394 29792 24400 29844
rect 24452 29832 24458 29844
rect 24489 29835 24547 29841
rect 24489 29832 24501 29835
rect 24452 29804 24501 29832
rect 24452 29792 24458 29804
rect 24489 29801 24501 29804
rect 24535 29801 24547 29835
rect 24489 29795 24547 29801
rect 25961 29835 26019 29841
rect 25961 29801 25973 29835
rect 26007 29832 26019 29835
rect 26050 29832 26056 29844
rect 26007 29804 26056 29832
rect 26007 29801 26019 29804
rect 25961 29795 26019 29801
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 27062 29832 27068 29844
rect 27023 29804 27068 29832
rect 27062 29792 27068 29804
rect 27120 29792 27126 29844
rect 27982 29792 27988 29844
rect 28040 29832 28046 29844
rect 28350 29832 28356 29844
rect 28040 29804 28356 29832
rect 28040 29792 28046 29804
rect 28350 29792 28356 29804
rect 28408 29792 28414 29844
rect 28534 29832 28540 29844
rect 28495 29804 28540 29832
rect 28534 29792 28540 29804
rect 28592 29792 28598 29844
rect 29914 29792 29920 29844
rect 29972 29832 29978 29844
rect 30193 29835 30251 29841
rect 30193 29832 30205 29835
rect 29972 29804 30205 29832
rect 29972 29792 29978 29804
rect 30193 29801 30205 29804
rect 30239 29801 30251 29835
rect 30926 29832 30932 29844
rect 30887 29804 30932 29832
rect 30193 29795 30251 29801
rect 30926 29792 30932 29804
rect 30984 29792 30990 29844
rect 46842 29832 46848 29844
rect 31726 29804 46848 29832
rect 26510 29724 26516 29776
rect 26568 29724 26574 29776
rect 26878 29724 26884 29776
rect 26936 29764 26942 29776
rect 31726 29764 31754 29804
rect 46842 29792 46848 29804
rect 46900 29792 46906 29844
rect 26936 29736 31754 29764
rect 26936 29724 26942 29736
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 22336 29600 22661 29628
rect 22336 29588 22342 29600
rect 22649 29597 22661 29600
rect 22695 29597 22707 29631
rect 22649 29591 22707 29597
rect 22833 29631 22891 29637
rect 22833 29597 22845 29631
rect 22879 29597 22891 29631
rect 22833 29591 22891 29597
rect 23385 29631 23443 29637
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 22848 29560 22876 29591
rect 24302 29588 24308 29640
rect 24360 29628 24366 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 24360 29600 24409 29628
rect 24360 29588 24366 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 26142 29588 26148 29640
rect 26200 29637 26206 29640
rect 26200 29631 26249 29637
rect 26200 29597 26203 29631
rect 26237 29597 26249 29631
rect 26323 29628 26329 29640
rect 26284 29600 26329 29628
rect 26200 29591 26249 29597
rect 26200 29588 26206 29591
rect 26323 29588 26329 29600
rect 26381 29588 26387 29640
rect 26426 29631 26484 29637
rect 26426 29597 26438 29631
rect 26472 29628 26484 29631
rect 26528 29628 26556 29724
rect 27798 29696 27804 29708
rect 26620 29668 27804 29696
rect 26620 29637 26648 29668
rect 27798 29656 27804 29668
rect 27856 29656 27862 29708
rect 30650 29696 30656 29708
rect 29564 29668 30656 29696
rect 26472 29600 26556 29628
rect 26605 29631 26663 29637
rect 26472 29597 26484 29600
rect 26426 29591 26484 29597
rect 26605 29597 26617 29631
rect 26651 29597 26663 29631
rect 26605 29591 26663 29597
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 27249 29631 27307 29637
rect 27249 29597 27261 29631
rect 27295 29628 27307 29631
rect 28718 29628 28724 29640
rect 27295 29600 28724 29628
rect 27295 29597 27307 29600
rect 27249 29591 27307 29597
rect 21140 29532 22048 29560
rect 22480 29532 22876 29560
rect 27080 29560 27108 29591
rect 28718 29588 28724 29600
rect 28776 29588 28782 29640
rect 29564 29637 29592 29668
rect 30650 29656 30656 29668
rect 30708 29656 30714 29708
rect 32858 29656 32864 29708
rect 32916 29696 32922 29708
rect 33229 29699 33287 29705
rect 33229 29696 33241 29699
rect 32916 29668 33241 29696
rect 32916 29656 32922 29668
rect 33229 29665 33241 29668
rect 33275 29665 33287 29699
rect 33229 29659 33287 29665
rect 29730 29637 29736 29640
rect 29549 29631 29607 29637
rect 29549 29597 29561 29631
rect 29595 29597 29607 29631
rect 29549 29591 29607 29597
rect 29697 29631 29736 29637
rect 29697 29597 29709 29631
rect 29697 29591 29736 29597
rect 29730 29588 29736 29591
rect 29788 29588 29794 29640
rect 30006 29628 30012 29640
rect 30064 29637 30070 29640
rect 29972 29600 30012 29628
rect 30006 29588 30012 29600
rect 30064 29591 30072 29637
rect 30190 29628 30196 29640
rect 30116 29600 30196 29628
rect 30064 29588 30070 29591
rect 28258 29560 28264 29572
rect 27080 29532 28264 29560
rect 21140 29520 21146 29532
rect 13136 29464 13308 29492
rect 13136 29452 13142 29464
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19392 29464 19441 29492
rect 19392 29452 19398 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 20165 29495 20223 29501
rect 20165 29461 20177 29495
rect 20211 29492 20223 29495
rect 20714 29492 20720 29504
rect 20211 29464 20720 29492
rect 20211 29461 20223 29464
rect 20165 29455 20223 29461
rect 20714 29452 20720 29464
rect 20772 29492 20778 29504
rect 20809 29495 20867 29501
rect 20809 29492 20821 29495
rect 20772 29464 20821 29492
rect 20772 29452 20778 29464
rect 20809 29461 20821 29464
rect 20855 29461 20867 29495
rect 20809 29455 20867 29461
rect 20901 29495 20959 29501
rect 20901 29461 20913 29495
rect 20947 29492 20959 29495
rect 21637 29495 21695 29501
rect 21637 29492 21649 29495
rect 20947 29464 21649 29492
rect 20947 29461 20959 29464
rect 20901 29455 20959 29461
rect 21637 29461 21649 29464
rect 21683 29461 21695 29495
rect 21637 29455 21695 29461
rect 22002 29452 22008 29504
rect 22060 29492 22066 29504
rect 22480 29492 22508 29532
rect 28258 29520 28264 29532
rect 28316 29520 28322 29572
rect 28442 29560 28448 29572
rect 28403 29532 28448 29560
rect 28442 29520 28448 29532
rect 28500 29520 28506 29572
rect 28534 29520 28540 29572
rect 28592 29560 28598 29572
rect 29825 29563 29883 29569
rect 29825 29560 29837 29563
rect 28592 29532 29837 29560
rect 28592 29520 28598 29532
rect 29825 29529 29837 29532
rect 29871 29529 29883 29563
rect 29825 29523 29883 29529
rect 29917 29563 29975 29569
rect 29917 29529 29929 29563
rect 29963 29560 29975 29563
rect 30116 29560 30144 29600
rect 30190 29588 30196 29600
rect 30248 29588 30254 29640
rect 30745 29631 30803 29637
rect 30745 29597 30757 29631
rect 30791 29628 30803 29631
rect 31478 29628 31484 29640
rect 30791 29600 31484 29628
rect 30791 29597 30803 29600
rect 30745 29591 30803 29597
rect 29963 29532 30144 29560
rect 29963 29529 29975 29532
rect 29917 29523 29975 29529
rect 22060 29464 22508 29492
rect 23477 29495 23535 29501
rect 22060 29452 22066 29464
rect 23477 29461 23489 29495
rect 23523 29492 23535 29495
rect 24394 29492 24400 29504
rect 23523 29464 24400 29492
rect 23523 29461 23535 29464
rect 23477 29455 23535 29461
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 26234 29452 26240 29504
rect 26292 29492 26298 29504
rect 27433 29495 27491 29501
rect 27433 29492 27445 29495
rect 26292 29464 27445 29492
rect 26292 29452 26298 29464
rect 27433 29461 27445 29464
rect 27479 29461 27491 29495
rect 27433 29455 27491 29461
rect 27522 29452 27528 29504
rect 27580 29492 27586 29504
rect 30760 29492 30788 29591
rect 31478 29588 31484 29600
rect 31536 29588 31542 29640
rect 48130 29628 48136 29640
rect 48091 29600 48136 29628
rect 48130 29588 48136 29600
rect 48188 29588 48194 29640
rect 32858 29520 32864 29572
rect 32916 29560 32922 29572
rect 33137 29563 33195 29569
rect 33137 29560 33149 29563
rect 32916 29532 33149 29560
rect 32916 29520 32922 29532
rect 33137 29529 33149 29532
rect 33183 29529 33195 29563
rect 33137 29523 33195 29529
rect 27580 29464 30788 29492
rect 32677 29495 32735 29501
rect 27580 29452 27586 29464
rect 32677 29461 32689 29495
rect 32723 29492 32735 29495
rect 32766 29492 32772 29504
rect 32723 29464 32772 29492
rect 32723 29461 32735 29464
rect 32677 29455 32735 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 33045 29495 33103 29501
rect 33045 29461 33057 29495
rect 33091 29492 33103 29495
rect 34054 29492 34060 29504
rect 33091 29464 34060 29492
rect 33091 29461 33103 29464
rect 33045 29455 33103 29461
rect 34054 29452 34060 29464
rect 34112 29452 34118 29504
rect 47394 29452 47400 29504
rect 47452 29492 47458 29504
rect 47949 29495 48007 29501
rect 47949 29492 47961 29495
rect 47452 29464 47961 29492
rect 47452 29452 47458 29464
rect 47949 29461 47961 29464
rect 47995 29461 48007 29495
rect 47949 29455 48007 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 9306 29288 9312 29300
rect 9267 29260 9312 29288
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 10505 29291 10563 29297
rect 10505 29288 10517 29291
rect 9824 29260 10517 29288
rect 9824 29248 9830 29260
rect 10505 29257 10517 29260
rect 10551 29257 10563 29291
rect 10505 29251 10563 29257
rect 12253 29291 12311 29297
rect 12253 29257 12265 29291
rect 12299 29288 12311 29291
rect 12434 29288 12440 29300
rect 12299 29260 12440 29288
rect 12299 29257 12311 29260
rect 12253 29251 12311 29257
rect 12434 29248 12440 29260
rect 12492 29248 12498 29300
rect 13078 29288 13084 29300
rect 12991 29260 13084 29288
rect 13078 29248 13084 29260
rect 13136 29288 13142 29300
rect 14274 29288 14280 29300
rect 13136 29260 14280 29288
rect 13136 29248 13142 29260
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 14366 29248 14372 29300
rect 14424 29248 14430 29300
rect 16574 29248 16580 29300
rect 16632 29288 16638 29300
rect 16761 29291 16819 29297
rect 16761 29288 16773 29291
rect 16632 29260 16773 29288
rect 16632 29248 16638 29260
rect 16761 29257 16773 29260
rect 16807 29257 16819 29291
rect 21821 29291 21879 29297
rect 16761 29251 16819 29257
rect 20732 29260 21220 29288
rect 11698 29180 11704 29232
rect 11756 29220 11762 29232
rect 12713 29223 12771 29229
rect 12713 29220 12725 29223
rect 11756 29192 12725 29220
rect 11756 29180 11762 29192
rect 12713 29189 12725 29192
rect 12759 29189 12771 29223
rect 12986 29220 12992 29232
rect 12899 29192 12992 29220
rect 12713 29183 12771 29189
rect 12986 29180 12992 29192
rect 13044 29220 13050 29232
rect 14384 29220 14412 29248
rect 13044 29192 14412 29220
rect 14461 29223 14519 29229
rect 13044 29180 13050 29192
rect 14461 29189 14473 29223
rect 14507 29220 14519 29223
rect 15746 29220 15752 29232
rect 14507 29192 15752 29220
rect 14507 29189 14519 29192
rect 14461 29183 14519 29189
rect 15746 29180 15752 29192
rect 15804 29180 15810 29232
rect 16117 29223 16175 29229
rect 16117 29189 16129 29223
rect 16163 29220 16175 29223
rect 20732 29220 20760 29260
rect 20898 29220 20904 29232
rect 16163 29192 20760 29220
rect 20859 29192 20904 29220
rect 16163 29189 16175 29192
rect 16117 29183 16175 29189
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 21082 29220 21088 29232
rect 21043 29192 21088 29220
rect 21082 29180 21088 29192
rect 21140 29180 21146 29232
rect 21192 29220 21220 29260
rect 21821 29257 21833 29291
rect 21867 29288 21879 29291
rect 22094 29288 22100 29300
rect 21867 29260 22100 29288
rect 21867 29257 21879 29260
rect 21821 29251 21879 29257
rect 22094 29248 22100 29260
rect 22152 29248 22158 29300
rect 22925 29291 22983 29297
rect 22925 29257 22937 29291
rect 22971 29288 22983 29291
rect 22971 29260 27016 29288
rect 22971 29257 22983 29260
rect 22925 29251 22983 29257
rect 26878 29220 26884 29232
rect 21192 29192 26884 29220
rect 26878 29180 26884 29192
rect 26936 29180 26942 29232
rect 26988 29220 27016 29260
rect 28994 29248 29000 29300
rect 29052 29288 29058 29300
rect 32398 29288 32404 29300
rect 29052 29260 32404 29288
rect 29052 29248 29058 29260
rect 26988 29192 27384 29220
rect 8478 29112 8484 29164
rect 8536 29152 8542 29164
rect 9217 29155 9275 29161
rect 9217 29152 9229 29155
rect 8536 29124 9229 29152
rect 8536 29112 8542 29124
rect 9217 29121 9229 29124
rect 9263 29121 9275 29155
rect 11882 29152 11888 29164
rect 11843 29124 11888 29152
rect 9217 29115 9275 29121
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 12066 29152 12072 29164
rect 12027 29124 12072 29152
rect 12066 29112 12072 29124
rect 12124 29112 12130 29164
rect 12897 29155 12955 29161
rect 12897 29121 12909 29155
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 9950 29044 9956 29096
rect 10008 29084 10014 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 10008 29056 10057 29084
rect 10008 29044 10014 29056
rect 10045 29053 10057 29056
rect 10091 29053 10103 29087
rect 10045 29047 10103 29053
rect 12158 29044 12164 29096
rect 12216 29084 12222 29096
rect 12912 29084 12940 29115
rect 16022 29112 16028 29164
rect 16080 29152 16086 29164
rect 16669 29155 16727 29161
rect 16669 29152 16681 29155
rect 16080 29124 16681 29152
rect 16080 29112 16086 29124
rect 16669 29121 16681 29124
rect 16715 29121 16727 29155
rect 19058 29152 19064 29164
rect 19019 29124 19064 29152
rect 16669 29115 16727 29121
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 20916 29152 20944 29180
rect 27356 29164 27384 29192
rect 22002 29152 22008 29164
rect 20916 29124 22008 29152
rect 22002 29112 22008 29124
rect 22060 29112 22066 29164
rect 22738 29152 22744 29164
rect 22699 29124 22744 29152
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 26970 29152 26976 29164
rect 22848 29124 26976 29152
rect 12216 29056 12940 29084
rect 12216 29044 12222 29056
rect 13354 29044 13360 29096
rect 13412 29084 13418 29096
rect 14277 29087 14335 29093
rect 14277 29084 14289 29087
rect 13412 29056 14289 29084
rect 13412 29044 13418 29056
rect 14277 29053 14289 29056
rect 14323 29053 14335 29087
rect 22278 29084 22284 29096
rect 22239 29056 22284 29084
rect 14277 29047 14335 29053
rect 22278 29044 22284 29056
rect 22336 29044 22342 29096
rect 22370 29044 22376 29096
rect 22428 29084 22434 29096
rect 22848 29084 22876 29124
rect 26970 29112 26976 29124
rect 27028 29112 27034 29164
rect 27065 29155 27123 29161
rect 27065 29121 27077 29155
rect 27111 29121 27123 29155
rect 27338 29152 27344 29164
rect 27299 29124 27344 29152
rect 27065 29115 27123 29121
rect 27080 29084 27108 29115
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 27798 29152 27804 29164
rect 27759 29124 27804 29152
rect 27798 29112 27804 29124
rect 27856 29112 27862 29164
rect 27982 29112 27988 29164
rect 28040 29152 28046 29164
rect 28077 29155 28135 29161
rect 28077 29152 28089 29155
rect 28040 29124 28089 29152
rect 28040 29112 28046 29124
rect 28077 29121 28089 29124
rect 28123 29121 28135 29155
rect 28718 29152 28724 29164
rect 28077 29115 28135 29121
rect 28460 29124 28724 29152
rect 28460 29093 28488 29124
rect 28718 29112 28724 29124
rect 28776 29112 28782 29164
rect 29089 29155 29147 29161
rect 29089 29121 29101 29155
rect 29135 29152 29147 29155
rect 29178 29152 29184 29164
rect 29135 29124 29184 29152
rect 29135 29121 29147 29124
rect 29089 29115 29147 29121
rect 29178 29112 29184 29124
rect 29236 29112 29242 29164
rect 29748 29161 29776 29260
rect 32398 29248 32404 29260
rect 32456 29248 32462 29300
rect 32677 29291 32735 29297
rect 32677 29257 32689 29291
rect 32723 29288 32735 29291
rect 32858 29288 32864 29300
rect 32723 29260 32864 29288
rect 32723 29257 32735 29260
rect 32677 29251 32735 29257
rect 32858 29248 32864 29260
rect 32916 29248 32922 29300
rect 33137 29291 33195 29297
rect 33137 29257 33149 29291
rect 33183 29288 33195 29291
rect 34425 29291 34483 29297
rect 34425 29288 34437 29291
rect 33183 29260 34437 29288
rect 33183 29257 33195 29260
rect 33137 29251 33195 29257
rect 34425 29257 34437 29260
rect 34471 29257 34483 29291
rect 34425 29251 34483 29257
rect 34514 29248 34520 29300
rect 34572 29288 34578 29300
rect 35161 29291 35219 29297
rect 35161 29288 35173 29291
rect 34572 29260 35173 29288
rect 34572 29248 34578 29260
rect 35161 29257 35173 29260
rect 35207 29257 35219 29291
rect 35161 29251 35219 29257
rect 29914 29180 29920 29232
rect 29972 29220 29978 29232
rect 30009 29223 30067 29229
rect 30009 29220 30021 29223
rect 29972 29192 30021 29220
rect 29972 29180 29978 29192
rect 30009 29189 30021 29192
rect 30055 29189 30067 29223
rect 30009 29183 30067 29189
rect 31018 29180 31024 29232
rect 31076 29180 31082 29232
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 32950 29112 32956 29164
rect 33008 29152 33014 29164
rect 33045 29155 33103 29161
rect 33045 29152 33057 29155
rect 33008 29124 33057 29152
rect 33008 29112 33014 29124
rect 33045 29121 33057 29124
rect 33091 29121 33103 29155
rect 34054 29152 34060 29164
rect 34015 29124 34060 29152
rect 33045 29115 33103 29121
rect 34054 29112 34060 29124
rect 34112 29152 34118 29164
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34112 29124 34897 29152
rect 34112 29112 34118 29124
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 22428 29056 22876 29084
rect 26436 29056 27108 29084
rect 28445 29087 28503 29093
rect 22428 29044 22434 29056
rect 26436 29028 26464 29056
rect 28445 29053 28457 29087
rect 28491 29053 28503 29087
rect 28445 29047 28503 29053
rect 28534 29044 28540 29096
rect 28592 29084 28598 29096
rect 28905 29087 28963 29093
rect 28905 29084 28917 29087
rect 28592 29056 28917 29084
rect 28592 29044 28598 29056
rect 28905 29053 28917 29056
rect 28951 29053 28963 29087
rect 28905 29047 28963 29053
rect 30006 29044 30012 29096
rect 30064 29084 30070 29096
rect 31481 29087 31539 29093
rect 31481 29084 31493 29087
rect 30064 29056 31493 29084
rect 30064 29044 30070 29056
rect 31481 29053 31493 29056
rect 31527 29053 31539 29087
rect 31481 29047 31539 29053
rect 32490 29044 32496 29096
rect 32548 29084 32554 29096
rect 33229 29087 33287 29093
rect 33229 29084 33241 29087
rect 32548 29056 33241 29084
rect 32548 29044 32554 29056
rect 33229 29053 33241 29056
rect 33275 29053 33287 29087
rect 33229 29047 33287 29053
rect 33962 29044 33968 29096
rect 34020 29084 34026 29096
rect 34149 29087 34207 29093
rect 34149 29084 34161 29087
rect 34020 29056 34161 29084
rect 34020 29044 34026 29056
rect 34149 29053 34161 29056
rect 34195 29084 34207 29087
rect 34977 29087 35035 29093
rect 34977 29084 34989 29087
rect 34195 29056 34989 29084
rect 34195 29053 34207 29056
rect 34149 29047 34207 29053
rect 34977 29053 34989 29056
rect 35023 29053 35035 29087
rect 34977 29047 35035 29053
rect 35161 29087 35219 29093
rect 35161 29053 35173 29087
rect 35207 29084 35219 29087
rect 35342 29084 35348 29096
rect 35207 29056 35348 29084
rect 35207 29053 35219 29056
rect 35161 29047 35219 29053
rect 35342 29044 35348 29056
rect 35400 29044 35406 29096
rect 10413 29019 10471 29025
rect 10413 28985 10425 29019
rect 10459 29016 10471 29019
rect 11238 29016 11244 29028
rect 10459 28988 11244 29016
rect 10459 28985 10471 28988
rect 10413 28979 10471 28985
rect 11238 28976 11244 28988
rect 11296 28976 11302 29028
rect 13265 29019 13323 29025
rect 13265 28985 13277 29019
rect 13311 29016 13323 29019
rect 17954 29016 17960 29028
rect 13311 28988 17960 29016
rect 13311 28985 13323 28988
rect 13265 28979 13323 28985
rect 17954 28976 17960 28988
rect 18012 28976 18018 29028
rect 18690 28976 18696 29028
rect 18748 29016 18754 29028
rect 19245 29019 19303 29025
rect 19245 29016 19257 29019
rect 18748 28988 19257 29016
rect 18748 28976 18754 28988
rect 19245 28985 19257 28988
rect 19291 29016 19303 29019
rect 22189 29019 22247 29025
rect 22189 29016 22201 29019
rect 19291 28988 22201 29016
rect 19291 28985 19303 28988
rect 19245 28979 19303 28985
rect 22189 28985 22201 28988
rect 22235 29016 22247 29019
rect 26142 29016 26148 29028
rect 22235 28988 26148 29016
rect 22235 28985 22247 28988
rect 22189 28979 22247 28985
rect 26142 28976 26148 28988
rect 26200 29016 26206 29028
rect 26418 29016 26424 29028
rect 26200 28988 26424 29016
rect 26200 28976 26206 28988
rect 26418 28976 26424 28988
rect 26476 28976 26482 29028
rect 28718 28976 28724 29028
rect 28776 29016 28782 29028
rect 29273 29019 29331 29025
rect 29273 29016 29285 29019
rect 28776 28988 29285 29016
rect 28776 28976 28782 28988
rect 29273 28985 29285 28988
rect 29319 28985 29331 29019
rect 29273 28979 29331 28985
rect 21266 28948 21272 28960
rect 21227 28920 21272 28948
rect 21266 28908 21272 28920
rect 21324 28908 21330 28960
rect 22830 28908 22836 28960
rect 22888 28948 22894 28960
rect 26234 28948 26240 28960
rect 22888 28920 26240 28948
rect 22888 28908 22894 28920
rect 26234 28908 26240 28920
rect 26292 28908 26298 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 12529 28747 12587 28753
rect 12529 28713 12541 28747
rect 12575 28744 12587 28747
rect 12618 28744 12624 28756
rect 12575 28716 12624 28744
rect 12575 28713 12587 28716
rect 12529 28707 12587 28713
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 15470 28704 15476 28756
rect 15528 28744 15534 28756
rect 18233 28747 18291 28753
rect 18233 28744 18245 28747
rect 15528 28716 18245 28744
rect 15528 28704 15534 28716
rect 18233 28713 18245 28716
rect 18279 28713 18291 28747
rect 18233 28707 18291 28713
rect 18322 28704 18328 28756
rect 18380 28744 18386 28756
rect 18601 28747 18659 28753
rect 18601 28744 18613 28747
rect 18380 28716 18613 28744
rect 18380 28704 18386 28716
rect 18601 28713 18613 28716
rect 18647 28744 18659 28747
rect 19797 28747 19855 28753
rect 19797 28744 19809 28747
rect 18647 28716 19809 28744
rect 18647 28713 18659 28716
rect 18601 28707 18659 28713
rect 19797 28713 19809 28716
rect 19843 28744 19855 28747
rect 22738 28744 22744 28756
rect 19843 28716 22744 28744
rect 19843 28713 19855 28716
rect 19797 28707 19855 28713
rect 22738 28704 22744 28716
rect 22796 28744 22802 28756
rect 26326 28744 26332 28756
rect 22796 28716 26332 28744
rect 22796 28704 22802 28716
rect 26326 28704 26332 28716
rect 26384 28744 26390 28756
rect 26421 28747 26479 28753
rect 26421 28744 26433 28747
rect 26384 28716 26433 28744
rect 26384 28704 26390 28716
rect 26421 28713 26433 28716
rect 26467 28713 26479 28747
rect 26421 28707 26479 28713
rect 29730 28704 29736 28756
rect 29788 28744 29794 28756
rect 30101 28747 30159 28753
rect 30101 28744 30113 28747
rect 29788 28716 30113 28744
rect 29788 28704 29794 28716
rect 30101 28713 30113 28716
rect 30147 28713 30159 28747
rect 30101 28707 30159 28713
rect 30929 28747 30987 28753
rect 30929 28713 30941 28747
rect 30975 28744 30987 28747
rect 31018 28744 31024 28756
rect 30975 28716 31024 28744
rect 30975 28713 30987 28716
rect 30929 28707 30987 28713
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 34054 28704 34060 28756
rect 34112 28744 34118 28756
rect 34149 28747 34207 28753
rect 34149 28744 34161 28747
rect 34112 28716 34161 28744
rect 34112 28704 34118 28716
rect 34149 28713 34161 28716
rect 34195 28744 34207 28747
rect 34701 28747 34759 28753
rect 34701 28744 34713 28747
rect 34195 28716 34713 28744
rect 34195 28713 34207 28716
rect 34149 28707 34207 28713
rect 34701 28713 34713 28716
rect 34747 28713 34759 28747
rect 34701 28707 34759 28713
rect 34790 28704 34796 28756
rect 34848 28744 34854 28756
rect 35161 28747 35219 28753
rect 35161 28744 35173 28747
rect 34848 28716 35173 28744
rect 34848 28704 34854 28716
rect 35161 28713 35173 28716
rect 35207 28713 35219 28747
rect 35161 28707 35219 28713
rect 3786 28636 3792 28688
rect 3844 28676 3850 28688
rect 21453 28679 21511 28685
rect 3844 28648 16620 28676
rect 3844 28636 3850 28648
rect 3970 28568 3976 28620
rect 4028 28608 4034 28620
rect 9769 28611 9827 28617
rect 9769 28608 9781 28611
rect 4028 28580 9781 28608
rect 4028 28568 4034 28580
rect 9769 28577 9781 28580
rect 9815 28577 9827 28611
rect 9769 28571 9827 28577
rect 15933 28611 15991 28617
rect 15933 28577 15945 28611
rect 15979 28608 15991 28611
rect 16390 28608 16396 28620
rect 15979 28580 16396 28608
rect 15979 28577 15991 28580
rect 15933 28571 15991 28577
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 16592 28617 16620 28648
rect 21453 28645 21465 28679
rect 21499 28676 21511 28679
rect 22278 28676 22284 28688
rect 21499 28648 22284 28676
rect 21499 28645 21511 28648
rect 21453 28639 21511 28645
rect 22278 28636 22284 28648
rect 22336 28636 22342 28688
rect 23106 28636 23112 28688
rect 23164 28676 23170 28688
rect 29178 28676 29184 28688
rect 23164 28648 23244 28676
rect 23164 28636 23170 28648
rect 16577 28611 16635 28617
rect 16577 28577 16589 28611
rect 16623 28577 16635 28611
rect 18690 28608 18696 28620
rect 18651 28580 18696 28608
rect 16577 28571 16635 28577
rect 18690 28568 18696 28580
rect 18748 28568 18754 28620
rect 21082 28568 21088 28620
rect 21140 28608 21146 28620
rect 23216 28617 23244 28648
rect 28736 28648 29184 28676
rect 23201 28611 23259 28617
rect 21140 28580 21680 28608
rect 21140 28568 21146 28580
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 9309 28503 9367 28509
rect 12529 28543 12587 28549
rect 12529 28509 12541 28543
rect 12575 28540 12587 28543
rect 14182 28540 14188 28552
rect 12575 28512 14188 28540
rect 12575 28509 12587 28512
rect 12529 28503 12587 28509
rect 9324 28404 9352 28503
rect 14182 28500 14188 28512
rect 14240 28500 14246 28552
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28540 18475 28543
rect 18506 28540 18512 28552
rect 18463 28512 18512 28540
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 18506 28500 18512 28512
rect 18564 28500 18570 28552
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 20349 28543 20407 28549
rect 20349 28540 20361 28543
rect 19392 28512 20361 28540
rect 19392 28500 19398 28512
rect 20349 28509 20361 28512
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 20898 28500 20904 28552
rect 20956 28540 20962 28552
rect 21361 28543 21419 28549
rect 21361 28540 21373 28543
rect 20956 28512 21373 28540
rect 20956 28500 20962 28512
rect 21361 28509 21373 28512
rect 21407 28509 21419 28543
rect 21542 28540 21548 28552
rect 21503 28512 21548 28540
rect 21361 28503 21419 28509
rect 21542 28500 21548 28512
rect 21600 28500 21606 28552
rect 21652 28549 21680 28580
rect 23201 28577 23213 28611
rect 23247 28577 23259 28611
rect 23201 28571 23259 28577
rect 26418 28568 26424 28620
rect 26476 28608 26482 28620
rect 26513 28611 26571 28617
rect 26513 28608 26525 28611
rect 26476 28580 26525 28608
rect 26476 28568 26482 28580
rect 26513 28577 26525 28580
rect 26559 28577 26571 28611
rect 28074 28608 28080 28620
rect 26513 28571 26571 28577
rect 27448 28580 28080 28608
rect 21637 28543 21695 28549
rect 21637 28509 21649 28543
rect 21683 28509 21695 28543
rect 22830 28540 22836 28552
rect 22791 28512 22836 28540
rect 21637 28503 21695 28509
rect 22830 28500 22836 28512
rect 22888 28500 22894 28552
rect 22922 28500 22928 28552
rect 22980 28540 22986 28552
rect 23021 28545 23079 28551
rect 23021 28540 23033 28545
rect 22980 28512 23033 28540
rect 22980 28500 22986 28512
rect 23021 28511 23033 28512
rect 23067 28511 23079 28545
rect 23021 28505 23079 28511
rect 23118 28543 23176 28549
rect 23118 28509 23130 28543
rect 23164 28534 23176 28543
rect 23290 28534 23296 28552
rect 23164 28509 23296 28534
rect 23118 28506 23296 28509
rect 23118 28503 23176 28506
rect 23290 28500 23296 28506
rect 23348 28500 23354 28552
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 23566 28540 23572 28552
rect 23431 28512 23572 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 24302 28500 24308 28552
rect 24360 28540 24366 28552
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 24360 28512 24409 28540
rect 24360 28500 24366 28512
rect 24397 28509 24409 28512
rect 24443 28509 24455 28543
rect 24397 28503 24455 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28540 26111 28543
rect 26326 28540 26332 28552
rect 26099 28512 26332 28540
rect 26099 28509 26111 28512
rect 26053 28503 26111 28509
rect 26326 28500 26332 28512
rect 26384 28500 26390 28552
rect 27246 28500 27252 28552
rect 27304 28540 27310 28552
rect 27448 28549 27476 28580
rect 28074 28568 28080 28580
rect 28132 28568 28138 28620
rect 27433 28543 27491 28549
rect 27433 28540 27445 28543
rect 27304 28512 27445 28540
rect 27304 28500 27310 28512
rect 27433 28509 27445 28512
rect 27479 28509 27491 28543
rect 27433 28503 27491 28509
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28540 27767 28543
rect 27985 28543 28043 28549
rect 27755 28512 27936 28540
rect 27755 28509 27767 28512
rect 27709 28503 27767 28509
rect 9493 28475 9551 28481
rect 9493 28441 9505 28475
rect 9539 28472 9551 28475
rect 10042 28472 10048 28484
rect 9539 28444 10048 28472
rect 9539 28441 9551 28444
rect 9493 28435 9551 28441
rect 10042 28432 10048 28444
rect 10100 28432 10106 28484
rect 14553 28475 14611 28481
rect 14553 28441 14565 28475
rect 14599 28472 14611 28475
rect 16114 28472 16120 28484
rect 14599 28444 15608 28472
rect 16075 28444 16120 28472
rect 14599 28441 14611 28444
rect 14553 28435 14611 28441
rect 10410 28404 10416 28416
rect 9324 28376 10416 28404
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 14642 28404 14648 28416
rect 14603 28376 14648 28404
rect 14642 28364 14648 28376
rect 14700 28364 14706 28416
rect 15580 28404 15608 28444
rect 16114 28432 16120 28444
rect 16172 28432 16178 28484
rect 18230 28432 18236 28484
rect 18288 28472 18294 28484
rect 19705 28475 19763 28481
rect 19705 28472 19717 28475
rect 18288 28444 19717 28472
rect 18288 28432 18294 28444
rect 19705 28441 19717 28444
rect 19751 28472 19763 28475
rect 21266 28472 21272 28484
rect 19751 28444 21272 28472
rect 19751 28441 19763 28444
rect 19705 28435 19763 28441
rect 21266 28432 21272 28444
rect 21324 28432 21330 28484
rect 26145 28475 26203 28481
rect 26145 28441 26157 28475
rect 26191 28472 26203 28475
rect 27614 28472 27620 28484
rect 26191 28444 27620 28472
rect 26191 28441 26203 28444
rect 26145 28435 26203 28441
rect 27614 28432 27620 28444
rect 27672 28472 27678 28484
rect 27798 28472 27804 28484
rect 27672 28444 27804 28472
rect 27672 28432 27678 28444
rect 27798 28432 27804 28444
rect 27856 28432 27862 28484
rect 19242 28404 19248 28416
rect 15580 28376 19248 28404
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 20441 28407 20499 28413
rect 20441 28373 20453 28407
rect 20487 28404 20499 28407
rect 20530 28404 20536 28416
rect 20487 28376 20536 28404
rect 20487 28373 20499 28376
rect 20441 28367 20499 28373
rect 20530 28364 20536 28376
rect 20588 28364 20594 28416
rect 21174 28404 21180 28416
rect 21135 28376 21180 28404
rect 21174 28364 21180 28376
rect 21232 28364 21238 28416
rect 22922 28364 22928 28416
rect 22980 28404 22986 28416
rect 23569 28407 23627 28413
rect 23569 28404 23581 28407
rect 22980 28376 23581 28404
rect 22980 28364 22986 28376
rect 23569 28373 23581 28376
rect 23615 28373 23627 28407
rect 24486 28404 24492 28416
rect 24447 28376 24492 28404
rect 23569 28367 23627 28373
rect 24486 28364 24492 28376
rect 24544 28364 24550 28416
rect 25314 28364 25320 28416
rect 25372 28404 25378 28416
rect 25777 28407 25835 28413
rect 25777 28404 25789 28407
rect 25372 28376 25789 28404
rect 25372 28364 25378 28376
rect 25777 28373 25789 28376
rect 25823 28373 25835 28407
rect 25777 28367 25835 28373
rect 26237 28407 26295 28413
rect 26237 28373 26249 28407
rect 26283 28404 26295 28407
rect 26510 28404 26516 28416
rect 26283 28376 26516 28404
rect 26283 28373 26295 28376
rect 26237 28367 26295 28373
rect 26510 28364 26516 28376
rect 26568 28404 26574 28416
rect 27062 28404 27068 28416
rect 26568 28376 27068 28404
rect 26568 28364 26574 28376
rect 27062 28364 27068 28376
rect 27120 28404 27126 28416
rect 27525 28407 27583 28413
rect 27525 28404 27537 28407
rect 27120 28376 27537 28404
rect 27120 28364 27126 28376
rect 27525 28373 27537 28376
rect 27571 28373 27583 28407
rect 27908 28404 27936 28512
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28540 28227 28543
rect 28736 28540 28764 28648
rect 29178 28636 29184 28648
rect 29236 28636 29242 28688
rect 28902 28608 28908 28620
rect 28815 28580 28908 28608
rect 28902 28568 28908 28580
rect 28960 28608 28966 28620
rect 29641 28611 29699 28617
rect 29641 28608 29653 28611
rect 28960 28580 29653 28608
rect 28960 28568 28966 28580
rect 29641 28577 29653 28580
rect 29687 28577 29699 28611
rect 32398 28608 32404 28620
rect 32359 28580 32404 28608
rect 29641 28571 29699 28577
rect 32398 28568 32404 28580
rect 32456 28568 32462 28620
rect 33870 28568 33876 28620
rect 33928 28608 33934 28620
rect 34793 28611 34851 28617
rect 34793 28608 34805 28611
rect 33928 28580 34805 28608
rect 33928 28568 33934 28580
rect 34793 28577 34805 28580
rect 34839 28577 34851 28611
rect 34793 28571 34851 28577
rect 28813 28543 28871 28549
rect 28813 28540 28825 28543
rect 28215 28512 28825 28540
rect 28215 28509 28227 28512
rect 28169 28503 28227 28509
rect 28813 28509 28825 28512
rect 28859 28509 28871 28543
rect 28813 28503 28871 28509
rect 28997 28543 29055 28549
rect 28997 28509 29009 28543
rect 29043 28509 29055 28543
rect 28997 28503 29055 28509
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 30006 28540 30012 28552
rect 29779 28512 30012 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 28000 28472 28028 28503
rect 28534 28472 28540 28484
rect 28000 28444 28540 28472
rect 28534 28432 28540 28444
rect 28592 28472 28598 28484
rect 29012 28472 29040 28503
rect 28592 28444 29040 28472
rect 28592 28432 28598 28444
rect 28350 28404 28356 28416
rect 27908 28376 28356 28404
rect 27525 28367 27583 28373
rect 28350 28364 28356 28376
rect 28408 28404 28414 28416
rect 29748 28404 29776 28503
rect 30006 28500 30012 28512
rect 30064 28500 30070 28552
rect 30837 28543 30895 28549
rect 30837 28509 30849 28543
rect 30883 28540 30895 28543
rect 30926 28540 30932 28552
rect 30883 28512 30932 28540
rect 30883 28509 30895 28512
rect 30837 28503 30895 28509
rect 30926 28500 30932 28512
rect 30984 28500 30990 28552
rect 31754 28500 31760 28552
rect 31812 28540 31818 28552
rect 34977 28543 35035 28549
rect 31812 28512 31857 28540
rect 31812 28500 31818 28512
rect 34977 28509 34989 28543
rect 35023 28540 35035 28543
rect 35342 28540 35348 28552
rect 35023 28512 35348 28540
rect 35023 28509 35035 28512
rect 34977 28503 35035 28509
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 46934 28500 46940 28552
rect 46992 28540 46998 28552
rect 47673 28543 47731 28549
rect 47673 28540 47685 28543
rect 46992 28512 47685 28540
rect 46992 28500 46998 28512
rect 47673 28509 47685 28512
rect 47719 28509 47731 28543
rect 47673 28503 47731 28509
rect 32582 28432 32588 28484
rect 32640 28472 32646 28484
rect 32677 28475 32735 28481
rect 32677 28472 32689 28475
rect 32640 28444 32689 28472
rect 32640 28432 32646 28444
rect 32677 28441 32689 28444
rect 32723 28441 32735 28475
rect 32677 28435 32735 28441
rect 33134 28432 33140 28484
rect 33192 28432 33198 28484
rect 34698 28472 34704 28484
rect 34659 28444 34704 28472
rect 34698 28432 34704 28444
rect 34756 28432 34762 28484
rect 31846 28404 31852 28416
rect 28408 28376 29776 28404
rect 31807 28376 31852 28404
rect 28408 28364 28414 28376
rect 31846 28364 31852 28376
rect 31904 28364 31910 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 10042 28200 10048 28212
rect 10003 28172 10048 28200
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 16025 28203 16083 28209
rect 16025 28169 16037 28203
rect 16071 28200 16083 28203
rect 16114 28200 16120 28212
rect 16071 28172 16120 28200
rect 16071 28169 16083 28172
rect 16025 28163 16083 28169
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 16758 28200 16764 28212
rect 16719 28172 16764 28200
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 17954 28200 17960 28212
rect 17915 28172 17960 28200
rect 17954 28160 17960 28172
rect 18012 28160 18018 28212
rect 18966 28160 18972 28212
rect 19024 28200 19030 28212
rect 22646 28200 22652 28212
rect 19024 28172 22652 28200
rect 19024 28160 19030 28172
rect 9968 28104 15332 28132
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28064 8263 28067
rect 8478 28064 8484 28076
rect 8251 28036 8484 28064
rect 8251 28033 8263 28036
rect 8205 28027 8263 28033
rect 8478 28024 8484 28036
rect 8536 28024 8542 28076
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 9309 28067 9367 28073
rect 9309 28064 9321 28067
rect 9272 28036 9321 28064
rect 9272 28024 9278 28036
rect 9309 28033 9321 28036
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 9766 28024 9772 28076
rect 9824 28064 9830 28076
rect 9968 28073 9996 28104
rect 15304 28076 15332 28104
rect 18046 28092 18052 28144
rect 18104 28132 18110 28144
rect 18104 28104 18460 28132
rect 18104 28092 18110 28104
rect 9953 28067 10011 28073
rect 9953 28064 9965 28067
rect 9824 28036 9965 28064
rect 9824 28024 9830 28036
rect 9953 28033 9965 28036
rect 9999 28033 10011 28067
rect 11882 28064 11888 28076
rect 11843 28036 11888 28064
rect 9953 28027 10011 28033
rect 11882 28024 11888 28036
rect 11940 28064 11946 28076
rect 12158 28064 12164 28076
rect 11940 28036 12164 28064
rect 11940 28024 11946 28036
rect 12158 28024 12164 28036
rect 12216 28024 12222 28076
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 13446 28064 13452 28076
rect 13407 28036 13452 28064
rect 12897 28027 12955 28033
rect 11974 27996 11980 28008
rect 11935 27968 11980 27996
rect 11974 27956 11980 27968
rect 12032 27956 12038 28008
rect 12912 27996 12940 28027
rect 13446 28024 13452 28036
rect 13504 28024 13510 28076
rect 15286 28024 15292 28076
rect 15344 28064 15350 28076
rect 15933 28067 15991 28073
rect 15933 28064 15945 28067
rect 15344 28036 15945 28064
rect 15344 28024 15350 28036
rect 15933 28033 15945 28036
rect 15979 28064 15991 28067
rect 16022 28064 16028 28076
rect 15979 28036 16028 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16669 28067 16727 28073
rect 16669 28033 16681 28067
rect 16715 28064 16727 28067
rect 17034 28064 17040 28076
rect 16715 28036 17040 28064
rect 16715 28033 16727 28036
rect 16669 28027 16727 28033
rect 17034 28024 17040 28036
rect 17092 28024 17098 28076
rect 18230 28064 18236 28076
rect 18191 28036 18236 28064
rect 18230 28024 18236 28036
rect 18288 28024 18294 28076
rect 18432 28073 18460 28104
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28064 18475 28067
rect 19058 28064 19064 28076
rect 18463 28036 19064 28064
rect 18463 28033 18475 28036
rect 18417 28027 18475 28033
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 19260 28073 19288 28172
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 23290 28160 23296 28212
rect 23348 28200 23354 28212
rect 24397 28203 24455 28209
rect 24397 28200 24409 28203
rect 23348 28172 24409 28200
rect 23348 28160 23354 28172
rect 24397 28169 24409 28172
rect 24443 28200 24455 28203
rect 27246 28200 27252 28212
rect 24443 28172 27252 28200
rect 24443 28169 24455 28172
rect 24397 28163 24455 28169
rect 27246 28160 27252 28172
rect 27304 28160 27310 28212
rect 28258 28200 28264 28212
rect 27356 28172 27660 28200
rect 28219 28172 28264 28200
rect 20530 28092 20536 28144
rect 20588 28092 20594 28144
rect 21266 28092 21272 28144
rect 21324 28132 21330 28144
rect 21821 28135 21879 28141
rect 21821 28132 21833 28135
rect 21324 28104 21833 28132
rect 21324 28092 21330 28104
rect 21821 28101 21833 28104
rect 21867 28101 21879 28135
rect 21821 28095 21879 28101
rect 22189 28135 22247 28141
rect 22189 28101 22201 28135
rect 22235 28132 22247 28135
rect 22370 28132 22376 28144
rect 22235 28104 22376 28132
rect 22235 28101 22247 28104
rect 22189 28095 22247 28101
rect 22370 28092 22376 28104
rect 22428 28092 22434 28144
rect 22922 28132 22928 28144
rect 22883 28104 22928 28132
rect 22922 28092 22928 28104
rect 22980 28092 22986 28144
rect 24486 28132 24492 28144
rect 24150 28104 24492 28132
rect 24486 28092 24492 28104
rect 24544 28092 24550 28144
rect 24857 28135 24915 28141
rect 24857 28101 24869 28135
rect 24903 28132 24915 28135
rect 25501 28135 25559 28141
rect 25501 28132 25513 28135
rect 24903 28104 25513 28132
rect 24903 28101 24915 28104
rect 24857 28095 24915 28101
rect 25501 28101 25513 28104
rect 25547 28132 25559 28135
rect 27356 28132 27384 28172
rect 25547 28104 27384 28132
rect 27632 28132 27660 28172
rect 28258 28160 28264 28172
rect 28316 28160 28322 28212
rect 32582 28200 32588 28212
rect 32543 28172 32588 28200
rect 32582 28160 32588 28172
rect 32640 28160 32646 28212
rect 47026 28200 47032 28212
rect 41386 28172 47032 28200
rect 41386 28132 41414 28172
rect 47026 28160 47032 28172
rect 47084 28160 47090 28212
rect 27632 28104 41414 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28033 19303 28067
rect 22002 28064 22008 28076
rect 19245 28027 19303 28033
rect 20732 28036 22008 28064
rect 14182 27996 14188 28008
rect 12912 27968 14188 27996
rect 14182 27956 14188 27968
rect 14240 27956 14246 28008
rect 17865 27999 17923 28005
rect 17865 27965 17877 27999
rect 17911 27965 17923 27999
rect 18138 27996 18144 28008
rect 18099 27968 18144 27996
rect 17865 27959 17923 27965
rect 17880 27928 17908 27959
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 19518 27996 19524 28008
rect 19479 27968 19524 27996
rect 19518 27956 19524 27968
rect 19576 27956 19582 28008
rect 18598 27928 18604 27940
rect 17880 27900 18604 27928
rect 18598 27888 18604 27900
rect 18656 27888 18662 27940
rect 8294 27860 8300 27872
rect 8255 27832 8300 27860
rect 8294 27820 8300 27832
rect 8352 27820 8358 27872
rect 9401 27863 9459 27869
rect 9401 27829 9413 27863
rect 9447 27860 9459 27863
rect 9674 27860 9680 27872
rect 9447 27832 9680 27860
rect 9447 27829 9459 27832
rect 9401 27823 9459 27829
rect 9674 27820 9680 27832
rect 9732 27820 9738 27872
rect 12158 27860 12164 27872
rect 12119 27832 12164 27860
rect 12158 27820 12164 27832
rect 12216 27820 12222 27872
rect 12710 27860 12716 27872
rect 12671 27832 12716 27860
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 13538 27860 13544 27872
rect 13499 27832 13544 27860
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 17310 27820 17316 27872
rect 17368 27860 17374 27872
rect 17681 27863 17739 27869
rect 17681 27860 17693 27863
rect 17368 27832 17693 27860
rect 17368 27820 17374 27832
rect 17681 27829 17693 27832
rect 17727 27829 17739 27863
rect 17681 27823 17739 27829
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 20732 27860 20760 28036
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27433 28067 27491 28073
rect 27356 28064 27445 28067
rect 27120 28039 27445 28064
rect 27120 28036 27384 28039
rect 27120 28024 27126 28036
rect 27433 28033 27445 28039
rect 27479 28033 27491 28067
rect 27433 28027 27491 28033
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28064 27583 28067
rect 27571 28033 27584 28064
rect 27525 28027 27584 28033
rect 20993 27999 21051 28005
rect 20993 27965 21005 27999
rect 21039 27996 21051 27999
rect 21082 27996 21088 28008
rect 21039 27968 21088 27996
rect 21039 27965 21051 27968
rect 20993 27959 21051 27965
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 22646 27996 22652 28008
rect 22607 27968 22652 27996
rect 22646 27956 22652 27968
rect 22704 27956 22710 28008
rect 25590 27996 25596 28008
rect 25551 27968 25596 27996
rect 25590 27956 25596 27968
rect 25648 27956 25654 28008
rect 25685 27999 25743 28005
rect 25685 27965 25697 27999
rect 25731 27965 25743 27999
rect 25685 27959 25743 27965
rect 25700 27928 25728 27959
rect 23952 27900 25728 27928
rect 19116 27832 20760 27860
rect 19116 27820 19122 27832
rect 21726 27820 21732 27872
rect 21784 27860 21790 27872
rect 23952 27860 23980 27900
rect 27338 27888 27344 27940
rect 27396 27928 27402 27940
rect 27556 27928 27584 28027
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 27801 28067 27859 28073
rect 27672 28036 27717 28064
rect 27672 28024 27678 28036
rect 27801 28033 27813 28067
rect 27847 28064 27859 28067
rect 27982 28064 27988 28076
rect 27847 28036 27988 28064
rect 27847 28033 27859 28036
rect 27801 28027 27859 28033
rect 27982 28024 27988 28036
rect 28040 28024 28046 28076
rect 28350 28024 28356 28076
rect 28408 28064 28414 28076
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 28408 28036 28457 28064
rect 28408 28024 28414 28036
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 28721 28067 28779 28073
rect 28721 28033 28733 28067
rect 28767 28033 28779 28067
rect 32766 28064 32772 28076
rect 32727 28036 32772 28064
rect 28721 28027 28779 28033
rect 28074 27956 28080 28008
rect 28132 27996 28138 28008
rect 28736 27996 28764 28027
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 47581 28067 47639 28073
rect 47581 28033 47593 28067
rect 47627 28064 47639 28067
rect 47670 28064 47676 28076
rect 47627 28036 47676 28064
rect 47627 28033 47639 28036
rect 47581 28027 47639 28033
rect 47670 28024 47676 28036
rect 47728 28024 47734 28076
rect 28132 27968 28764 27996
rect 28132 27956 28138 27968
rect 27396 27900 27584 27928
rect 27396 27888 27402 27900
rect 28258 27888 28264 27940
rect 28316 27928 28322 27940
rect 28534 27928 28540 27940
rect 28316 27900 28540 27928
rect 28316 27888 28322 27900
rect 28534 27888 28540 27900
rect 28592 27888 28598 27940
rect 28629 27931 28687 27937
rect 28629 27897 28641 27931
rect 28675 27928 28687 27931
rect 29178 27928 29184 27940
rect 28675 27900 29184 27928
rect 28675 27897 28687 27900
rect 28629 27891 28687 27897
rect 29178 27888 29184 27900
rect 29236 27888 29242 27940
rect 25130 27860 25136 27872
rect 21784 27832 23980 27860
rect 25091 27832 25136 27860
rect 21784 27820 21790 27832
rect 25130 27820 25136 27832
rect 25188 27820 25194 27872
rect 27157 27863 27215 27869
rect 27157 27829 27169 27863
rect 27203 27860 27215 27863
rect 28442 27860 28448 27872
rect 27203 27832 28448 27860
rect 27203 27829 27215 27832
rect 27157 27823 27215 27829
rect 28442 27820 28448 27832
rect 28500 27820 28506 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 11964 27659 12022 27665
rect 11964 27625 11976 27659
rect 12010 27656 12022 27659
rect 12158 27656 12164 27668
rect 12010 27628 12164 27656
rect 12010 27625 12022 27628
rect 11964 27619 12022 27625
rect 12158 27616 12164 27628
rect 12216 27616 12222 27668
rect 19518 27616 19524 27668
rect 19576 27656 19582 27668
rect 19981 27659 20039 27665
rect 19981 27656 19993 27659
rect 19576 27628 19993 27656
rect 19576 27616 19582 27628
rect 19981 27625 19993 27628
rect 20027 27625 20039 27659
rect 25590 27656 25596 27668
rect 25551 27628 25596 27656
rect 19981 27619 20039 27625
rect 25590 27616 25596 27628
rect 25648 27616 25654 27668
rect 26602 27656 26608 27668
rect 26436 27628 26608 27656
rect 26326 27588 26332 27600
rect 26287 27560 26332 27588
rect 26326 27548 26332 27560
rect 26384 27548 26390 27600
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 8941 27523 8999 27529
rect 8941 27520 8953 27523
rect 8352 27492 8953 27520
rect 8352 27480 8358 27492
rect 8941 27489 8953 27492
rect 8987 27489 8999 27523
rect 8941 27483 8999 27489
rect 11701 27523 11759 27529
rect 11701 27489 11713 27523
rect 11747 27520 11759 27523
rect 12710 27520 12716 27532
rect 11747 27492 12716 27520
rect 11747 27489 11759 27492
rect 11701 27483 11759 27489
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 15194 27480 15200 27532
rect 15252 27520 15258 27532
rect 15838 27520 15844 27532
rect 15252 27492 15844 27520
rect 15252 27480 15258 27492
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 17954 27480 17960 27532
rect 18012 27520 18018 27532
rect 18012 27492 18460 27520
rect 18012 27480 18018 27492
rect 8386 27452 8392 27464
rect 8347 27424 8392 27452
rect 8386 27412 8392 27424
rect 8444 27412 8450 27464
rect 14182 27452 14188 27464
rect 14143 27424 14188 27452
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27452 14427 27455
rect 14829 27455 14887 27461
rect 14829 27452 14841 27455
rect 14415 27424 14841 27452
rect 14415 27421 14427 27424
rect 14369 27415 14427 27421
rect 14829 27421 14841 27424
rect 14875 27421 14887 27455
rect 17034 27452 17040 27464
rect 16995 27424 17040 27452
rect 14829 27415 14887 27421
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 18046 27412 18052 27464
rect 18104 27452 18110 27464
rect 18432 27461 18460 27492
rect 21174 27480 21180 27532
rect 21232 27520 21238 27532
rect 21269 27523 21327 27529
rect 21269 27520 21281 27523
rect 21232 27492 21281 27520
rect 21232 27480 21238 27492
rect 21269 27489 21281 27492
rect 21315 27489 21327 27523
rect 21269 27483 21327 27489
rect 21453 27523 21511 27529
rect 21453 27489 21465 27523
rect 21499 27520 21511 27523
rect 21726 27520 21732 27532
rect 21499 27492 21732 27520
rect 21499 27489 21511 27492
rect 21453 27483 21511 27489
rect 21726 27480 21732 27492
rect 21784 27480 21790 27532
rect 25314 27520 25320 27532
rect 25275 27492 25320 27520
rect 25314 27480 25320 27492
rect 25372 27480 25378 27532
rect 26436 27520 26464 27628
rect 26602 27616 26608 27628
rect 26660 27656 26666 27668
rect 27249 27659 27307 27665
rect 27249 27656 27261 27659
rect 26660 27628 27261 27656
rect 26660 27616 26666 27628
rect 27249 27625 27261 27628
rect 27295 27625 27307 27659
rect 27249 27619 27307 27625
rect 26694 27548 26700 27600
rect 26752 27588 26758 27600
rect 27706 27588 27712 27600
rect 26752 27560 27568 27588
rect 27667 27560 27712 27588
rect 26752 27548 26758 27560
rect 26252 27492 26464 27520
rect 18233 27455 18291 27461
rect 18233 27452 18245 27455
rect 18104 27424 18245 27452
rect 18104 27412 18110 27424
rect 18233 27421 18245 27424
rect 18279 27421 18291 27455
rect 18233 27415 18291 27421
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18417 27455 18475 27461
rect 18417 27421 18429 27455
rect 18463 27421 18475 27455
rect 18598 27452 18604 27464
rect 18559 27424 18604 27452
rect 18417 27415 18475 27421
rect 9217 27387 9275 27393
rect 9217 27384 9229 27387
rect 8220 27356 9229 27384
rect 8220 27325 8248 27356
rect 9217 27353 9229 27356
rect 9263 27353 9275 27387
rect 9217 27347 9275 27353
rect 9674 27344 9680 27396
rect 9732 27344 9738 27396
rect 13538 27384 13544 27396
rect 13202 27356 13544 27384
rect 13538 27344 13544 27356
rect 13596 27344 13602 27396
rect 14200 27384 14228 27412
rect 14550 27384 14556 27396
rect 14200 27356 14556 27384
rect 14550 27344 14556 27356
rect 14608 27344 14614 27396
rect 15105 27387 15163 27393
rect 15105 27353 15117 27387
rect 15151 27384 15163 27387
rect 15194 27384 15200 27396
rect 15151 27356 15200 27384
rect 15151 27353 15163 27356
rect 15105 27347 15163 27353
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 17129 27387 17187 27393
rect 17129 27384 17141 27387
rect 16330 27356 17141 27384
rect 17129 27353 17141 27356
rect 17175 27353 17187 27387
rect 17129 27347 17187 27353
rect 18340 27328 18368 27415
rect 18598 27412 18604 27424
rect 18656 27412 18662 27464
rect 19334 27452 19340 27464
rect 19295 27424 19340 27452
rect 19334 27412 19340 27424
rect 19392 27412 19398 27464
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27452 20223 27455
rect 20211 27424 20852 27452
rect 20211 27421 20223 27424
rect 20165 27415 20223 27421
rect 8205 27319 8263 27325
rect 8205 27285 8217 27319
rect 8251 27285 8263 27319
rect 8205 27279 8263 27285
rect 10689 27319 10747 27325
rect 10689 27285 10701 27319
rect 10735 27316 10747 27319
rect 11330 27316 11336 27328
rect 10735 27288 11336 27316
rect 10735 27285 10747 27288
rect 10689 27279 10747 27285
rect 11330 27276 11336 27288
rect 11388 27276 11394 27328
rect 11882 27276 11888 27328
rect 11940 27316 11946 27328
rect 13449 27319 13507 27325
rect 13449 27316 13461 27319
rect 11940 27288 13461 27316
rect 11940 27276 11946 27288
rect 13449 27285 13461 27288
rect 13495 27285 13507 27319
rect 13449 27279 13507 27285
rect 15838 27276 15844 27328
rect 15896 27316 15902 27328
rect 16577 27319 16635 27325
rect 16577 27316 16589 27319
rect 15896 27288 16589 27316
rect 15896 27276 15902 27288
rect 16577 27285 16589 27288
rect 16623 27316 16635 27319
rect 16758 27316 16764 27328
rect 16623 27288 16764 27316
rect 16623 27285 16635 27288
rect 16577 27279 16635 27285
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 17954 27316 17960 27328
rect 17915 27288 17960 27316
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 18322 27276 18328 27328
rect 18380 27276 18386 27328
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 20070 27316 20076 27328
rect 19475 27288 20076 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 20070 27276 20076 27288
rect 20128 27276 20134 27328
rect 20824 27325 20852 27424
rect 22002 27412 22008 27464
rect 22060 27452 22066 27464
rect 22097 27455 22155 27461
rect 22097 27452 22109 27455
rect 22060 27424 22109 27452
rect 22060 27412 22066 27424
rect 22097 27421 22109 27424
rect 22143 27421 22155 27455
rect 22097 27415 22155 27421
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 25130 27452 25136 27464
rect 24627 27424 25136 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 26252 27461 26280 27492
rect 27246 27480 27252 27532
rect 27304 27520 27310 27532
rect 27341 27523 27399 27529
rect 27341 27520 27353 27523
rect 27304 27492 27353 27520
rect 27304 27480 27310 27492
rect 27341 27489 27353 27492
rect 27387 27489 27399 27523
rect 27540 27520 27568 27560
rect 27706 27548 27712 27560
rect 27764 27548 27770 27600
rect 28718 27588 28724 27600
rect 28679 27560 28724 27588
rect 28718 27548 28724 27560
rect 28776 27548 28782 27600
rect 33045 27591 33103 27597
rect 33045 27557 33057 27591
rect 33091 27588 33103 27591
rect 33134 27588 33140 27600
rect 33091 27560 33140 27588
rect 33091 27557 33103 27560
rect 33045 27551 33103 27557
rect 33134 27548 33140 27560
rect 33192 27548 33198 27600
rect 46934 27588 46940 27600
rect 33520 27560 40356 27588
rect 28813 27523 28871 27529
rect 27540 27492 28672 27520
rect 27341 27483 27399 27489
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 26237 27455 26295 27461
rect 26237 27421 26249 27455
rect 26283 27421 26295 27455
rect 27525 27455 27583 27461
rect 27525 27452 27537 27455
rect 26237 27415 26295 27421
rect 26344 27424 27537 27452
rect 21542 27344 21548 27396
rect 21600 27384 21606 27396
rect 22281 27387 22339 27393
rect 22281 27384 22293 27387
rect 21600 27356 22293 27384
rect 21600 27344 21606 27356
rect 22281 27353 22293 27356
rect 22327 27384 22339 27387
rect 25240 27384 25268 27415
rect 25314 27384 25320 27396
rect 22327 27356 24532 27384
rect 25227 27356 25320 27384
rect 22327 27353 22339 27356
rect 22281 27347 22339 27353
rect 20809 27319 20867 27325
rect 20809 27285 20821 27319
rect 20855 27285 20867 27319
rect 20809 27279 20867 27285
rect 21082 27276 21088 27328
rect 21140 27316 21146 27328
rect 21177 27319 21235 27325
rect 21177 27316 21189 27319
rect 21140 27288 21189 27316
rect 21140 27276 21146 27288
rect 21177 27285 21189 27288
rect 21223 27285 21235 27319
rect 21177 27279 21235 27285
rect 23842 27276 23848 27328
rect 23900 27316 23906 27328
rect 24397 27319 24455 27325
rect 24397 27316 24409 27319
rect 23900 27288 24409 27316
rect 23900 27276 23906 27288
rect 24397 27285 24409 27288
rect 24443 27285 24455 27319
rect 24504 27316 24532 27356
rect 25314 27344 25320 27356
rect 25372 27384 25378 27396
rect 26344 27384 26372 27424
rect 27525 27421 27537 27424
rect 27571 27421 27583 27455
rect 27525 27415 27583 27421
rect 28350 27412 28356 27464
rect 28408 27412 28414 27464
rect 28442 27412 28448 27464
rect 28500 27452 28506 27464
rect 28537 27455 28595 27461
rect 28537 27452 28549 27455
rect 28500 27424 28549 27452
rect 28500 27412 28506 27424
rect 28537 27421 28549 27424
rect 28583 27421 28595 27455
rect 28537 27415 28595 27421
rect 25372 27356 26372 27384
rect 27249 27387 27307 27393
rect 25372 27344 25378 27356
rect 27249 27353 27261 27387
rect 27295 27384 27307 27387
rect 28368 27384 28396 27412
rect 27295 27356 28396 27384
rect 28644 27384 28672 27492
rect 28813 27489 28825 27523
rect 28859 27520 28871 27523
rect 28902 27520 28908 27532
rect 28859 27492 28908 27520
rect 28859 27489 28871 27492
rect 28813 27483 28871 27489
rect 28902 27480 28908 27492
rect 28960 27480 28966 27532
rect 30561 27523 30619 27529
rect 30561 27489 30573 27523
rect 30607 27520 30619 27523
rect 31570 27520 31576 27532
rect 30607 27492 31576 27520
rect 30607 27489 30619 27492
rect 30561 27483 30619 27489
rect 31570 27480 31576 27492
rect 31628 27520 31634 27532
rect 31846 27520 31852 27532
rect 31628 27492 31852 27520
rect 31628 27480 31634 27492
rect 31846 27480 31852 27492
rect 31904 27480 31910 27532
rect 30742 27452 30748 27464
rect 30703 27424 30748 27452
rect 30742 27412 30748 27424
rect 30800 27412 30806 27464
rect 31662 27412 31668 27464
rect 31720 27452 31726 27464
rect 32953 27455 33011 27461
rect 32953 27452 32965 27455
rect 31720 27424 32965 27452
rect 31720 27412 31726 27424
rect 32953 27421 32965 27424
rect 32999 27421 33011 27455
rect 32953 27415 33011 27421
rect 33520 27384 33548 27560
rect 33962 27520 33968 27532
rect 33923 27492 33968 27520
rect 33962 27480 33968 27492
rect 34020 27480 34026 27532
rect 36170 27520 36176 27532
rect 36131 27492 36176 27520
rect 36170 27480 36176 27492
rect 36228 27480 36234 27532
rect 39853 27523 39911 27529
rect 39853 27489 39865 27523
rect 39899 27520 39911 27523
rect 40126 27520 40132 27532
rect 39899 27492 40132 27520
rect 39899 27489 39911 27492
rect 39853 27483 39911 27489
rect 40126 27480 40132 27492
rect 40184 27480 40190 27532
rect 40328 27529 40356 27560
rect 46308 27560 46940 27588
rect 46308 27529 46336 27560
rect 46934 27548 46940 27560
rect 46992 27548 46998 27600
rect 40313 27523 40371 27529
rect 40313 27489 40325 27523
rect 40359 27489 40371 27523
rect 40313 27483 40371 27489
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46293 27483 46351 27489
rect 46477 27523 46535 27529
rect 46477 27489 46489 27523
rect 46523 27520 46535 27523
rect 47670 27520 47676 27532
rect 46523 27492 47676 27520
rect 46523 27489 46535 27492
rect 46477 27483 46535 27489
rect 47670 27480 47676 27492
rect 47728 27480 47734 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 33781 27455 33839 27461
rect 33781 27421 33793 27455
rect 33827 27452 33839 27455
rect 33870 27452 33876 27464
rect 33827 27424 33876 27452
rect 33827 27421 33839 27424
rect 33781 27415 33839 27421
rect 33870 27412 33876 27424
rect 33928 27412 33934 27464
rect 35342 27452 35348 27464
rect 35303 27424 35348 27452
rect 35342 27412 35348 27424
rect 35400 27412 35406 27464
rect 28644 27356 33548 27384
rect 33597 27387 33655 27393
rect 27295 27353 27307 27356
rect 27249 27347 27307 27353
rect 33597 27353 33609 27387
rect 33643 27384 33655 27387
rect 34054 27384 34060 27396
rect 33643 27356 34060 27384
rect 33643 27353 33655 27356
rect 33597 27347 33655 27353
rect 34054 27344 34060 27356
rect 34112 27384 34118 27396
rect 34698 27384 34704 27396
rect 34112 27356 34704 27384
rect 34112 27344 34118 27356
rect 34698 27344 34704 27356
rect 34756 27344 34762 27396
rect 40034 27384 40040 27396
rect 39995 27356 40040 27384
rect 40034 27344 40040 27356
rect 40092 27344 40098 27396
rect 27062 27316 27068 27328
rect 24504 27288 27068 27316
rect 24397 27279 24455 27285
rect 27062 27276 27068 27288
rect 27120 27276 27126 27328
rect 28074 27276 28080 27328
rect 28132 27316 28138 27328
rect 28353 27319 28411 27325
rect 28353 27316 28365 27319
rect 28132 27288 28365 27316
rect 28132 27276 28138 27288
rect 28353 27285 28365 27288
rect 28399 27285 28411 27319
rect 28353 27279 28411 27285
rect 30929 27319 30987 27325
rect 30929 27285 30941 27319
rect 30975 27316 30987 27319
rect 31386 27316 31392 27328
rect 30975 27288 31392 27316
rect 30975 27285 30987 27288
rect 30929 27279 30987 27285
rect 31386 27276 31392 27288
rect 31444 27276 31450 27328
rect 36170 27276 36176 27328
rect 36228 27316 36234 27328
rect 47578 27316 47584 27328
rect 36228 27288 47584 27316
rect 36228 27276 36234 27288
rect 47578 27276 47584 27288
rect 47636 27276 47642 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 9677 27115 9735 27121
rect 9677 27112 9689 27115
rect 8444 27084 9689 27112
rect 8444 27072 8450 27084
rect 9677 27081 9689 27084
rect 9723 27081 9735 27115
rect 9677 27075 9735 27081
rect 10689 27115 10747 27121
rect 10689 27081 10701 27115
rect 10735 27112 10747 27115
rect 10778 27112 10784 27124
rect 10735 27084 10784 27112
rect 10735 27081 10747 27084
rect 10689 27075 10747 27081
rect 10778 27072 10784 27084
rect 10836 27072 10842 27124
rect 13173 27115 13231 27121
rect 13173 27112 13185 27115
rect 10888 27084 13185 27112
rect 10410 27044 10416 27056
rect 10371 27016 10416 27044
rect 10410 27004 10416 27016
rect 10468 27004 10474 27056
rect 10888 27044 10916 27084
rect 13173 27081 13185 27084
rect 13219 27112 13231 27115
rect 13446 27112 13452 27124
rect 13219 27084 13452 27112
rect 13219 27081 13231 27084
rect 13173 27075 13231 27081
rect 13446 27072 13452 27084
rect 13504 27072 13510 27124
rect 15194 27072 15200 27124
rect 15252 27112 15258 27124
rect 15289 27115 15347 27121
rect 15289 27112 15301 27115
rect 15252 27084 15301 27112
rect 15252 27072 15258 27084
rect 15289 27081 15301 27084
rect 15335 27081 15347 27115
rect 17954 27112 17960 27124
rect 15289 27075 15347 27081
rect 16546 27084 17960 27112
rect 16546 27044 16574 27084
rect 17954 27072 17960 27084
rect 18012 27072 18018 27124
rect 18417 27115 18475 27121
rect 18417 27081 18429 27115
rect 18463 27081 18475 27115
rect 25314 27112 25320 27124
rect 25275 27084 25320 27112
rect 18417 27075 18475 27081
rect 10704 27016 10916 27044
rect 11532 27016 16574 27044
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 9214 26976 9220 26988
rect 8711 26948 9220 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 9214 26936 9220 26948
rect 9272 26976 9278 26988
rect 9493 26979 9551 26985
rect 9272 26948 9444 26976
rect 9272 26936 9278 26948
rect 9306 26908 9312 26920
rect 9267 26880 9312 26908
rect 9306 26868 9312 26880
rect 9364 26868 9370 26920
rect 9416 26908 9444 26948
rect 9493 26945 9505 26979
rect 9539 26976 9551 26979
rect 10318 26976 10324 26988
rect 9539 26948 10324 26976
rect 9539 26945 9551 26948
rect 9493 26939 9551 26945
rect 10318 26936 10324 26948
rect 10376 26936 10382 26988
rect 10594 26976 10600 26988
rect 10555 26948 10600 26976
rect 10594 26936 10600 26948
rect 10652 26936 10658 26988
rect 10704 26908 10732 27016
rect 10781 26979 10839 26985
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 11330 26976 11336 26988
rect 10827 26948 11336 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 11330 26936 11336 26948
rect 11388 26936 11394 26988
rect 9416 26880 10732 26908
rect 11238 26868 11244 26920
rect 11296 26908 11302 26920
rect 11532 26917 11560 27016
rect 17034 27004 17040 27056
rect 17092 27044 17098 27056
rect 17770 27044 17776 27056
rect 17092 27016 17776 27044
rect 17092 27004 17098 27016
rect 17770 27004 17776 27016
rect 17828 27044 17834 27056
rect 18432 27044 18460 27075
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 33413 27115 33471 27121
rect 27672 27084 31754 27112
rect 27672 27072 27678 27084
rect 23842 27044 23848 27056
rect 17828 27016 18460 27044
rect 23803 27016 23848 27044
rect 17828 27004 17834 27016
rect 23842 27004 23848 27016
rect 23900 27004 23906 27056
rect 25222 27044 25228 27056
rect 25070 27016 25228 27044
rect 25222 27004 25228 27016
rect 25280 27004 25286 27056
rect 27890 27004 27896 27056
rect 27948 27044 27954 27056
rect 27948 27016 31064 27044
rect 27948 27004 27954 27016
rect 31036 26988 31064 27016
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26976 13047 26979
rect 13814 26976 13820 26988
rect 13035 26948 13820 26976
rect 13035 26945 13047 26948
rect 12989 26939 13047 26945
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 15470 26976 15476 26988
rect 15431 26948 15476 26976
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15749 26979 15807 26985
rect 15749 26945 15761 26979
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 11517 26911 11575 26917
rect 11517 26908 11529 26911
rect 11296 26880 11529 26908
rect 11296 26868 11302 26880
rect 11517 26877 11529 26880
rect 11563 26877 11575 26911
rect 11517 26871 11575 26877
rect 11606 26868 11612 26920
rect 11664 26908 11670 26920
rect 11793 26911 11851 26917
rect 11793 26908 11805 26911
rect 11664 26880 11805 26908
rect 11664 26868 11670 26880
rect 11793 26877 11805 26880
rect 11839 26877 11851 26911
rect 15764 26908 15792 26939
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 15933 26979 15991 26985
rect 15933 26976 15945 26979
rect 15896 26948 15945 26976
rect 15896 26936 15902 26948
rect 15933 26945 15945 26948
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 16114 26908 16120 26920
rect 15764 26880 16120 26908
rect 11793 26871 11851 26877
rect 16114 26868 16120 26880
rect 16172 26868 16178 26920
rect 10965 26843 11023 26849
rect 10965 26809 10977 26843
rect 11011 26840 11023 26843
rect 18138 26840 18144 26852
rect 11011 26812 18144 26840
rect 11011 26809 11023 26812
rect 10965 26803 11023 26809
rect 18138 26800 18144 26812
rect 18196 26800 18202 26852
rect 8754 26772 8760 26784
rect 8715 26744 8760 26772
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 13814 26732 13820 26784
rect 13872 26772 13878 26784
rect 14642 26772 14648 26784
rect 13872 26744 14648 26772
rect 13872 26732 13878 26744
rect 14642 26732 14648 26744
rect 14700 26772 14706 26784
rect 18248 26772 18276 26939
rect 22646 26936 22652 26988
rect 22704 26976 22710 26988
rect 23569 26979 23627 26985
rect 23569 26976 23581 26979
rect 22704 26948 23581 26976
rect 22704 26936 22710 26948
rect 23569 26945 23581 26948
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 29273 26979 29331 26985
rect 29273 26976 29285 26979
rect 28316 26948 29285 26976
rect 28316 26936 28322 26948
rect 29273 26945 29285 26948
rect 29319 26945 29331 26979
rect 29273 26939 29331 26945
rect 30285 26979 30343 26985
rect 30285 26945 30297 26979
rect 30331 26976 30343 26979
rect 30926 26976 30932 26988
rect 30331 26948 30932 26976
rect 30331 26945 30343 26948
rect 30285 26939 30343 26945
rect 30926 26936 30932 26948
rect 30984 26936 30990 26988
rect 31018 26936 31024 26988
rect 31076 26976 31082 26988
rect 31113 26979 31171 26985
rect 31113 26976 31125 26979
rect 31076 26948 31125 26976
rect 31076 26936 31082 26948
rect 31113 26945 31125 26948
rect 31159 26945 31171 26979
rect 31113 26939 31171 26945
rect 31202 26936 31208 26988
rect 31260 26985 31266 26988
rect 31491 26985 31549 26991
rect 31260 26979 31295 26985
rect 31283 26945 31295 26979
rect 31260 26939 31295 26945
rect 31389 26979 31447 26985
rect 31389 26945 31401 26979
rect 31435 26945 31447 26979
rect 31491 26951 31503 26985
rect 31537 26951 31549 26985
rect 31491 26945 31549 26951
rect 31726 26976 31754 27084
rect 33413 27081 33425 27115
rect 33459 27112 33471 27115
rect 33962 27112 33968 27124
rect 33459 27084 33968 27112
rect 33459 27081 33471 27084
rect 33413 27075 33471 27081
rect 33962 27072 33968 27084
rect 34020 27072 34026 27124
rect 39945 27115 40003 27121
rect 39945 27081 39957 27115
rect 39991 27112 40003 27115
rect 40034 27112 40040 27124
rect 39991 27084 40040 27112
rect 39991 27081 40003 27084
rect 39945 27075 40003 27081
rect 40034 27072 40040 27084
rect 40092 27072 40098 27124
rect 33229 27047 33287 27053
rect 33229 27044 33241 27047
rect 32140 27016 33241 27044
rect 32140 26985 32168 27016
rect 33229 27013 33241 27016
rect 33275 27013 33287 27047
rect 33229 27007 33287 27013
rect 33336 27016 33640 27044
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 31726 26948 32137 26976
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 31389 26939 31447 26945
rect 31260 26936 31266 26939
rect 28350 26868 28356 26920
rect 28408 26908 28414 26920
rect 28810 26908 28816 26920
rect 28408 26880 28816 26908
rect 28408 26868 28414 26880
rect 28810 26868 28816 26880
rect 28868 26868 28874 26920
rect 28997 26911 29055 26917
rect 28997 26877 29009 26911
rect 29043 26908 29055 26911
rect 29086 26908 29092 26920
rect 29043 26880 29092 26908
rect 29043 26877 29055 26880
rect 28997 26871 29055 26877
rect 29086 26868 29092 26880
rect 29144 26868 29150 26920
rect 31404 26784 31432 26939
rect 31506 26908 31534 26945
rect 32125 26939 32183 26945
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26976 32367 26979
rect 32490 26976 32496 26988
rect 32355 26948 32496 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 32490 26936 32496 26948
rect 32548 26976 32554 26988
rect 33336 26976 33364 27016
rect 32548 26948 33364 26976
rect 33505 26979 33563 26985
rect 32548 26936 32554 26948
rect 33505 26945 33517 26979
rect 33551 26945 33563 26979
rect 33612 26976 33640 27016
rect 33870 27004 33876 27056
rect 33928 27044 33934 27056
rect 33928 27016 34192 27044
rect 33928 27004 33934 27016
rect 33962 26976 33968 26988
rect 33612 26948 33968 26976
rect 33505 26939 33563 26945
rect 32217 26911 32275 26917
rect 32217 26908 32229 26911
rect 31506 26880 32229 26908
rect 32217 26877 32229 26880
rect 32263 26877 32275 26911
rect 33520 26908 33548 26939
rect 33962 26936 33968 26948
rect 34020 26936 34026 26988
rect 34164 26985 34192 27016
rect 34149 26979 34207 26985
rect 34149 26945 34161 26979
rect 34195 26976 34207 26979
rect 34238 26976 34244 26988
rect 34195 26948 34244 26976
rect 34195 26945 34207 26948
rect 34149 26939 34207 26945
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 35253 26979 35311 26985
rect 35253 26945 35265 26979
rect 35299 26976 35311 26979
rect 35526 26976 35532 26988
rect 35299 26948 35532 26976
rect 35299 26945 35311 26948
rect 35253 26939 35311 26945
rect 35526 26936 35532 26948
rect 35584 26936 35590 26988
rect 39850 26976 39856 26988
rect 39811 26948 39856 26976
rect 39850 26936 39856 26948
rect 39908 26936 39914 26988
rect 34057 26911 34115 26917
rect 34057 26908 34069 26911
rect 33520 26880 34069 26908
rect 32217 26871 32275 26877
rect 34057 26877 34069 26880
rect 34103 26877 34115 26911
rect 34057 26871 34115 26877
rect 30374 26772 30380 26784
rect 14700 26744 18276 26772
rect 30335 26744 30380 26772
rect 14700 26732 14706 26744
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 30926 26772 30932 26784
rect 30887 26744 30932 26772
rect 30926 26732 30932 26744
rect 30984 26732 30990 26784
rect 31386 26732 31392 26784
rect 31444 26732 31450 26784
rect 33229 26775 33287 26781
rect 33229 26741 33241 26775
rect 33275 26772 33287 26775
rect 33318 26772 33324 26784
rect 33275 26744 33324 26772
rect 33275 26741 33287 26744
rect 33229 26735 33287 26741
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 35342 26772 35348 26784
rect 35303 26744 35348 26772
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 15470 26568 15476 26580
rect 2746 26540 15476 26568
rect 14 26392 20 26444
rect 72 26432 78 26444
rect 2746 26432 2774 26540
rect 15470 26528 15476 26540
rect 15528 26528 15534 26580
rect 22922 26568 22928 26580
rect 15764 26540 22928 26568
rect 10318 26500 10324 26512
rect 10279 26472 10324 26500
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 11609 26503 11667 26509
rect 11609 26500 11621 26503
rect 10612 26472 11621 26500
rect 72 26404 2774 26432
rect 72 26392 78 26404
rect 9306 26392 9312 26444
rect 9364 26432 9370 26444
rect 10612 26432 10640 26472
rect 11609 26469 11621 26472
rect 11655 26469 11667 26503
rect 15286 26500 15292 26512
rect 11609 26463 11667 26469
rect 13372 26472 15292 26500
rect 9364 26404 10640 26432
rect 9364 26392 9370 26404
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26364 8263 26367
rect 8478 26364 8484 26376
rect 8251 26336 8484 26364
rect 8251 26333 8263 26336
rect 8205 26327 8263 26333
rect 8478 26324 8484 26336
rect 8536 26364 8542 26376
rect 9122 26364 9128 26376
rect 8536 26336 9128 26364
rect 8536 26324 8542 26336
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 9508 26373 9536 26404
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9217 26327 9275 26333
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9950 26364 9956 26376
rect 9911 26336 9956 26364
rect 9493 26327 9551 26333
rect 9232 26296 9260 26327
rect 9950 26324 9956 26336
rect 10008 26324 10014 26376
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26364 10195 26367
rect 10502 26364 10508 26376
rect 10183 26336 10508 26364
rect 10183 26333 10195 26336
rect 10137 26327 10195 26333
rect 10502 26324 10508 26336
rect 10560 26364 10566 26376
rect 11057 26367 11115 26373
rect 10560 26336 10916 26364
rect 11057 26354 11069 26367
rect 11103 26354 11115 26367
rect 11514 26364 11520 26376
rect 10560 26324 10566 26336
rect 9858 26296 9864 26308
rect 9232 26268 9864 26296
rect 9858 26256 9864 26268
rect 9916 26256 9922 26308
rect 9968 26296 9996 26324
rect 10686 26296 10692 26308
rect 9968 26268 10692 26296
rect 10686 26256 10692 26268
rect 10744 26296 10750 26308
rect 10781 26299 10839 26305
rect 10781 26296 10793 26299
rect 10744 26268 10793 26296
rect 10744 26256 10750 26268
rect 10781 26265 10793 26268
rect 10827 26265 10839 26299
rect 10888 26296 10916 26336
rect 10965 26299 11023 26305
rect 11054 26302 11060 26354
rect 11112 26302 11118 26354
rect 11475 26336 11520 26364
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 13372 26373 13400 26472
rect 15286 26460 15292 26472
rect 15344 26460 15350 26512
rect 15764 26500 15792 26540
rect 22922 26528 22928 26540
rect 22980 26528 22986 26580
rect 24302 26528 24308 26580
rect 24360 26568 24366 26580
rect 24581 26571 24639 26577
rect 24581 26568 24593 26571
rect 24360 26540 24593 26568
rect 24360 26528 24366 26540
rect 24581 26537 24593 26540
rect 24627 26537 24639 26571
rect 25222 26568 25228 26580
rect 25183 26540 25228 26568
rect 24581 26531 24639 26537
rect 15396 26472 15792 26500
rect 14093 26435 14151 26441
rect 14093 26401 14105 26435
rect 14139 26432 14151 26435
rect 15396 26432 15424 26472
rect 15838 26460 15844 26512
rect 15896 26500 15902 26512
rect 16393 26503 16451 26509
rect 16393 26500 16405 26503
rect 15896 26472 16405 26500
rect 15896 26460 15902 26472
rect 16393 26469 16405 26472
rect 16439 26469 16451 26503
rect 16393 26463 16451 26469
rect 14139 26404 15424 26432
rect 14139 26401 14151 26404
rect 14093 26395 14151 26401
rect 15470 26392 15476 26444
rect 15528 26432 15534 26444
rect 15528 26404 15573 26432
rect 15528 26392 15534 26404
rect 11701 26367 11759 26373
rect 11701 26333 11713 26367
rect 11747 26333 11759 26367
rect 11701 26327 11759 26333
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 10965 26296 10977 26299
rect 10888 26268 10977 26296
rect 10781 26259 10839 26265
rect 10965 26265 10977 26268
rect 11011 26265 11023 26299
rect 10965 26259 11023 26265
rect 11606 26256 11612 26308
rect 11664 26296 11670 26308
rect 11716 26296 11744 26327
rect 15746 26324 15752 26376
rect 15804 26364 15810 26376
rect 16390 26364 16396 26376
rect 15804 26336 16396 26364
rect 15804 26324 15810 26336
rect 16390 26324 16396 26336
rect 16448 26324 16454 26376
rect 16666 26364 16672 26376
rect 16627 26336 16672 26364
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 24394 26364 24400 26376
rect 24355 26336 24400 26364
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24596 26364 24624 26531
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 31662 26528 31668 26580
rect 31720 26568 31726 26580
rect 31720 26540 32628 26568
rect 31720 26528 31726 26540
rect 26973 26503 27031 26509
rect 26973 26469 26985 26503
rect 27019 26469 27031 26503
rect 26973 26463 27031 26469
rect 26510 26432 26516 26444
rect 26471 26404 26516 26432
rect 26510 26392 26516 26404
rect 26568 26392 26574 26444
rect 25038 26364 25044 26376
rect 24596 26336 25044 26364
rect 25038 26324 25044 26336
rect 25096 26364 25102 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 25096 26336 25145 26364
rect 25096 26324 25102 26336
rect 25133 26333 25145 26336
rect 25179 26333 25191 26367
rect 26602 26364 26608 26376
rect 26563 26336 26608 26364
rect 25133 26327 25191 26333
rect 26602 26324 26608 26336
rect 26660 26324 26666 26376
rect 26988 26364 27016 26463
rect 27982 26392 27988 26444
rect 28040 26432 28046 26444
rect 32398 26432 32404 26444
rect 28040 26404 28396 26432
rect 28040 26392 28046 26404
rect 27433 26367 27491 26373
rect 27433 26364 27445 26367
rect 26988 26336 27445 26364
rect 27433 26333 27445 26336
rect 27479 26333 27491 26367
rect 27614 26364 27620 26376
rect 27575 26336 27620 26364
rect 27433 26327 27491 26333
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 28074 26364 28080 26376
rect 28035 26336 28080 26364
rect 28074 26324 28080 26336
rect 28132 26324 28138 26376
rect 28258 26373 28264 26376
rect 28225 26367 28264 26373
rect 28225 26333 28237 26367
rect 28225 26327 28264 26333
rect 28258 26324 28264 26327
rect 28316 26324 28322 26376
rect 28368 26364 28396 26404
rect 30668 26404 32404 26432
rect 30668 26373 30696 26404
rect 32398 26392 32404 26404
rect 32456 26392 32462 26444
rect 32600 26432 32628 26540
rect 32674 26528 32680 26580
rect 32732 26568 32738 26580
rect 39850 26568 39856 26580
rect 32732 26540 39856 26568
rect 32732 26528 32738 26540
rect 35452 26432 35480 26540
rect 39850 26528 39856 26540
rect 39908 26528 39914 26580
rect 35529 26435 35587 26441
rect 35529 26432 35541 26435
rect 32600 26404 33548 26432
rect 35452 26404 35541 26432
rect 28542 26367 28600 26373
rect 28542 26364 28554 26367
rect 28368 26336 28554 26364
rect 28542 26333 28554 26336
rect 28588 26333 28600 26367
rect 30653 26367 30711 26373
rect 30653 26364 30665 26367
rect 28542 26327 28600 26333
rect 30392 26336 30665 26364
rect 11664 26268 11744 26296
rect 13449 26299 13507 26305
rect 11664 26256 11670 26268
rect 13449 26265 13461 26299
rect 13495 26296 13507 26299
rect 14277 26299 14335 26305
rect 14277 26296 14289 26299
rect 13495 26268 14289 26296
rect 13495 26265 13507 26268
rect 13449 26259 13507 26265
rect 14277 26265 14289 26268
rect 14323 26265 14335 26299
rect 24412 26296 24440 26324
rect 26694 26296 26700 26308
rect 24412 26268 26700 26296
rect 14277 26259 14335 26265
rect 26694 26256 26700 26268
rect 26752 26296 26758 26308
rect 27154 26296 27160 26308
rect 26752 26268 27160 26296
rect 26752 26256 26758 26268
rect 27154 26256 27160 26268
rect 27212 26256 27218 26308
rect 27246 26256 27252 26308
rect 27304 26296 27310 26308
rect 27890 26296 27896 26308
rect 27304 26268 27896 26296
rect 27304 26256 27310 26268
rect 27890 26256 27896 26268
rect 27948 26296 27954 26308
rect 28353 26299 28411 26305
rect 28353 26296 28365 26299
rect 27948 26268 28365 26296
rect 27948 26256 27954 26268
rect 28353 26265 28365 26268
rect 28399 26265 28411 26299
rect 28353 26259 28411 26265
rect 28442 26256 28448 26308
rect 28500 26296 28506 26308
rect 28500 26268 28545 26296
rect 28500 26256 28506 26268
rect 7926 26188 7932 26240
rect 7984 26228 7990 26240
rect 8205 26231 8263 26237
rect 8205 26228 8217 26231
rect 7984 26200 8217 26228
rect 7984 26188 7990 26200
rect 8205 26197 8217 26200
rect 8251 26197 8263 26231
rect 8205 26191 8263 26197
rect 8294 26188 8300 26240
rect 8352 26228 8358 26240
rect 9033 26231 9091 26237
rect 9033 26228 9045 26231
rect 8352 26200 9045 26228
rect 8352 26188 8358 26200
rect 9033 26197 9045 26200
rect 9079 26197 9091 26231
rect 9033 26191 9091 26197
rect 9401 26231 9459 26237
rect 9401 26197 9413 26231
rect 9447 26228 9459 26231
rect 9674 26228 9680 26240
rect 9447 26200 9680 26228
rect 9447 26197 9459 26200
rect 9401 26191 9459 26197
rect 9674 26188 9680 26200
rect 9732 26188 9738 26240
rect 11057 26231 11115 26237
rect 11057 26197 11069 26231
rect 11103 26228 11115 26231
rect 11422 26228 11428 26240
rect 11103 26200 11428 26228
rect 11103 26197 11115 26200
rect 11057 26191 11115 26197
rect 11422 26188 11428 26200
rect 11480 26188 11486 26240
rect 16577 26231 16635 26237
rect 16577 26197 16589 26231
rect 16623 26228 16635 26231
rect 17034 26228 17040 26240
rect 16623 26200 17040 26228
rect 16623 26197 16635 26200
rect 16577 26191 16635 26197
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 26970 26188 26976 26240
rect 27028 26228 27034 26240
rect 27525 26231 27583 26237
rect 27525 26228 27537 26231
rect 27028 26200 27537 26228
rect 27028 26188 27034 26200
rect 27525 26197 27537 26200
rect 27571 26197 27583 26231
rect 28718 26228 28724 26240
rect 28679 26200 28724 26228
rect 27525 26191 27583 26197
rect 28718 26188 28724 26200
rect 28776 26188 28782 26240
rect 28902 26188 28908 26240
rect 28960 26228 28966 26240
rect 30392 26228 30420 26336
rect 30653 26333 30665 26336
rect 30699 26333 30711 26367
rect 30653 26327 30711 26333
rect 33045 26367 33103 26373
rect 33045 26333 33057 26367
rect 33091 26333 33103 26367
rect 33045 26327 33103 26333
rect 33137 26367 33195 26373
rect 33137 26333 33149 26367
rect 33183 26333 33195 26367
rect 33318 26364 33324 26376
rect 33279 26336 33324 26364
rect 33137 26327 33195 26333
rect 30926 26296 30932 26308
rect 30887 26268 30932 26296
rect 30926 26256 30932 26268
rect 30984 26256 30990 26308
rect 31938 26256 31944 26308
rect 31996 26256 32002 26308
rect 33060 26296 33088 26327
rect 32232 26268 33088 26296
rect 28960 26200 30420 26228
rect 28960 26188 28966 26200
rect 31018 26188 31024 26240
rect 31076 26228 31082 26240
rect 32232 26228 32260 26268
rect 31076 26200 32260 26228
rect 32401 26231 32459 26237
rect 31076 26188 31082 26200
rect 32401 26197 32413 26231
rect 32447 26228 32459 26231
rect 32490 26228 32496 26240
rect 32447 26200 32496 26228
rect 32447 26197 32459 26200
rect 32401 26191 32459 26197
rect 32490 26188 32496 26200
rect 32548 26188 32554 26240
rect 32858 26228 32864 26240
rect 32819 26200 32864 26228
rect 32858 26188 32864 26200
rect 32916 26188 32922 26240
rect 33152 26228 33180 26327
rect 33318 26324 33324 26336
rect 33376 26324 33382 26376
rect 33413 26367 33471 26373
rect 33413 26333 33425 26367
rect 33459 26333 33471 26367
rect 33520 26364 33548 26404
rect 35529 26401 35541 26404
rect 35575 26401 35587 26435
rect 35529 26395 35587 26401
rect 33873 26367 33931 26373
rect 33873 26364 33885 26367
rect 33520 26336 33885 26364
rect 33413 26327 33471 26333
rect 33873 26333 33885 26336
rect 33919 26333 33931 26367
rect 35342 26364 35348 26376
rect 35303 26336 35348 26364
rect 33873 26327 33931 26333
rect 33428 26296 33456 26327
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 39868 26364 39896 26528
rect 45005 26367 45063 26373
rect 45005 26364 45017 26367
rect 39868 26336 45017 26364
rect 45005 26333 45017 26336
rect 45051 26333 45063 26367
rect 47670 26364 47676 26376
rect 47631 26336 47676 26364
rect 45005 26327 45063 26333
rect 47670 26324 47676 26336
rect 47728 26324 47734 26376
rect 33594 26296 33600 26308
rect 33428 26268 33600 26296
rect 33594 26256 33600 26268
rect 33652 26256 33658 26308
rect 33778 26256 33784 26308
rect 33836 26296 33842 26308
rect 33965 26299 34023 26305
rect 33965 26296 33977 26299
rect 33836 26268 33977 26296
rect 33836 26256 33842 26268
rect 33965 26265 33977 26268
rect 34011 26265 34023 26299
rect 33965 26259 34023 26265
rect 34238 26228 34244 26240
rect 33152 26200 34244 26228
rect 34238 26188 34244 26200
rect 34296 26188 34302 26240
rect 45094 26228 45100 26240
rect 45055 26200 45100 26228
rect 45094 26188 45100 26200
rect 45152 26188 45158 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 9858 25984 9864 26036
rect 9916 26024 9922 26036
rect 10781 26027 10839 26033
rect 10781 26024 10793 26027
rect 9916 25996 10793 26024
rect 9916 25984 9922 25996
rect 10781 25993 10793 25996
rect 10827 25993 10839 26027
rect 16114 26024 16120 26036
rect 16075 25996 16120 26024
rect 10781 25987 10839 25993
rect 16114 25984 16120 25996
rect 16172 25984 16178 26036
rect 16390 25984 16396 26036
rect 16448 26024 16454 26036
rect 16945 26027 17003 26033
rect 16945 26024 16957 26027
rect 16448 25996 16957 26024
rect 16448 25984 16454 25996
rect 16945 25993 16957 25996
rect 16991 25993 17003 26027
rect 16945 25987 17003 25993
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 23477 26027 23535 26033
rect 23477 26024 23489 26027
rect 18656 25996 23489 26024
rect 18656 25984 18662 25996
rect 23477 25993 23489 25996
rect 23523 25993 23535 26027
rect 28902 26024 28908 26036
rect 23477 25987 23535 25993
rect 24688 25996 28908 26024
rect 8205 25959 8263 25965
rect 8205 25925 8217 25959
rect 8251 25956 8263 25959
rect 8294 25956 8300 25968
rect 8251 25928 8300 25956
rect 8251 25925 8263 25928
rect 8205 25919 8263 25925
rect 8294 25916 8300 25928
rect 8352 25916 8358 25968
rect 8754 25916 8760 25968
rect 8812 25916 8818 25968
rect 10597 25959 10655 25965
rect 10597 25925 10609 25959
rect 10643 25956 10655 25959
rect 10686 25956 10692 25968
rect 10643 25928 10692 25956
rect 10643 25925 10655 25928
rect 10597 25919 10655 25925
rect 10686 25916 10692 25928
rect 10744 25956 10750 25968
rect 11514 25956 11520 25968
rect 10744 25928 11520 25956
rect 10744 25916 10750 25928
rect 11514 25916 11520 25928
rect 11572 25916 11578 25968
rect 15746 25956 15752 25968
rect 15707 25928 15752 25956
rect 15746 25916 15752 25928
rect 15804 25916 15810 25968
rect 15965 25959 16023 25965
rect 15965 25925 15977 25959
rect 16011 25956 16023 25959
rect 16758 25956 16764 25968
rect 16011 25928 16574 25956
rect 16719 25928 16764 25956
rect 16011 25925 16023 25928
rect 15965 25919 16023 25925
rect 7926 25888 7932 25900
rect 7887 25860 7932 25888
rect 7926 25848 7932 25860
rect 7984 25848 7990 25900
rect 11330 25848 11336 25900
rect 11388 25888 11394 25900
rect 11698 25888 11704 25900
rect 11388 25860 11704 25888
rect 11388 25848 11394 25860
rect 11698 25848 11704 25860
rect 11756 25848 11762 25900
rect 14642 25888 14648 25900
rect 14603 25860 14648 25888
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 16546 25888 16574 25928
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 17313 25959 17371 25965
rect 16868 25928 17172 25956
rect 16666 25888 16672 25900
rect 16546 25860 16672 25888
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 15378 25780 15384 25832
rect 15436 25820 15442 25832
rect 16868 25820 16896 25928
rect 17034 25888 17040 25900
rect 16995 25860 17040 25888
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17144 25897 17172 25928
rect 17313 25925 17325 25959
rect 17359 25956 17371 25959
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 17359 25928 23305 25956
rect 17359 25925 17371 25928
rect 17313 25919 17371 25925
rect 23293 25925 23305 25928
rect 23339 25925 23351 25959
rect 23293 25919 23351 25925
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17402 25888 17408 25900
rect 17175 25860 17408 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 17770 25888 17776 25900
rect 17731 25860 17776 25888
rect 17770 25848 17776 25860
rect 17828 25888 17834 25900
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 17828 25860 19073 25888
rect 17828 25848 17834 25860
rect 19061 25857 19073 25860
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19242 25848 19248 25900
rect 19300 25888 19306 25900
rect 19889 25891 19947 25897
rect 19889 25888 19901 25891
rect 19300 25860 19901 25888
rect 19300 25848 19306 25860
rect 19889 25857 19901 25860
rect 19935 25888 19947 25891
rect 20990 25888 20996 25900
rect 19935 25860 20996 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 21542 25848 21548 25900
rect 21600 25888 21606 25900
rect 22051 25891 22109 25897
rect 22051 25888 22063 25891
rect 21600 25860 22063 25888
rect 21600 25848 21606 25860
rect 22051 25857 22063 25860
rect 22097 25857 22109 25891
rect 22051 25851 22109 25857
rect 22186 25891 22244 25897
rect 22186 25857 22198 25891
rect 22232 25857 22244 25891
rect 22186 25851 22244 25857
rect 15436 25792 16896 25820
rect 15436 25780 15442 25792
rect 17494 25780 17500 25832
rect 17552 25820 17558 25832
rect 19978 25820 19984 25832
rect 17552 25792 19748 25820
rect 19939 25792 19984 25820
rect 17552 25780 17558 25792
rect 9674 25752 9680 25764
rect 9587 25724 9680 25752
rect 9674 25712 9680 25724
rect 9732 25752 9738 25764
rect 10229 25755 10287 25761
rect 10229 25752 10241 25755
rect 9732 25724 10241 25752
rect 9732 25712 9738 25724
rect 10229 25721 10241 25724
rect 10275 25752 10287 25755
rect 10778 25752 10784 25764
rect 10275 25724 10784 25752
rect 10275 25721 10287 25724
rect 10229 25715 10287 25721
rect 10778 25712 10784 25724
rect 10836 25712 10842 25764
rect 17034 25752 17040 25764
rect 15948 25724 17040 25752
rect 10502 25644 10508 25696
rect 10560 25684 10566 25696
rect 10597 25687 10655 25693
rect 10597 25684 10609 25687
rect 10560 25656 10609 25684
rect 10560 25644 10566 25656
rect 10597 25653 10609 25656
rect 10643 25684 10655 25687
rect 11517 25687 11575 25693
rect 11517 25684 11529 25687
rect 10643 25656 11529 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 11517 25653 11529 25656
rect 11563 25684 11575 25687
rect 11606 25684 11612 25696
rect 11563 25656 11612 25684
rect 11563 25653 11575 25656
rect 11517 25647 11575 25653
rect 11606 25644 11612 25656
rect 11664 25644 11670 25696
rect 14829 25687 14887 25693
rect 14829 25653 14841 25687
rect 14875 25684 14887 25687
rect 15010 25684 15016 25696
rect 14875 25656 15016 25684
rect 14875 25653 14887 25656
rect 14829 25647 14887 25653
rect 15010 25644 15016 25656
rect 15068 25644 15074 25696
rect 15948 25693 15976 25724
rect 17034 25712 17040 25724
rect 17092 25712 17098 25764
rect 17865 25755 17923 25761
rect 17865 25752 17877 25755
rect 17236 25724 17877 25752
rect 15933 25687 15991 25693
rect 15933 25653 15945 25687
rect 15979 25653 15991 25687
rect 15933 25647 15991 25653
rect 16390 25644 16396 25696
rect 16448 25684 16454 25696
rect 17236 25684 17264 25724
rect 17865 25721 17877 25724
rect 17911 25721 17923 25755
rect 17865 25715 17923 25721
rect 19153 25755 19211 25761
rect 19153 25721 19165 25755
rect 19199 25752 19211 25755
rect 19610 25752 19616 25764
rect 19199 25724 19616 25752
rect 19199 25721 19211 25724
rect 19153 25715 19211 25721
rect 19610 25712 19616 25724
rect 19668 25712 19674 25764
rect 19720 25752 19748 25792
rect 19978 25780 19984 25792
rect 20036 25780 20042 25832
rect 22204 25820 22232 25851
rect 22278 25848 22284 25900
rect 22336 25888 22342 25900
rect 22465 25891 22523 25897
rect 22336 25860 22381 25888
rect 22336 25848 22342 25860
rect 22465 25857 22477 25891
rect 22511 25888 22523 25891
rect 22554 25888 22560 25900
rect 22511 25860 22560 25888
rect 22511 25857 22523 25860
rect 22465 25851 22523 25857
rect 22554 25848 22560 25860
rect 22612 25848 22618 25900
rect 22922 25888 22928 25900
rect 22883 25860 22928 25888
rect 22922 25848 22928 25860
rect 22980 25848 22986 25900
rect 23109 25891 23167 25897
rect 23109 25857 23121 25891
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 23124 25820 23152 25851
rect 23198 25848 23204 25900
rect 23256 25888 23262 25900
rect 24688 25897 24716 25996
rect 25406 25916 25412 25968
rect 25464 25916 25470 25968
rect 26602 25916 26608 25968
rect 26660 25956 26666 25968
rect 28442 25956 28448 25968
rect 26660 25928 27108 25956
rect 26660 25916 26666 25928
rect 24673 25891 24731 25897
rect 23256 25860 23301 25888
rect 23256 25848 23262 25860
rect 24673 25857 24685 25891
rect 24719 25857 24731 25891
rect 26970 25888 26976 25900
rect 26931 25860 26976 25888
rect 24673 25851 24731 25857
rect 26970 25848 26976 25860
rect 27028 25848 27034 25900
rect 27080 25897 27108 25928
rect 27356 25928 28448 25956
rect 27066 25891 27124 25897
rect 27066 25857 27078 25891
rect 27112 25857 27124 25891
rect 27246 25888 27252 25900
rect 27207 25860 27252 25888
rect 27066 25851 27124 25857
rect 27246 25848 27252 25860
rect 27304 25848 27310 25900
rect 27356 25897 27384 25928
rect 28442 25916 28448 25928
rect 28500 25916 28506 25968
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 27430 25848 27436 25900
rect 27488 25897 27494 25900
rect 28552 25897 28580 25996
rect 28902 25984 28908 25996
rect 28960 25984 28966 26036
rect 29086 25984 29092 26036
rect 29144 26024 29150 26036
rect 30285 26027 30343 26033
rect 30285 26024 30297 26027
rect 29144 25996 30297 26024
rect 29144 25984 29150 25996
rect 30285 25993 30297 25996
rect 30331 25993 30343 26027
rect 30285 25987 30343 25993
rect 31481 26027 31539 26033
rect 31481 25993 31493 26027
rect 31527 26024 31539 26027
rect 31938 26024 31944 26036
rect 31527 25996 31944 26024
rect 31527 25993 31539 25996
rect 31481 25987 31539 25993
rect 31938 25984 31944 25996
rect 31996 25984 32002 26036
rect 34238 26024 34244 26036
rect 34199 25996 34244 26024
rect 34238 25984 34244 25996
rect 34296 25984 34302 26036
rect 28718 25916 28724 25968
rect 28776 25956 28782 25968
rect 28813 25959 28871 25965
rect 28813 25956 28825 25959
rect 28776 25928 28825 25956
rect 28776 25916 28782 25928
rect 28813 25925 28825 25928
rect 28859 25925 28871 25959
rect 30374 25956 30380 25968
rect 30038 25928 30380 25956
rect 28813 25919 28871 25925
rect 30374 25916 30380 25928
rect 30432 25916 30438 25968
rect 32769 25959 32827 25965
rect 32769 25925 32781 25959
rect 32815 25956 32827 25959
rect 32858 25956 32864 25968
rect 32815 25928 32864 25956
rect 32815 25925 32827 25928
rect 32769 25919 32827 25925
rect 32858 25916 32864 25928
rect 32916 25916 32922 25968
rect 33778 25916 33784 25968
rect 33836 25916 33842 25968
rect 35434 25916 35440 25968
rect 35492 25956 35498 25968
rect 35529 25959 35587 25965
rect 35529 25956 35541 25959
rect 35492 25928 35541 25956
rect 35492 25916 35498 25928
rect 35529 25925 35541 25928
rect 35575 25925 35587 25959
rect 35529 25919 35587 25925
rect 45094 25916 45100 25968
rect 45152 25956 45158 25968
rect 45281 25959 45339 25965
rect 45281 25956 45293 25959
rect 45152 25928 45293 25956
rect 45152 25916 45158 25928
rect 45281 25925 45293 25928
rect 45327 25925 45339 25959
rect 45281 25919 45339 25925
rect 27488 25888 27496 25897
rect 28537 25891 28595 25897
rect 27488 25860 27533 25888
rect 27488 25851 27496 25860
rect 28537 25857 28549 25891
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25888 31447 25891
rect 31662 25888 31668 25900
rect 31435 25860 31668 25888
rect 31435 25857 31447 25860
rect 31389 25851 31447 25857
rect 27488 25848 27494 25851
rect 31662 25848 31668 25860
rect 31720 25848 31726 25900
rect 32398 25848 32404 25900
rect 32456 25888 32462 25900
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 32456 25860 32505 25888
rect 32456 25848 32462 25860
rect 32493 25857 32505 25860
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 35253 25891 35311 25897
rect 35253 25888 35265 25891
rect 34848 25860 35265 25888
rect 34848 25848 34854 25860
rect 35253 25857 35265 25860
rect 35299 25888 35311 25891
rect 35342 25888 35348 25900
rect 35299 25860 35348 25888
rect 35299 25857 35311 25860
rect 35253 25851 35311 25857
rect 35342 25848 35348 25860
rect 35400 25888 35406 25900
rect 36173 25891 36231 25897
rect 36173 25888 36185 25891
rect 35400 25860 36185 25888
rect 35400 25848 35406 25860
rect 36173 25857 36185 25860
rect 36219 25857 36231 25891
rect 36173 25851 36231 25857
rect 24026 25820 24032 25832
rect 22204 25792 22324 25820
rect 23124 25792 24032 25820
rect 21821 25755 21879 25761
rect 21821 25752 21833 25755
rect 19720 25724 21833 25752
rect 21821 25721 21833 25724
rect 21867 25721 21879 25755
rect 21821 25715 21879 25721
rect 16448 25656 17264 25684
rect 16448 25644 16454 25656
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 19242 25684 19248 25696
rect 17460 25656 19248 25684
rect 17460 25644 17466 25656
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 20257 25687 20315 25693
rect 20257 25684 20269 25687
rect 19576 25656 20269 25684
rect 19576 25644 19582 25656
rect 20257 25653 20269 25656
rect 20303 25653 20315 25687
rect 22296 25684 22324 25792
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 24949 25823 25007 25829
rect 24949 25789 24961 25823
rect 24995 25820 25007 25823
rect 45094 25820 45100 25832
rect 24995 25792 26740 25820
rect 45055 25792 45100 25820
rect 24995 25789 25007 25792
rect 24949 25783 25007 25789
rect 26421 25755 26479 25761
rect 26421 25721 26433 25755
rect 26467 25752 26479 25755
rect 26602 25752 26608 25764
rect 26467 25724 26608 25752
rect 26467 25721 26479 25724
rect 26421 25715 26479 25721
rect 26602 25712 26608 25724
rect 26660 25712 26666 25764
rect 26712 25752 26740 25792
rect 45094 25780 45100 25792
rect 45152 25780 45158 25832
rect 46842 25820 46848 25832
rect 46803 25792 46848 25820
rect 46842 25780 46848 25792
rect 46900 25780 46906 25832
rect 27617 25755 27675 25761
rect 27617 25752 27629 25755
rect 26712 25724 27629 25752
rect 27617 25721 27629 25724
rect 27663 25721 27675 25755
rect 27617 25715 27675 25721
rect 27338 25684 27344 25696
rect 22296 25656 27344 25684
rect 20257 25647 20315 25653
rect 27338 25644 27344 25656
rect 27396 25644 27402 25696
rect 35894 25644 35900 25696
rect 35952 25684 35958 25696
rect 36265 25687 36323 25693
rect 36265 25684 36277 25687
rect 35952 25656 36277 25684
rect 35952 25644 35958 25656
rect 36265 25653 36277 25656
rect 36311 25653 36323 25687
rect 47762 25684 47768 25696
rect 47723 25656 47768 25684
rect 36265 25647 36323 25653
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 10502 25440 10508 25492
rect 10560 25440 10566 25492
rect 14277 25483 14335 25489
rect 14277 25449 14289 25483
rect 14323 25480 14335 25483
rect 14642 25480 14648 25492
rect 14323 25452 14648 25480
rect 14323 25449 14335 25452
rect 14277 25443 14335 25449
rect 14642 25440 14648 25452
rect 14700 25440 14706 25492
rect 16482 25440 16488 25492
rect 16540 25480 16546 25492
rect 16761 25483 16819 25489
rect 16761 25480 16773 25483
rect 16540 25452 16773 25480
rect 16540 25440 16546 25452
rect 16761 25449 16773 25452
rect 16807 25449 16819 25483
rect 16761 25443 16819 25449
rect 19978 25440 19984 25492
rect 20036 25480 20042 25492
rect 22002 25480 22008 25492
rect 20036 25452 22008 25480
rect 20036 25440 20042 25452
rect 22002 25440 22008 25452
rect 22060 25440 22066 25492
rect 22649 25483 22707 25489
rect 22649 25449 22661 25483
rect 22695 25480 22707 25483
rect 24026 25480 24032 25492
rect 22695 25452 24032 25480
rect 22695 25449 22707 25452
rect 22649 25443 22707 25449
rect 24026 25440 24032 25452
rect 24084 25440 24090 25492
rect 25133 25483 25191 25489
rect 25133 25449 25145 25483
rect 25179 25480 25191 25483
rect 25406 25480 25412 25492
rect 25179 25452 25412 25480
rect 25179 25449 25191 25452
rect 25133 25443 25191 25449
rect 25406 25440 25412 25452
rect 25464 25440 25470 25492
rect 26786 25440 26792 25492
rect 26844 25480 26850 25492
rect 29917 25483 29975 25489
rect 29917 25480 29929 25483
rect 26844 25452 29929 25480
rect 26844 25440 26850 25452
rect 29917 25449 29929 25452
rect 29963 25449 29975 25483
rect 33594 25480 33600 25492
rect 33555 25452 33600 25480
rect 29917 25443 29975 25449
rect 33594 25440 33600 25452
rect 33652 25440 33658 25492
rect 10520 25412 10548 25440
rect 20990 25412 20996 25424
rect 10520 25384 10732 25412
rect 20903 25384 20996 25412
rect 10410 25344 10416 25356
rect 10371 25316 10416 25344
rect 10410 25304 10416 25316
rect 10468 25304 10474 25356
rect 10505 25347 10563 25353
rect 10505 25313 10517 25347
rect 10551 25344 10563 25347
rect 10594 25344 10600 25356
rect 10551 25316 10600 25344
rect 10551 25313 10563 25316
rect 10505 25307 10563 25313
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 10612 25208 10640 25304
rect 10704 25276 10732 25384
rect 20990 25372 20996 25384
rect 21048 25412 21054 25424
rect 22554 25412 22560 25424
rect 21048 25384 22560 25412
rect 21048 25372 21054 25384
rect 22554 25372 22560 25384
rect 22612 25372 22618 25424
rect 22833 25415 22891 25421
rect 22833 25381 22845 25415
rect 22879 25381 22891 25415
rect 22833 25375 22891 25381
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25344 10931 25347
rect 11238 25344 11244 25356
rect 10919 25316 11244 25344
rect 10919 25313 10931 25316
rect 10873 25307 10931 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11422 25344 11428 25356
rect 11383 25316 11428 25344
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 15010 25344 15016 25356
rect 14971 25316 15016 25344
rect 15010 25304 15016 25316
rect 15068 25304 15074 25356
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 17494 25344 17500 25356
rect 16724 25316 17500 25344
rect 16724 25304 16730 25316
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 18046 25344 18052 25356
rect 17819 25316 18052 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 18046 25304 18052 25316
rect 18104 25304 18110 25356
rect 19518 25344 19524 25356
rect 19479 25316 19524 25344
rect 19518 25304 19524 25316
rect 19576 25304 19582 25356
rect 22278 25344 22284 25356
rect 21836 25316 22284 25344
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 10704 25248 10793 25276
rect 10781 25245 10793 25248
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25245 11575 25279
rect 12434 25276 12440 25288
rect 12395 25248 12440 25276
rect 11517 25239 11575 25245
rect 11532 25208 11560 25239
rect 12434 25236 12440 25248
rect 12492 25236 12498 25288
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 12676 25248 14105 25276
rect 12676 25236 12682 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 16390 25236 16396 25288
rect 16448 25236 16454 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17402 25276 17408 25288
rect 17092 25248 17408 25276
rect 17092 25236 17098 25248
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 17862 25236 17868 25288
rect 17920 25276 17926 25288
rect 21836 25285 21864 25316
rect 22278 25304 22284 25316
rect 22336 25344 22342 25356
rect 22848 25344 22876 25375
rect 27246 25372 27252 25424
rect 27304 25412 27310 25424
rect 27430 25412 27436 25424
rect 27304 25384 27436 25412
rect 27304 25372 27310 25384
rect 27430 25372 27436 25384
rect 27488 25372 27494 25424
rect 22336 25316 22876 25344
rect 22336 25304 22342 25316
rect 28442 25304 28448 25356
rect 28500 25344 28506 25356
rect 29549 25347 29607 25353
rect 29549 25344 29561 25347
rect 28500 25316 29561 25344
rect 28500 25304 28506 25316
rect 29549 25313 29561 25316
rect 29595 25344 29607 25347
rect 31570 25344 31576 25356
rect 29595 25316 31576 25344
rect 29595 25313 29607 25316
rect 29549 25307 29607 25313
rect 31570 25304 31576 25316
rect 31628 25344 31634 25356
rect 33229 25347 33287 25353
rect 33229 25344 33241 25347
rect 31628 25316 33241 25344
rect 31628 25304 31634 25316
rect 33229 25313 33241 25316
rect 33275 25313 33287 25347
rect 35894 25344 35900 25356
rect 35855 25316 35900 25344
rect 33229 25307 33287 25313
rect 35894 25304 35900 25316
rect 35952 25304 35958 25356
rect 46293 25347 46351 25353
rect 46293 25313 46305 25347
rect 46339 25344 46351 25347
rect 47670 25344 47676 25356
rect 46339 25316 47676 25344
rect 46339 25313 46351 25316
rect 46293 25307 46351 25313
rect 47670 25304 47676 25316
rect 47728 25304 47734 25356
rect 18509 25279 18567 25285
rect 18509 25276 18521 25279
rect 17920 25248 18521 25276
rect 17920 25236 17926 25248
rect 18509 25245 18521 25248
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 21729 25239 21787 25245
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25245 21879 25279
rect 25038 25276 25044 25288
rect 24999 25248 25044 25276
rect 21821 25239 21879 25245
rect 13354 25208 13360 25220
rect 10612 25180 13360 25208
rect 13354 25168 13360 25180
rect 13412 25168 13418 25220
rect 15286 25208 15292 25220
rect 15247 25180 15292 25208
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 19260 25208 19288 25239
rect 19426 25208 19432 25220
rect 19260 25180 19432 25208
rect 19426 25168 19432 25180
rect 19484 25168 19490 25220
rect 19610 25168 19616 25220
rect 19668 25208 19674 25220
rect 21744 25208 21772 25239
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25276 29791 25279
rect 29914 25276 29920 25288
rect 29779 25248 29920 25276
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 29914 25236 29920 25248
rect 29972 25236 29978 25288
rect 33410 25276 33416 25288
rect 33371 25248 33416 25276
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 34790 25236 34796 25288
rect 34848 25276 34854 25288
rect 34885 25279 34943 25285
rect 34885 25276 34897 25279
rect 34848 25248 34897 25276
rect 34848 25236 34854 25248
rect 34885 25245 34897 25248
rect 34931 25245 34943 25279
rect 34885 25239 34943 25245
rect 35713 25279 35771 25285
rect 35713 25245 35725 25279
rect 35759 25245 35771 25279
rect 35713 25239 35771 25245
rect 22370 25208 22376 25220
rect 19668 25180 20010 25208
rect 21744 25180 22376 25208
rect 19668 25168 19674 25180
rect 22370 25168 22376 25180
rect 22428 25168 22434 25220
rect 22465 25211 22523 25217
rect 22465 25177 22477 25211
rect 22511 25208 22523 25211
rect 22922 25208 22928 25220
rect 22511 25180 22928 25208
rect 22511 25177 22523 25180
rect 22465 25171 22523 25177
rect 22922 25168 22928 25180
rect 22980 25168 22986 25220
rect 32122 25168 32128 25220
rect 32180 25208 32186 25220
rect 35728 25208 35756 25239
rect 32180 25180 35756 25208
rect 37553 25211 37611 25217
rect 32180 25168 32186 25180
rect 37553 25177 37565 25211
rect 37599 25208 37611 25211
rect 45554 25208 45560 25220
rect 37599 25180 45560 25208
rect 37599 25177 37611 25180
rect 37553 25171 37611 25177
rect 45554 25168 45560 25180
rect 45612 25168 45618 25220
rect 46477 25211 46535 25217
rect 46477 25177 46489 25211
rect 46523 25208 46535 25211
rect 46934 25208 46940 25220
rect 46523 25180 46940 25208
rect 46523 25177 46535 25180
rect 46477 25171 46535 25177
rect 46934 25168 46940 25180
rect 46992 25168 46998 25220
rect 48130 25208 48136 25220
rect 48091 25180 48136 25208
rect 48130 25168 48136 25180
rect 48188 25168 48194 25220
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2038 25140 2044 25152
rect 1995 25112 2044 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 10042 25100 10048 25152
rect 10100 25140 10106 25152
rect 10229 25143 10287 25149
rect 10229 25140 10241 25143
rect 10100 25112 10241 25140
rect 10100 25100 10106 25112
rect 10229 25109 10241 25112
rect 10275 25109 10287 25143
rect 10229 25103 10287 25109
rect 10689 25143 10747 25149
rect 10689 25109 10701 25143
rect 10735 25140 10747 25143
rect 10778 25140 10784 25152
rect 10735 25112 10784 25140
rect 10735 25109 10747 25112
rect 10689 25103 10747 25109
rect 10778 25100 10784 25112
rect 10836 25100 10842 25152
rect 11885 25143 11943 25149
rect 11885 25109 11897 25143
rect 11931 25140 11943 25143
rect 12066 25140 12072 25152
rect 11931 25112 12072 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 12066 25100 12072 25112
rect 12124 25100 12130 25152
rect 12526 25140 12532 25152
rect 12487 25112 12532 25140
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 18598 25140 18604 25152
rect 18559 25112 18604 25140
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 22675 25143 22733 25149
rect 22675 25109 22687 25143
rect 22721 25140 22733 25143
rect 23198 25140 23204 25152
rect 22721 25112 23204 25140
rect 22721 25109 22733 25112
rect 22675 25103 22733 25109
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 33594 25100 33600 25152
rect 33652 25140 33658 25152
rect 34977 25143 35035 25149
rect 34977 25140 34989 25143
rect 33652 25112 34989 25140
rect 33652 25100 33658 25112
rect 34977 25109 34989 25112
rect 35023 25109 35035 25143
rect 34977 25103 35035 25109
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 13354 24896 13360 24948
rect 13412 24936 13418 24948
rect 13541 24939 13599 24945
rect 13541 24936 13553 24939
rect 13412 24908 13553 24936
rect 13412 24896 13418 24908
rect 13541 24905 13553 24908
rect 13587 24905 13599 24939
rect 13541 24899 13599 24905
rect 15286 24896 15292 24948
rect 15344 24936 15350 24948
rect 15933 24939 15991 24945
rect 15933 24936 15945 24939
rect 15344 24908 15945 24936
rect 15344 24896 15350 24908
rect 15933 24905 15945 24908
rect 15979 24905 15991 24939
rect 15933 24899 15991 24905
rect 22922 24896 22928 24948
rect 22980 24936 22986 24948
rect 23474 24936 23480 24948
rect 22980 24908 23480 24936
rect 22980 24896 22986 24908
rect 23474 24896 23480 24908
rect 23532 24936 23538 24948
rect 23569 24939 23627 24945
rect 23569 24936 23581 24939
rect 23532 24908 23581 24936
rect 23532 24896 23538 24908
rect 23569 24905 23581 24908
rect 23615 24905 23627 24939
rect 23569 24899 23627 24905
rect 33410 24896 33416 24948
rect 33468 24936 33474 24948
rect 42886 24936 42892 24948
rect 33468 24908 42892 24936
rect 33468 24896 33474 24908
rect 42886 24896 42892 24908
rect 42944 24896 42950 24948
rect 12066 24868 12072 24880
rect 12027 24840 12072 24868
rect 12066 24828 12072 24840
rect 12124 24828 12130 24880
rect 18598 24828 18604 24880
rect 18656 24828 18662 24880
rect 22554 24828 22560 24880
rect 22612 24828 22618 24880
rect 34425 24871 34483 24877
rect 34425 24868 34437 24871
rect 28368 24840 28948 24868
rect 13170 24760 13176 24812
rect 13228 24760 13234 24812
rect 14093 24803 14151 24809
rect 14093 24769 14105 24803
rect 14139 24769 14151 24803
rect 14918 24800 14924 24812
rect 14879 24772 14924 24800
rect 14093 24763 14151 24769
rect 11793 24735 11851 24741
rect 11793 24701 11805 24735
rect 11839 24732 11851 24735
rect 12526 24732 12532 24744
rect 11839 24704 12532 24732
rect 11839 24701 11851 24704
rect 11793 24695 11851 24701
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 14108 24732 14136 24763
rect 14918 24760 14924 24772
rect 14976 24760 14982 24812
rect 15838 24800 15844 24812
rect 15799 24772 15844 24800
rect 15838 24760 15844 24772
rect 15896 24760 15902 24812
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16114 24800 16120 24812
rect 16071 24772 16120 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 16114 24760 16120 24772
rect 16172 24760 16178 24812
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24800 20131 24803
rect 20806 24800 20812 24812
rect 20119 24772 20812 24800
rect 20119 24769 20131 24772
rect 20073 24763 20131 24769
rect 20806 24760 20812 24772
rect 20864 24760 20870 24812
rect 21266 24800 21272 24812
rect 21227 24772 21272 24800
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 25041 24803 25099 24809
rect 25041 24769 25053 24803
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 14182 24732 14188 24744
rect 14095 24704 14188 24732
rect 14182 24692 14188 24704
rect 14240 24732 14246 24744
rect 17773 24735 17831 24741
rect 14240 24704 15148 24732
rect 14240 24692 14246 24704
rect 15120 24608 15148 24704
rect 17773 24701 17785 24735
rect 17819 24701 17831 24735
rect 18046 24732 18052 24744
rect 18007 24704 18052 24732
rect 17773 24695 17831 24701
rect 14185 24599 14243 24605
rect 14185 24565 14197 24599
rect 14231 24596 14243 24599
rect 14274 24596 14280 24608
rect 14231 24568 14280 24596
rect 14231 24565 14243 24568
rect 14185 24559 14243 24565
rect 14274 24556 14280 24568
rect 14332 24556 14338 24608
rect 15102 24596 15108 24608
rect 15063 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 17788 24596 17816 24695
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 21174 24692 21180 24744
rect 21232 24732 21238 24744
rect 21821 24735 21879 24741
rect 21821 24732 21833 24735
rect 21232 24704 21833 24732
rect 21232 24692 21238 24704
rect 21821 24701 21833 24704
rect 21867 24701 21879 24735
rect 22097 24735 22155 24741
rect 22097 24732 22109 24735
rect 21821 24695 21879 24701
rect 21928 24704 22109 24732
rect 20165 24667 20223 24673
rect 20165 24664 20177 24667
rect 19076 24636 20177 24664
rect 19076 24596 19104 24636
rect 20165 24633 20177 24636
rect 20211 24633 20223 24667
rect 20165 24627 20223 24633
rect 21085 24667 21143 24673
rect 21085 24633 21097 24667
rect 21131 24664 21143 24667
rect 21928 24664 21956 24704
rect 22097 24701 22109 24704
rect 22143 24701 22155 24735
rect 25056 24732 25084 24763
rect 26694 24760 26700 24812
rect 26752 24800 26758 24812
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26752 24772 26985 24800
rect 26752 24760 26758 24772
rect 26973 24769 26985 24772
rect 27019 24800 27031 24803
rect 28368 24800 28396 24840
rect 27019 24772 28396 24800
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 28442 24760 28448 24812
rect 28500 24800 28506 24812
rect 28629 24803 28687 24809
rect 28629 24800 28641 24803
rect 28500 24772 28641 24800
rect 28500 24760 28506 24772
rect 28629 24769 28641 24772
rect 28675 24769 28687 24803
rect 28629 24763 28687 24769
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 28813 24803 28871 24809
rect 28813 24800 28825 24803
rect 28776 24772 28825 24800
rect 28776 24760 28782 24772
rect 28813 24769 28825 24772
rect 28859 24769 28871 24803
rect 28920 24800 28948 24840
rect 34256 24840 34437 24868
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 28920 24772 32137 24800
rect 28813 24763 28871 24769
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 33594 24800 33600 24812
rect 33555 24772 33600 24800
rect 32125 24763 32183 24769
rect 33594 24760 33600 24772
rect 33652 24760 33658 24812
rect 33689 24803 33747 24809
rect 33689 24769 33701 24803
rect 33735 24800 33747 24803
rect 34256 24800 34284 24840
rect 34425 24837 34437 24840
rect 34471 24837 34483 24871
rect 34425 24831 34483 24837
rect 33735 24772 34284 24800
rect 36081 24803 36139 24809
rect 33735 24769 33747 24772
rect 33689 24763 33747 24769
rect 36081 24769 36093 24803
rect 36127 24800 36139 24803
rect 38654 24800 38660 24812
rect 36127 24772 38660 24800
rect 36127 24769 36139 24772
rect 36081 24763 36139 24769
rect 38654 24760 38660 24772
rect 38712 24760 38718 24812
rect 46290 24800 46296 24812
rect 41386 24772 46296 24800
rect 25222 24732 25228 24744
rect 25056 24704 25228 24732
rect 22097 24695 22155 24701
rect 25222 24692 25228 24704
rect 25280 24732 25286 24744
rect 33962 24732 33968 24744
rect 25280 24704 33968 24732
rect 25280 24692 25286 24704
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 34238 24732 34244 24744
rect 34199 24704 34244 24732
rect 34238 24692 34244 24704
rect 34296 24692 34302 24744
rect 21131 24636 21956 24664
rect 21131 24633 21143 24636
rect 21085 24627 21143 24633
rect 24670 24624 24676 24676
rect 24728 24664 24734 24676
rect 41386 24664 41414 24772
rect 46290 24760 46296 24772
rect 46348 24760 46354 24812
rect 46382 24760 46388 24812
rect 46440 24800 46446 24812
rect 46842 24800 46848 24812
rect 46440 24772 46485 24800
rect 46803 24772 46848 24800
rect 46440 24760 46446 24772
rect 46842 24760 46848 24772
rect 46900 24760 46906 24812
rect 46934 24760 46940 24812
rect 46992 24800 46998 24812
rect 46992 24772 47037 24800
rect 46992 24760 46998 24772
rect 47486 24760 47492 24812
rect 47544 24800 47550 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47544 24772 47593 24800
rect 47544 24760 47550 24772
rect 47581 24769 47593 24772
rect 47627 24800 47639 24803
rect 47946 24800 47952 24812
rect 47627 24772 47952 24800
rect 47627 24769 47639 24772
rect 47581 24763 47639 24769
rect 47946 24760 47952 24772
rect 48004 24760 48010 24812
rect 45922 24692 45928 24744
rect 45980 24732 45986 24744
rect 46474 24732 46480 24744
rect 45980 24704 46480 24732
rect 45980 24692 45986 24704
rect 46474 24692 46480 24704
rect 46532 24692 46538 24744
rect 24728 24636 41414 24664
rect 46201 24667 46259 24673
rect 24728 24624 24734 24636
rect 46201 24633 46213 24667
rect 46247 24664 46259 24667
rect 47578 24664 47584 24676
rect 46247 24636 47584 24664
rect 46247 24633 46259 24636
rect 46201 24627 46259 24633
rect 47578 24624 47584 24636
rect 47636 24624 47642 24676
rect 19518 24596 19524 24608
rect 17788 24568 19104 24596
rect 19431 24568 19524 24596
rect 19518 24556 19524 24568
rect 19576 24596 19582 24608
rect 20254 24596 20260 24608
rect 19576 24568 20260 24596
rect 19576 24556 19582 24568
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 25130 24596 25136 24608
rect 25091 24568 25136 24596
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 27154 24596 27160 24608
rect 27115 24568 27160 24596
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 28721 24599 28779 24605
rect 28721 24565 28733 24599
rect 28767 24596 28779 24599
rect 29546 24596 29552 24608
rect 28767 24568 29552 24596
rect 28767 24565 28779 24568
rect 28721 24559 28779 24565
rect 29546 24556 29552 24568
rect 29604 24556 29610 24608
rect 31662 24556 31668 24608
rect 31720 24596 31726 24608
rect 32309 24599 32367 24605
rect 32309 24596 32321 24599
rect 31720 24568 32321 24596
rect 31720 24556 31726 24568
rect 32309 24565 32321 24568
rect 32355 24565 32367 24599
rect 32309 24559 32367 24565
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 47673 24599 47731 24605
rect 47673 24596 47685 24599
rect 46532 24568 47685 24596
rect 46532 24556 46538 24568
rect 47673 24565 47685 24568
rect 47719 24565 47731 24599
rect 47673 24559 47731 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 13170 24352 13176 24404
rect 13228 24392 13234 24404
rect 13265 24395 13323 24401
rect 13265 24392 13277 24395
rect 13228 24364 13277 24392
rect 13228 24352 13234 24364
rect 13265 24361 13277 24364
rect 13311 24361 13323 24395
rect 19426 24392 19432 24404
rect 19387 24364 19432 24392
rect 13265 24355 13323 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 21174 24392 21180 24404
rect 21135 24364 21180 24392
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 22465 24395 22523 24401
rect 22465 24392 22477 24395
rect 21324 24364 22477 24392
rect 21324 24352 21330 24364
rect 22465 24361 22477 24364
rect 22511 24361 22523 24395
rect 33597 24395 33655 24401
rect 22465 24355 22523 24361
rect 23308 24364 31754 24392
rect 10042 24324 10048 24336
rect 10003 24296 10048 24324
rect 10042 24284 10048 24296
rect 10100 24284 10106 24336
rect 12434 24324 12440 24336
rect 10152 24296 12440 24324
rect 9122 24188 9128 24200
rect 9035 24160 9128 24188
rect 9122 24148 9128 24160
rect 9180 24188 9186 24200
rect 10152 24188 10180 24296
rect 12434 24284 12440 24296
rect 12492 24324 12498 24336
rect 12621 24327 12679 24333
rect 12621 24324 12633 24327
rect 12492 24296 12633 24324
rect 12492 24284 12498 24296
rect 12621 24293 12633 24296
rect 12667 24293 12679 24327
rect 15378 24324 15384 24336
rect 12621 24287 12679 24293
rect 14108 24296 15384 24324
rect 13078 24256 13084 24268
rect 10612 24228 13084 24256
rect 10612 24197 10640 24228
rect 13078 24216 13084 24228
rect 13136 24256 13142 24268
rect 14108 24265 14136 24296
rect 15378 24284 15384 24296
rect 15436 24284 15442 24336
rect 17402 24284 17408 24336
rect 17460 24324 17466 24336
rect 19518 24324 19524 24336
rect 17460 24296 19524 24324
rect 17460 24284 17466 24296
rect 19518 24284 19524 24296
rect 19576 24284 19582 24336
rect 22373 24327 22431 24333
rect 22373 24293 22385 24327
rect 22419 24324 22431 24327
rect 23017 24327 23075 24333
rect 23017 24324 23029 24327
rect 22419 24296 23029 24324
rect 22419 24293 22431 24296
rect 22373 24287 22431 24293
rect 23017 24293 23029 24296
rect 23063 24293 23075 24327
rect 23017 24287 23075 24293
rect 14093 24259 14151 24265
rect 13136 24228 13216 24256
rect 13136 24216 13142 24228
rect 9180 24160 10180 24188
rect 10597 24191 10655 24197
rect 9180 24148 9186 24160
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 12526 24188 12532 24200
rect 12483 24160 12532 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 13188 24197 13216 24228
rect 14093 24225 14105 24259
rect 14139 24225 14151 24259
rect 14274 24256 14280 24268
rect 14235 24228 14280 24256
rect 14093 24219 14151 24225
rect 14274 24216 14280 24228
rect 14332 24216 14338 24268
rect 15562 24256 15568 24268
rect 15523 24228 15568 24256
rect 15562 24216 15568 24228
rect 15620 24216 15626 24268
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24256 18291 24259
rect 23308 24256 23336 24364
rect 24394 24324 24400 24336
rect 23400 24296 24400 24324
rect 23400 24265 23428 24296
rect 24394 24284 24400 24296
rect 24452 24284 24458 24336
rect 29086 24284 29092 24336
rect 29144 24324 29150 24336
rect 29549 24327 29607 24333
rect 29549 24324 29561 24327
rect 29144 24296 29561 24324
rect 29144 24284 29150 24296
rect 29549 24293 29561 24296
rect 29595 24293 29607 24327
rect 31726 24324 31754 24364
rect 33597 24361 33609 24395
rect 33643 24392 33655 24395
rect 34238 24392 34244 24404
rect 33643 24364 34244 24392
rect 33643 24361 33655 24364
rect 33597 24355 33655 24361
rect 34238 24352 34244 24364
rect 34296 24352 34302 24404
rect 43070 24352 43076 24404
rect 43128 24392 43134 24404
rect 43438 24392 43444 24404
rect 43128 24364 43444 24392
rect 43128 24352 43134 24364
rect 43438 24352 43444 24364
rect 43496 24392 43502 24404
rect 48222 24392 48228 24404
rect 43496 24364 48228 24392
rect 43496 24352 43502 24364
rect 48222 24352 48228 24364
rect 48280 24352 48286 24404
rect 40218 24324 40224 24336
rect 31726 24296 40224 24324
rect 29549 24287 29607 24293
rect 40218 24284 40224 24296
rect 40276 24284 40282 24336
rect 47762 24324 47768 24336
rect 46308 24296 47768 24324
rect 18279 24228 23336 24256
rect 23385 24259 23443 24265
rect 18279 24225 18291 24228
rect 18233 24219 18291 24225
rect 23385 24225 23397 24259
rect 23431 24225 23443 24259
rect 25130 24256 25136 24268
rect 25091 24228 25136 24256
rect 23385 24219 23443 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 26789 24259 26847 24265
rect 26789 24225 26801 24259
rect 26835 24256 26847 24259
rect 46014 24256 46020 24268
rect 26835 24228 46020 24256
rect 26835 24225 26847 24228
rect 26789 24219 26847 24225
rect 46014 24216 46020 24228
rect 46072 24216 46078 24268
rect 46308 24265 46336 24296
rect 47762 24284 47768 24296
rect 47820 24284 47826 24336
rect 46293 24259 46351 24265
rect 46293 24225 46305 24259
rect 46339 24225 46351 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46293 24219 46351 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 16393 24191 16451 24197
rect 16393 24157 16405 24191
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 20806 24188 20812 24200
rect 19475 24160 20812 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 3878 24080 3884 24132
rect 3936 24120 3942 24132
rect 9674 24120 9680 24132
rect 3936 24092 9260 24120
rect 9635 24092 9680 24120
rect 3936 24080 3942 24092
rect 9030 24012 9036 24064
rect 9088 24052 9094 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 9088 24024 9137 24052
rect 9088 24012 9094 24024
rect 9125 24021 9137 24024
rect 9171 24021 9183 24055
rect 9232 24052 9260 24092
rect 9674 24080 9680 24092
rect 9732 24080 9738 24132
rect 13998 24120 14004 24132
rect 9784 24092 14004 24120
rect 9784 24052 9812 24092
rect 13998 24080 14004 24092
rect 14056 24080 14062 24132
rect 14734 24080 14740 24132
rect 14792 24120 14798 24132
rect 16408 24120 16436 24151
rect 20806 24148 20812 24160
rect 20864 24188 20870 24200
rect 21177 24191 21235 24197
rect 21177 24188 21189 24191
rect 20864 24160 21189 24188
rect 20864 24148 20870 24160
rect 21177 24157 21189 24160
rect 21223 24188 21235 24191
rect 21726 24188 21732 24200
rect 21223 24160 21732 24188
rect 21223 24157 21235 24160
rect 21177 24151 21235 24157
rect 21726 24148 21732 24160
rect 21784 24148 21790 24200
rect 22002 24188 22008 24200
rect 21963 24160 22008 24188
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 23198 24188 23204 24200
rect 23159 24160 23204 24188
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 23474 24188 23480 24200
rect 23348 24160 23393 24188
rect 23435 24160 23480 24188
rect 23348 24148 23354 24160
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 24946 24188 24952 24200
rect 24907 24160 24952 24188
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 26878 24148 26884 24200
rect 26936 24188 26942 24200
rect 27249 24191 27307 24197
rect 27249 24188 27261 24191
rect 26936 24160 27261 24188
rect 26936 24148 26942 24160
rect 27249 24157 27261 24160
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 27525 24191 27583 24197
rect 27525 24157 27537 24191
rect 27571 24157 27583 24191
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 27525 24151 27583 24157
rect 28828 24160 29745 24188
rect 14792 24092 16436 24120
rect 16577 24123 16635 24129
rect 14792 24080 14798 24092
rect 16577 24089 16589 24123
rect 16623 24120 16635 24123
rect 16758 24120 16764 24132
rect 16623 24092 16764 24120
rect 16623 24089 16635 24092
rect 16577 24083 16635 24089
rect 16758 24080 16764 24092
rect 16816 24080 16822 24132
rect 24394 24080 24400 24132
rect 24452 24120 24458 24132
rect 27540 24120 27568 24151
rect 28442 24120 28448 24132
rect 24452 24092 28448 24120
rect 24452 24080 24458 24092
rect 28442 24080 28448 24092
rect 28500 24120 28506 24132
rect 28629 24123 28687 24129
rect 28629 24120 28641 24123
rect 28500 24092 28641 24120
rect 28500 24080 28506 24092
rect 28629 24089 28641 24092
rect 28675 24089 28687 24123
rect 28629 24083 28687 24089
rect 28718 24080 28724 24132
rect 28776 24120 28782 24132
rect 28828 24129 28856 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29834 24191 29892 24197
rect 29834 24157 29846 24191
rect 29880 24188 29892 24191
rect 30006 24188 30012 24200
rect 29880 24160 30012 24188
rect 29880 24157 29892 24160
rect 29834 24151 29892 24157
rect 30006 24148 30012 24160
rect 30064 24188 30070 24200
rect 30064 24160 30328 24188
rect 30064 24148 30070 24160
rect 28813 24123 28871 24129
rect 28813 24120 28825 24123
rect 28776 24092 28825 24120
rect 28776 24080 28782 24092
rect 28813 24089 28825 24092
rect 28859 24089 28871 24123
rect 28813 24083 28871 24089
rect 29270 24080 29276 24132
rect 29328 24120 29334 24132
rect 29549 24123 29607 24129
rect 29549 24120 29561 24123
rect 29328 24092 29561 24120
rect 29328 24080 29334 24092
rect 29549 24089 29561 24092
rect 29595 24089 29607 24123
rect 30300 24120 30328 24160
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 30469 24191 30527 24197
rect 30469 24188 30481 24191
rect 30432 24160 30481 24188
rect 30432 24148 30438 24160
rect 30469 24157 30481 24160
rect 30515 24157 30527 24191
rect 31662 24188 31668 24200
rect 31623 24160 31668 24188
rect 30469 24151 30527 24157
rect 31662 24148 31668 24160
rect 31720 24148 31726 24200
rect 33505 24191 33563 24197
rect 33505 24157 33517 24191
rect 33551 24157 33563 24191
rect 35066 24188 35072 24200
rect 35027 24160 35072 24188
rect 33505 24151 33563 24157
rect 33520 24120 33548 24151
rect 35066 24148 35072 24160
rect 35124 24148 35130 24200
rect 36906 24188 36912 24200
rect 36867 24160 36912 24188
rect 36906 24148 36912 24160
rect 36964 24148 36970 24200
rect 43070 24188 43076 24200
rect 43031 24160 43076 24188
rect 43070 24148 43076 24160
rect 43128 24148 43134 24200
rect 43254 24188 43260 24200
rect 43215 24160 43260 24188
rect 43254 24148 43260 24160
rect 43312 24148 43318 24200
rect 43898 24188 43904 24200
rect 43859 24160 43904 24188
rect 43898 24148 43904 24160
rect 43956 24148 43962 24200
rect 44085 24191 44143 24197
rect 44085 24157 44097 24191
rect 44131 24157 44143 24191
rect 44085 24151 44143 24157
rect 30300 24092 33548 24120
rect 35253 24123 35311 24129
rect 29549 24083 29607 24089
rect 35253 24089 35265 24123
rect 35299 24120 35311 24123
rect 35802 24120 35808 24132
rect 35299 24092 35808 24120
rect 35299 24089 35311 24092
rect 35253 24083 35311 24089
rect 35802 24080 35808 24092
rect 35860 24080 35866 24132
rect 43441 24123 43499 24129
rect 43441 24089 43453 24123
rect 43487 24120 43499 24123
rect 44100 24120 44128 24151
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45649 24191 45707 24197
rect 45649 24188 45661 24191
rect 45612 24160 45661 24188
rect 45612 24148 45618 24160
rect 45649 24157 45661 24160
rect 45695 24157 45707 24191
rect 45649 24151 45707 24157
rect 45833 24191 45891 24197
rect 45833 24157 45845 24191
rect 45879 24157 45891 24191
rect 45833 24151 45891 24157
rect 43487 24092 44128 24120
rect 45848 24120 45876 24151
rect 47394 24120 47400 24132
rect 45848 24092 47400 24120
rect 43487 24089 43499 24092
rect 43441 24083 43499 24089
rect 47394 24080 47400 24092
rect 47452 24080 47458 24132
rect 10134 24052 10140 24064
rect 9232 24024 9812 24052
rect 10095 24024 10140 24052
rect 9125 24015 9183 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10686 24052 10692 24064
rect 10647 24024 10692 24052
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 28997 24055 29055 24061
rect 28997 24021 29009 24055
rect 29043 24052 29055 24055
rect 29638 24052 29644 24064
rect 29043 24024 29644 24052
rect 29043 24021 29055 24024
rect 28997 24015 29055 24021
rect 29638 24012 29644 24024
rect 29696 24012 29702 24064
rect 30285 24055 30343 24061
rect 30285 24021 30297 24055
rect 30331 24052 30343 24055
rect 30650 24052 30656 24064
rect 30331 24024 30656 24052
rect 30331 24021 30343 24024
rect 30285 24015 30343 24021
rect 30650 24012 30656 24024
rect 30708 24012 30714 24064
rect 31754 24012 31760 24064
rect 31812 24052 31818 24064
rect 43990 24052 43996 24064
rect 31812 24024 31857 24052
rect 43951 24024 43996 24052
rect 31812 24012 31818 24024
rect 43990 24012 43996 24024
rect 44048 24012 44054 24064
rect 45833 24055 45891 24061
rect 45833 24021 45845 24055
rect 45879 24052 45891 24055
rect 47670 24052 47676 24064
rect 45879 24024 47676 24052
rect 45879 24021 45891 24024
rect 45833 24015 45891 24021
rect 47670 24012 47676 24024
rect 47728 24012 47734 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 9766 23848 9772 23860
rect 8404 23820 9772 23848
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 8404 23721 8432 23820
rect 9766 23808 9772 23820
rect 9824 23848 9830 23860
rect 15841 23851 15899 23857
rect 15841 23848 15853 23851
rect 9824 23820 15853 23848
rect 9824 23808 9830 23820
rect 15841 23817 15853 23820
rect 15887 23817 15899 23851
rect 16758 23848 16764 23860
rect 16719 23820 16764 23848
rect 15841 23811 15899 23817
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 22373 23851 22431 23857
rect 22373 23817 22385 23851
rect 22419 23848 22431 23851
rect 22554 23848 22560 23860
rect 22419 23820 22560 23848
rect 22419 23817 22431 23820
rect 22373 23811 22431 23817
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 29270 23808 29276 23860
rect 29328 23848 29334 23860
rect 31481 23851 31539 23857
rect 31481 23848 31493 23851
rect 29328 23820 31493 23848
rect 29328 23808 29334 23820
rect 31481 23817 31493 23820
rect 31527 23848 31539 23851
rect 35066 23848 35072 23860
rect 31527 23820 35072 23848
rect 31527 23817 31539 23820
rect 31481 23811 31539 23817
rect 35066 23808 35072 23820
rect 35124 23808 35130 23860
rect 35802 23848 35808 23860
rect 35763 23820 35808 23848
rect 35802 23808 35808 23820
rect 35860 23808 35866 23860
rect 43898 23848 43904 23860
rect 42444 23820 43904 23848
rect 8481 23783 8539 23789
rect 8481 23749 8493 23783
rect 8527 23780 8539 23783
rect 9217 23783 9275 23789
rect 9217 23780 9229 23783
rect 8527 23752 9229 23780
rect 8527 23749 8539 23752
rect 8481 23743 8539 23749
rect 9217 23749 9229 23752
rect 9263 23749 9275 23783
rect 15378 23780 15384 23792
rect 9217 23743 9275 23749
rect 13096 23752 15384 23780
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23681 8447 23715
rect 11698 23712 11704 23724
rect 8389 23675 8447 23681
rect 10704 23684 11704 23712
rect 9033 23647 9091 23653
rect 9033 23613 9045 23647
rect 9079 23644 9091 23647
rect 10704 23644 10732 23684
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 13096 23721 13124 23752
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 15749 23783 15807 23789
rect 15749 23749 15761 23783
rect 15795 23780 15807 23783
rect 15795 23752 17540 23780
rect 15795 23749 15807 23752
rect 15749 23743 15807 23749
rect 17512 23724 17540 23752
rect 23290 23740 23296 23792
rect 23348 23780 23354 23792
rect 23842 23780 23848 23792
rect 23348 23752 23848 23780
rect 23348 23740 23354 23752
rect 23842 23740 23848 23752
rect 23900 23780 23906 23792
rect 25593 23783 25651 23789
rect 23900 23752 23980 23780
rect 23900 23740 23906 23752
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 15102 23672 15108 23724
rect 15160 23712 15166 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 15160 23684 16681 23712
rect 15160 23672 15166 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 17494 23712 17500 23724
rect 17455 23684 17500 23712
rect 16669 23675 16727 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23712 19579 23715
rect 20346 23712 20352 23724
rect 19567 23684 20352 23712
rect 19567 23681 19579 23684
rect 19521 23675 19579 23681
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 22278 23712 22284 23724
rect 22239 23684 22284 23712
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 23017 23715 23075 23721
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 23198 23712 23204 23724
rect 23063 23684 23204 23712
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 23198 23672 23204 23684
rect 23256 23712 23262 23724
rect 23952 23721 23980 23752
rect 25593 23749 25605 23783
rect 25639 23780 25651 23783
rect 26878 23780 26884 23792
rect 25639 23752 26884 23780
rect 25639 23749 25651 23752
rect 25593 23743 25651 23749
rect 26878 23740 26884 23752
rect 26936 23740 26942 23792
rect 29178 23740 29184 23792
rect 29236 23780 29242 23792
rect 30009 23783 30067 23789
rect 30009 23780 30021 23783
rect 29236 23752 30021 23780
rect 29236 23740 29242 23752
rect 30009 23749 30021 23752
rect 30055 23749 30067 23783
rect 32217 23783 32275 23789
rect 32217 23780 32229 23783
rect 31234 23752 32229 23780
rect 30009 23743 30067 23749
rect 32217 23749 32229 23752
rect 32263 23749 32275 23783
rect 32217 23743 32275 23749
rect 34698 23740 34704 23792
rect 34756 23780 34762 23792
rect 35253 23783 35311 23789
rect 35253 23780 35265 23783
rect 34756 23752 35265 23780
rect 34756 23740 34762 23752
rect 35253 23749 35265 23752
rect 35299 23780 35311 23783
rect 41046 23780 41052 23792
rect 35299 23752 41052 23780
rect 35299 23749 35311 23752
rect 35253 23743 35311 23749
rect 41046 23740 41052 23752
rect 41104 23740 41110 23792
rect 42444 23789 42472 23820
rect 43898 23808 43904 23820
rect 43956 23808 43962 23860
rect 45554 23808 45560 23860
rect 45612 23848 45618 23860
rect 45612 23820 47624 23848
rect 45612 23808 45618 23820
rect 42429 23783 42487 23789
rect 42429 23749 42441 23783
rect 42475 23749 42487 23783
rect 42429 23743 42487 23749
rect 42613 23783 42671 23789
rect 42613 23749 42625 23783
rect 42659 23780 42671 23783
rect 43070 23780 43076 23792
rect 42659 23752 43076 23780
rect 42659 23749 42671 23752
rect 42613 23743 42671 23749
rect 43070 23740 43076 23752
rect 43128 23740 43134 23792
rect 45097 23783 45155 23789
rect 45097 23749 45109 23783
rect 45143 23780 45155 23783
rect 45646 23780 45652 23792
rect 45143 23752 45652 23780
rect 45143 23749 45155 23752
rect 45097 23743 45155 23749
rect 45646 23740 45652 23752
rect 45704 23780 45710 23792
rect 46106 23780 46112 23792
rect 45704 23752 46112 23780
rect 45704 23740 45710 23752
rect 46106 23740 46112 23752
rect 46164 23740 46170 23792
rect 23937 23715 23995 23721
rect 23256 23684 23428 23712
rect 23256 23672 23262 23684
rect 10870 23644 10876 23656
rect 9079 23616 10732 23644
rect 10831 23616 10876 23644
rect 9079 23613 9091 23616
rect 9033 23607 9091 23613
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 13265 23647 13323 23653
rect 13265 23613 13277 23647
rect 13311 23644 13323 23647
rect 13906 23644 13912 23656
rect 13311 23616 13912 23644
rect 13311 23613 13323 23616
rect 13265 23607 13323 23613
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 13998 23604 14004 23656
rect 14056 23644 14062 23656
rect 17862 23644 17868 23656
rect 14056 23616 14101 23644
rect 17823 23616 17868 23644
rect 14056 23604 14062 23616
rect 17862 23604 17868 23616
rect 17920 23644 17926 23656
rect 18782 23644 18788 23656
rect 17920 23616 18788 23644
rect 17920 23604 17926 23616
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 23106 23644 23112 23656
rect 19306 23616 23112 23644
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 19306 23576 19334 23616
rect 23106 23604 23112 23616
rect 23164 23604 23170 23656
rect 2087 23548 19334 23576
rect 23400 23576 23428 23684
rect 23937 23681 23949 23715
rect 23983 23681 23995 23715
rect 27430 23712 27436 23724
rect 27391 23684 27436 23712
rect 23937 23675 23995 23681
rect 27430 23672 27436 23684
rect 27488 23672 27494 23724
rect 28353 23715 28411 23721
rect 28353 23681 28365 23715
rect 28399 23712 28411 23715
rect 28810 23712 28816 23724
rect 28399 23684 28816 23712
rect 28399 23681 28411 23684
rect 28353 23675 28411 23681
rect 28810 23672 28816 23684
rect 28868 23672 28874 23724
rect 28994 23712 29000 23724
rect 28920 23684 29000 23712
rect 23661 23647 23719 23653
rect 23661 23613 23673 23647
rect 23707 23644 23719 23647
rect 24026 23644 24032 23656
rect 23707 23616 24032 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24026 23604 24032 23616
rect 24084 23604 24090 23656
rect 27525 23647 27583 23653
rect 27525 23613 27537 23647
rect 27571 23644 27583 23647
rect 28258 23644 28264 23656
rect 27571 23616 28264 23644
rect 27571 23613 27583 23616
rect 27525 23607 27583 23613
rect 28258 23604 28264 23616
rect 28316 23604 28322 23656
rect 28629 23647 28687 23653
rect 28629 23613 28641 23647
rect 28675 23644 28687 23647
rect 28718 23644 28724 23656
rect 28675 23616 28724 23644
rect 28675 23613 28687 23616
rect 28629 23607 28687 23613
rect 28718 23604 28724 23616
rect 28776 23604 28782 23656
rect 25682 23576 25688 23588
rect 23400 23548 25688 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 25682 23536 25688 23548
rect 25740 23536 25746 23588
rect 25777 23579 25835 23585
rect 25777 23545 25789 23579
rect 25823 23576 25835 23579
rect 28920 23576 28948 23684
rect 28994 23672 29000 23684
rect 29052 23672 29058 23724
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29656 23684 29745 23712
rect 25823 23548 28948 23576
rect 25823 23545 25835 23548
rect 25777 23539 25835 23545
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 19576 23480 19625 23508
rect 19576 23468 19582 23480
rect 19613 23477 19625 23480
rect 19659 23477 19671 23511
rect 19613 23471 19671 23477
rect 23109 23511 23167 23517
rect 23109 23477 23121 23511
rect 23155 23508 23167 23511
rect 24670 23508 24676 23520
rect 23155 23480 24676 23508
rect 23155 23477 23167 23480
rect 23109 23471 23167 23477
rect 24670 23468 24676 23480
rect 24728 23468 24734 23520
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25792 23508 25820 23539
rect 27798 23508 27804 23520
rect 24912 23480 25820 23508
rect 27759 23480 27804 23508
rect 24912 23468 24918 23480
rect 27798 23468 27804 23480
rect 27856 23468 27862 23520
rect 29656 23508 29684 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 31662 23672 31668 23724
rect 31720 23712 31726 23724
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31720 23684 32137 23712
rect 31720 23672 31726 23684
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 33502 23712 33508 23724
rect 33463 23684 33508 23712
rect 32125 23675 32183 23681
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 35434 23672 35440 23724
rect 35492 23712 35498 23724
rect 35713 23715 35771 23721
rect 35713 23712 35725 23715
rect 35492 23684 35725 23712
rect 35492 23672 35498 23684
rect 35713 23681 35725 23684
rect 35759 23712 35771 23715
rect 35802 23712 35808 23724
rect 35759 23684 35808 23712
rect 35759 23681 35771 23684
rect 35713 23675 35771 23681
rect 35802 23672 35808 23684
rect 35860 23672 35866 23724
rect 39206 23712 39212 23724
rect 39167 23684 39212 23712
rect 39206 23672 39212 23684
rect 39264 23672 39270 23724
rect 40034 23712 40040 23724
rect 39995 23684 40040 23712
rect 40034 23672 40040 23684
rect 40092 23672 40098 23724
rect 42705 23715 42763 23721
rect 42705 23681 42717 23715
rect 42751 23712 42763 23715
rect 43162 23712 43168 23724
rect 42751 23684 43168 23712
rect 42751 23681 42763 23684
rect 42705 23675 42763 23681
rect 43162 23672 43168 23684
rect 43220 23712 43226 23724
rect 43257 23715 43315 23721
rect 43257 23712 43269 23715
rect 43220 23684 43269 23712
rect 43220 23672 43226 23684
rect 43257 23681 43269 23684
rect 43303 23681 43315 23715
rect 43990 23712 43996 23724
rect 43951 23684 43996 23712
rect 43257 23675 43315 23681
rect 43990 23672 43996 23684
rect 44048 23672 44054 23724
rect 47596 23721 47624 23820
rect 45741 23715 45799 23721
rect 45741 23681 45753 23715
rect 45787 23712 45799 23715
rect 47581 23715 47639 23721
rect 45787 23684 46888 23712
rect 45787 23681 45799 23684
rect 45741 23675 45799 23681
rect 38378 23604 38384 23656
rect 38436 23644 38442 23656
rect 39117 23647 39175 23653
rect 39117 23644 39129 23647
rect 38436 23616 39129 23644
rect 38436 23604 38442 23616
rect 39117 23613 39129 23616
rect 39163 23613 39175 23647
rect 40218 23644 40224 23656
rect 40179 23616 40224 23644
rect 39117 23607 39175 23613
rect 40218 23604 40224 23616
rect 40276 23604 40282 23656
rect 41874 23644 41880 23656
rect 41835 23616 41880 23644
rect 41874 23604 41880 23616
rect 41932 23604 41938 23656
rect 46106 23604 46112 23656
rect 46164 23644 46170 23656
rect 46201 23647 46259 23653
rect 46201 23644 46213 23647
rect 46164 23616 46213 23644
rect 46164 23604 46170 23616
rect 46201 23613 46213 23616
rect 46247 23613 46259 23647
rect 46201 23607 46259 23613
rect 46477 23647 46535 23653
rect 46477 23613 46489 23647
rect 46523 23613 46535 23647
rect 46860 23644 46888 23684
rect 47581 23681 47593 23715
rect 47627 23712 47639 23715
rect 47946 23712 47952 23724
rect 47627 23684 47952 23712
rect 47627 23681 47639 23684
rect 47581 23675 47639 23681
rect 47946 23672 47952 23684
rect 48004 23672 48010 23724
rect 48041 23647 48099 23653
rect 48041 23644 48053 23647
rect 46860 23616 48053 23644
rect 46477 23607 46535 23613
rect 48041 23613 48053 23616
rect 48087 23613 48099 23647
rect 48041 23607 48099 23613
rect 42886 23536 42892 23588
rect 42944 23576 42950 23588
rect 46492 23576 46520 23607
rect 42944 23548 46520 23576
rect 42944 23536 42950 23548
rect 30006 23508 30012 23520
rect 29656 23480 30012 23508
rect 30006 23468 30012 23480
rect 30064 23468 30070 23520
rect 39485 23511 39543 23517
rect 39485 23477 39497 23511
rect 39531 23508 39543 23511
rect 40034 23508 40040 23520
rect 39531 23480 40040 23508
rect 39531 23477 39543 23480
rect 39485 23471 39543 23477
rect 40034 23468 40040 23480
rect 40092 23468 40098 23520
rect 41414 23468 41420 23520
rect 41472 23508 41478 23520
rect 42429 23511 42487 23517
rect 42429 23508 42441 23511
rect 41472 23480 42441 23508
rect 41472 23468 41478 23480
rect 42429 23477 42441 23480
rect 42475 23477 42487 23511
rect 42429 23471 42487 23477
rect 45554 23468 45560 23520
rect 45612 23508 45618 23520
rect 45612 23480 45657 23508
rect 45612 23468 45618 23480
rect 47394 23468 47400 23520
rect 47452 23508 47458 23520
rect 47673 23511 47731 23517
rect 47673 23508 47685 23511
rect 47452 23480 47685 23508
rect 47452 23468 47458 23480
rect 47673 23477 47685 23480
rect 47719 23477 47731 23511
rect 47673 23471 47731 23477
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 10410 23264 10416 23316
rect 10468 23304 10474 23316
rect 10781 23307 10839 23313
rect 10781 23304 10793 23307
rect 10468 23276 10793 23304
rect 10468 23264 10474 23276
rect 10781 23273 10793 23276
rect 10827 23273 10839 23307
rect 13078 23304 13084 23316
rect 13039 23276 13084 23304
rect 10781 23267 10839 23273
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23304 18475 23307
rect 18506 23304 18512 23316
rect 18463 23276 18512 23304
rect 18463 23273 18475 23276
rect 18417 23267 18475 23273
rect 18506 23264 18512 23276
rect 18564 23264 18570 23316
rect 25406 23304 25412 23316
rect 19168 23276 25412 23304
rect 9030 23168 9036 23180
rect 8991 23140 9036 23168
rect 9030 23128 9036 23140
rect 9088 23128 9094 23180
rect 14918 23128 14924 23180
rect 14976 23168 14982 23180
rect 14976 23140 18184 23168
rect 14976 23128 14982 23140
rect 11330 23100 11336 23112
rect 11291 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 13814 23100 13820 23112
rect 12943 23072 13820 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 13814 23060 13820 23072
rect 13872 23100 13878 23112
rect 15102 23100 15108 23112
rect 13872 23072 15108 23100
rect 13872 23060 13878 23072
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 15746 23100 15752 23112
rect 15707 23072 15752 23100
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 17586 23100 17592 23112
rect 17547 23072 17592 23100
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 18156 23109 18184 23140
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 19168 23100 19196 23276
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 25501 23307 25559 23313
rect 25501 23273 25513 23307
rect 25547 23273 25559 23307
rect 25501 23267 25559 23273
rect 24210 23196 24216 23248
rect 24268 23236 24274 23248
rect 24765 23239 24823 23245
rect 24765 23236 24777 23239
rect 24268 23208 24777 23236
rect 24268 23196 24274 23208
rect 24765 23205 24777 23208
rect 24811 23205 24823 23239
rect 24765 23199 24823 23205
rect 25038 23196 25044 23248
rect 25096 23236 25102 23248
rect 25516 23236 25544 23267
rect 25590 23264 25596 23316
rect 25648 23304 25654 23316
rect 28718 23304 28724 23316
rect 25648 23276 27936 23304
rect 28679 23276 28724 23304
rect 25648 23264 25654 23276
rect 25682 23236 25688 23248
rect 25096 23208 25544 23236
rect 25643 23208 25688 23236
rect 25096 23196 25102 23208
rect 25682 23196 25688 23208
rect 25740 23196 25746 23248
rect 19518 23168 19524 23180
rect 19479 23140 19524 23168
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 22097 23171 22155 23177
rect 22097 23137 22109 23171
rect 22143 23168 22155 23171
rect 24397 23171 24455 23177
rect 24397 23168 24409 23171
rect 22143 23140 24409 23168
rect 22143 23137 22155 23140
rect 22097 23131 22155 23137
rect 24397 23137 24409 23140
rect 24443 23137 24455 23171
rect 24397 23131 24455 23137
rect 24670 23128 24676 23180
rect 24728 23168 24734 23180
rect 24857 23171 24915 23177
rect 24857 23168 24869 23171
rect 24728 23140 24869 23168
rect 24728 23128 24734 23140
rect 24857 23137 24869 23140
rect 24903 23137 24915 23171
rect 24857 23131 24915 23137
rect 26513 23171 26571 23177
rect 26513 23137 26525 23171
rect 26559 23168 26571 23171
rect 27798 23168 27804 23180
rect 26559 23140 27804 23168
rect 26559 23137 26571 23140
rect 26513 23131 26571 23137
rect 27798 23128 27804 23140
rect 27856 23128 27862 23180
rect 18187 23072 19196 23100
rect 19245 23103 19303 23109
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 21818 23100 21824 23112
rect 21779 23072 21824 23100
rect 19245 23063 19303 23069
rect 9309 23035 9367 23041
rect 9309 23001 9321 23035
rect 9355 23032 9367 23035
rect 9582 23032 9588 23044
rect 9355 23004 9588 23032
rect 9355 23001 9367 23004
rect 9309 22995 9367 23001
rect 9582 22992 9588 23004
rect 9640 22992 9646 23044
rect 10686 23032 10692 23044
rect 10534 23004 10692 23032
rect 10686 22992 10692 23004
rect 10744 22992 10750 23044
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23032 14611 23035
rect 15930 23032 15936 23044
rect 14599 23004 15608 23032
rect 15891 23004 15936 23032
rect 14599 23001 14611 23004
rect 14553 22995 14611 23001
rect 11425 22967 11483 22973
rect 11425 22933 11437 22967
rect 11471 22964 11483 22967
rect 11698 22964 11704 22976
rect 11471 22936 11704 22964
rect 11471 22933 11483 22936
rect 11425 22927 11483 22933
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 13630 22924 13636 22976
rect 13688 22964 13694 22976
rect 14645 22967 14703 22973
rect 14645 22964 14657 22967
rect 13688 22936 14657 22964
rect 13688 22924 13694 22936
rect 14645 22933 14657 22936
rect 14691 22933 14703 22967
rect 15580 22964 15608 23004
rect 15930 22992 15936 23004
rect 15988 22992 15994 23044
rect 18690 22992 18696 23044
rect 18748 23032 18754 23044
rect 19260 23032 19288 23063
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 23382 23060 23388 23112
rect 23440 23100 23446 23112
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 23440 23072 24593 23100
rect 23440 23060 23446 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 26234 23100 26240 23112
rect 26195 23072 26240 23100
rect 24581 23063 24639 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 27908 23100 27936 23276
rect 28718 23264 28724 23276
rect 28776 23264 28782 23316
rect 28810 23264 28816 23316
rect 28868 23304 28874 23316
rect 29917 23307 29975 23313
rect 28868 23276 29040 23304
rect 28868 23264 28874 23276
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 28902 23236 28908 23248
rect 28316 23208 28908 23236
rect 28316 23196 28322 23208
rect 28902 23196 28908 23208
rect 28960 23196 28966 23248
rect 29012 23236 29040 23276
rect 29917 23273 29929 23307
rect 29963 23304 29975 23307
rect 30374 23304 30380 23316
rect 29963 23276 30380 23304
rect 29963 23273 29975 23276
rect 29917 23267 29975 23273
rect 30374 23264 30380 23276
rect 30432 23264 30438 23316
rect 32122 23304 32128 23316
rect 30484 23276 32128 23304
rect 30484 23236 30512 23276
rect 32122 23264 32128 23276
rect 32180 23264 32186 23316
rect 46750 23304 46756 23316
rect 41386 23276 46756 23304
rect 29012 23208 30512 23236
rect 33962 23196 33968 23248
rect 34020 23236 34026 23248
rect 41386 23236 41414 23276
rect 46750 23264 46756 23276
rect 46808 23264 46814 23316
rect 34020 23208 41414 23236
rect 43257 23239 43315 23245
rect 34020 23196 34026 23208
rect 43257 23205 43269 23239
rect 43303 23236 43315 23239
rect 43898 23236 43904 23248
rect 43303 23208 43904 23236
rect 43303 23205 43315 23208
rect 43257 23199 43315 23205
rect 43898 23196 43904 23208
rect 43956 23196 43962 23248
rect 44269 23239 44327 23245
rect 44269 23205 44281 23239
rect 44315 23236 44327 23239
rect 44315 23208 45968 23236
rect 44315 23205 44327 23208
rect 44269 23199 44327 23205
rect 29546 23168 29552 23180
rect 29507 23140 29552 23168
rect 29546 23128 29552 23140
rect 29604 23128 29610 23180
rect 30650 23168 30656 23180
rect 30611 23140 30656 23168
rect 30650 23128 30656 23140
rect 30708 23128 30714 23180
rect 40034 23168 40040 23180
rect 39995 23140 40040 23168
rect 40034 23128 40040 23140
rect 40092 23128 40098 23180
rect 40126 23128 40132 23180
rect 40184 23168 40190 23180
rect 40865 23171 40923 23177
rect 40865 23168 40877 23171
rect 40184 23140 40877 23168
rect 40184 23128 40190 23140
rect 40865 23137 40877 23140
rect 40911 23137 40923 23171
rect 42613 23171 42671 23177
rect 40865 23131 40923 23137
rect 41524 23140 42472 23168
rect 27908 23072 29408 23100
rect 18748 23004 19288 23032
rect 18748 22992 18754 23004
rect 20070 22992 20076 23044
rect 20128 22992 20134 23044
rect 22830 22992 22836 23044
rect 22888 22992 22894 23044
rect 24946 23032 24952 23044
rect 23584 23004 24952 23032
rect 23584 22976 23612 23004
rect 24946 22992 24952 23004
rect 25004 23032 25010 23044
rect 25317 23035 25375 23041
rect 25317 23032 25329 23035
rect 25004 23004 25329 23032
rect 25004 22992 25010 23004
rect 25317 23001 25329 23004
rect 25363 23001 25375 23035
rect 25317 22995 25375 23001
rect 26970 22992 26976 23044
rect 27028 22992 27034 23044
rect 27798 22992 27804 23044
rect 27856 23032 27862 23044
rect 28537 23035 28595 23041
rect 28537 23032 28549 23035
rect 27856 23004 28549 23032
rect 27856 22992 27862 23004
rect 28537 23001 28549 23004
rect 28583 23032 28595 23035
rect 29270 23032 29276 23044
rect 28583 23004 29276 23032
rect 28583 23001 28595 23004
rect 28537 22995 28595 23001
rect 29270 22992 29276 23004
rect 29328 22992 29334 23044
rect 16666 22964 16672 22976
rect 15580 22936 16672 22964
rect 14645 22927 14703 22933
rect 16666 22924 16672 22936
rect 16724 22964 16730 22976
rect 17310 22964 17316 22976
rect 16724 22936 17316 22964
rect 16724 22924 16730 22936
rect 17310 22924 17316 22936
rect 17368 22924 17374 22976
rect 19150 22924 19156 22976
rect 19208 22964 19214 22976
rect 20993 22967 21051 22973
rect 20993 22964 21005 22967
rect 19208 22936 21005 22964
rect 19208 22924 19214 22936
rect 20993 22933 21005 22936
rect 21039 22933 21051 22967
rect 23566 22964 23572 22976
rect 23479 22936 23572 22964
rect 20993 22927 21051 22933
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 24486 22924 24492 22976
rect 24544 22964 24550 22976
rect 25517 22967 25575 22973
rect 25517 22964 25529 22967
rect 24544 22936 25529 22964
rect 24544 22924 24550 22936
rect 25517 22933 25529 22936
rect 25563 22933 25575 22967
rect 25517 22927 25575 22933
rect 25682 22924 25688 22976
rect 25740 22964 25746 22976
rect 27338 22964 27344 22976
rect 25740 22936 27344 22964
rect 25740 22924 25746 22936
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 27430 22924 27436 22976
rect 27488 22964 27494 22976
rect 27985 22967 28043 22973
rect 27985 22964 27997 22967
rect 27488 22936 27997 22964
rect 27488 22924 27494 22936
rect 27985 22933 27997 22936
rect 28031 22933 28043 22967
rect 27985 22927 28043 22933
rect 28442 22924 28448 22976
rect 28500 22964 28506 22976
rect 28737 22967 28795 22973
rect 28737 22964 28749 22967
rect 28500 22936 28749 22964
rect 28500 22924 28506 22936
rect 28737 22933 28749 22936
rect 28783 22933 28795 22967
rect 29380 22964 29408 23072
rect 29638 23060 29644 23112
rect 29696 23100 29702 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29696 23072 29745 23100
rect 29696 23060 29702 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 30098 23060 30104 23112
rect 30156 23100 30162 23112
rect 30377 23103 30435 23109
rect 30377 23100 30389 23103
rect 30156 23072 30389 23100
rect 30156 23060 30162 23072
rect 30377 23069 30389 23072
rect 30423 23069 30435 23103
rect 30377 23063 30435 23069
rect 31754 23060 31760 23112
rect 31812 23060 31818 23112
rect 33962 23100 33968 23112
rect 33923 23072 33968 23100
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 34701 23103 34759 23109
rect 34701 23069 34713 23103
rect 34747 23069 34759 23103
rect 34701 23063 34759 23069
rect 40313 23103 40371 23109
rect 40313 23069 40325 23103
rect 40359 23100 40371 23103
rect 41414 23100 41420 23112
rect 40359 23072 41420 23100
rect 40359 23069 40371 23072
rect 40313 23063 40371 23069
rect 33229 23035 33287 23041
rect 33229 23032 33241 23035
rect 32048 23004 33241 23032
rect 32048 22964 32076 23004
rect 33229 23001 33241 23004
rect 33275 23032 33287 23035
rect 33502 23032 33508 23044
rect 33275 23004 33508 23032
rect 33275 23001 33287 23004
rect 33229 22995 33287 23001
rect 33502 22992 33508 23004
rect 33560 22992 33566 23044
rect 34716 23032 34744 23063
rect 41414 23060 41420 23072
rect 41472 23060 41478 23112
rect 35526 23032 35532 23044
rect 34716 23004 35532 23032
rect 35526 22992 35532 23004
rect 35584 23032 35590 23044
rect 41524 23041 41552 23140
rect 42337 23103 42395 23109
rect 42337 23100 42349 23103
rect 41616 23072 42349 23100
rect 41509 23035 41567 23041
rect 41509 23032 41521 23035
rect 35584 23004 41521 23032
rect 35584 22992 35590 23004
rect 41509 23001 41521 23004
rect 41555 23001 41567 23035
rect 41509 22995 41567 23001
rect 29380 22936 32076 22964
rect 33520 22964 33548 22992
rect 41616 22976 41644 23072
rect 42337 23069 42349 23072
rect 42383 23069 42395 23103
rect 42337 23063 42395 23069
rect 42444 23032 42472 23140
rect 42613 23137 42625 23171
rect 42659 23168 42671 23171
rect 42659 23140 45554 23168
rect 42659 23137 42671 23140
rect 42613 23131 42671 23137
rect 43254 23100 43260 23112
rect 43215 23072 43260 23100
rect 43254 23060 43260 23072
rect 43312 23060 43318 23112
rect 43438 23100 43444 23112
rect 43399 23072 43444 23100
rect 43438 23060 43444 23072
rect 43496 23060 43502 23112
rect 44450 23100 44456 23112
rect 44411 23072 44456 23100
rect 44450 23060 44456 23072
rect 44508 23060 44514 23112
rect 45097 23035 45155 23041
rect 45097 23032 45109 23035
rect 42444 23004 45109 23032
rect 45097 23001 45109 23004
rect 45143 23001 45155 23035
rect 45278 23032 45284 23044
rect 45239 23004 45284 23032
rect 45097 22995 45155 23001
rect 34885 22967 34943 22973
rect 34885 22964 34897 22967
rect 33520 22936 34897 22964
rect 28737 22927 28795 22933
rect 34885 22933 34897 22936
rect 34931 22933 34943 22967
rect 41598 22964 41604 22976
rect 41559 22936 41604 22964
rect 34885 22927 34943 22933
rect 41598 22924 41604 22936
rect 41656 22924 41662 22976
rect 45112 22964 45140 22995
rect 45278 22992 45284 23004
rect 45336 22992 45342 23044
rect 45526 23032 45554 23140
rect 45646 23128 45652 23180
rect 45704 23168 45710 23180
rect 45940 23177 45968 23208
rect 45741 23171 45799 23177
rect 45741 23168 45753 23171
rect 45704 23140 45753 23168
rect 45704 23128 45710 23140
rect 45741 23137 45753 23140
rect 45787 23137 45799 23171
rect 45741 23131 45799 23137
rect 45925 23171 45983 23177
rect 45925 23137 45937 23171
rect 45971 23137 45983 23171
rect 46934 23168 46940 23180
rect 46895 23140 46940 23168
rect 45925 23131 45983 23137
rect 46934 23128 46940 23140
rect 46992 23128 46998 23180
rect 47486 23032 47492 23044
rect 45526 23004 47492 23032
rect 47486 22992 47492 23004
rect 47544 22992 47550 23044
rect 46566 22964 46572 22976
rect 45112 22936 46572 22964
rect 46566 22924 46572 22936
rect 46624 22924 46630 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 9582 22760 9588 22772
rect 9543 22732 9588 22760
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 13906 22760 13912 22772
rect 13867 22732 13912 22760
rect 13906 22720 13912 22732
rect 13964 22720 13970 22772
rect 21085 22763 21143 22769
rect 16546 22732 20944 22760
rect 11698 22692 11704 22704
rect 11659 22664 11704 22692
rect 11698 22652 11704 22664
rect 11756 22652 11762 22704
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 10134 22624 10140 22636
rect 9815 22596 10140 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 10778 22584 10784 22636
rect 10836 22624 10842 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10836 22596 11529 22624
rect 10836 22584 10842 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 11517 22587 11575 22593
rect 12912 22596 13829 22624
rect 11330 22448 11336 22500
rect 11388 22488 11394 22500
rect 12912 22488 12940 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 13354 22556 13360 22568
rect 13315 22528 13360 22556
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 11388 22460 12940 22488
rect 13832 22488 13860 22587
rect 14918 22584 14924 22636
rect 14976 22624 14982 22636
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14976 22596 15025 22624
rect 14976 22584 14982 22596
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 15013 22587 15071 22593
rect 15102 22584 15108 22636
rect 15160 22624 15166 22636
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 15160 22596 15853 22624
rect 15160 22584 15166 22596
rect 15841 22593 15853 22596
rect 15887 22624 15899 22627
rect 16546 22624 16574 22732
rect 18598 22692 18604 22704
rect 18446 22664 18604 22692
rect 18598 22652 18604 22664
rect 18656 22652 18662 22704
rect 19150 22624 19156 22636
rect 15887 22596 16574 22624
rect 19111 22596 19156 22624
rect 15887 22593 15899 22596
rect 15841 22587 15899 22593
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19886 22624 19892 22636
rect 19847 22596 19892 22624
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 20916 22633 20944 22732
rect 21085 22729 21097 22763
rect 21131 22729 21143 22763
rect 21085 22723 21143 22729
rect 21100 22692 21128 22723
rect 21818 22720 21824 22772
rect 21876 22760 21882 22772
rect 22005 22763 22063 22769
rect 22005 22760 22017 22763
rect 21876 22732 22017 22760
rect 21876 22720 21882 22732
rect 22005 22729 22017 22732
rect 22051 22729 22063 22763
rect 22830 22760 22836 22772
rect 22791 22732 22836 22760
rect 22005 22723 22063 22729
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 23382 22760 23388 22772
rect 23343 22732 23388 22760
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 23845 22763 23903 22769
rect 23845 22729 23857 22763
rect 23891 22729 23903 22763
rect 23845 22723 23903 22729
rect 23937 22763 23995 22769
rect 23937 22729 23949 22763
rect 23983 22760 23995 22763
rect 24854 22760 24860 22772
rect 23983 22732 24860 22760
rect 23983 22729 23995 22732
rect 23937 22723 23995 22729
rect 23860 22692 23888 22723
rect 24854 22720 24860 22732
rect 24912 22720 24918 22772
rect 26329 22763 26387 22769
rect 26329 22729 26341 22763
rect 26375 22760 26387 22763
rect 26970 22760 26976 22772
rect 26375 22732 26976 22760
rect 26375 22729 26387 22732
rect 26329 22723 26387 22729
rect 26970 22720 26976 22732
rect 27028 22720 27034 22772
rect 27255 22763 27313 22769
rect 27255 22729 27267 22763
rect 27301 22729 27313 22763
rect 27255 22723 27313 22729
rect 24486 22692 24492 22704
rect 21100 22664 22094 22692
rect 23860 22664 24492 22692
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22593 20959 22627
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 20901 22587 20959 22593
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22066 22624 22094 22664
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 24719 22661 24777 22667
rect 24719 22658 24731 22661
rect 22278 22624 22284 22636
rect 22066 22596 22284 22624
rect 22278 22584 22284 22596
rect 22336 22624 22342 22636
rect 22741 22627 22799 22633
rect 22741 22624 22753 22627
rect 22336 22596 22753 22624
rect 22336 22584 22342 22596
rect 22741 22593 22753 22596
rect 22787 22624 22799 22627
rect 22830 22624 22836 22636
rect 22787 22596 22836 22624
rect 22787 22593 22799 22596
rect 22741 22587 22799 22593
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 23566 22624 23572 22636
rect 23527 22596 23572 22624
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 23842 22584 23848 22636
rect 23900 22624 23906 22636
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23900 22596 24041 22624
rect 23900 22584 23906 22596
rect 24029 22593 24041 22596
rect 24075 22624 24087 22627
rect 24704 22627 24731 22658
rect 24765 22627 24777 22661
rect 26878 22652 26884 22704
rect 26936 22692 26942 22704
rect 27270 22692 27298 22723
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 29178 22760 29184 22772
rect 27488 22732 27533 22760
rect 29139 22732 29184 22760
rect 27488 22720 27494 22732
rect 29178 22720 29184 22732
rect 29236 22720 29242 22772
rect 30098 22760 30104 22772
rect 30059 22732 30104 22760
rect 30098 22720 30104 22732
rect 30156 22720 30162 22772
rect 40218 22720 40224 22772
rect 40276 22760 40282 22772
rect 40865 22763 40923 22769
rect 40865 22760 40877 22763
rect 40276 22732 40877 22760
rect 40276 22720 40282 22732
rect 40865 22729 40877 22732
rect 40911 22729 40923 22763
rect 43070 22760 43076 22772
rect 43031 22732 43076 22760
rect 40865 22723 40923 22729
rect 43070 22720 43076 22732
rect 43128 22720 43134 22772
rect 44450 22720 44456 22772
rect 44508 22760 44514 22772
rect 48133 22763 48191 22769
rect 48133 22760 48145 22763
rect 44508 22732 48145 22760
rect 44508 22720 44514 22732
rect 48133 22729 48145 22732
rect 48179 22729 48191 22763
rect 48133 22723 48191 22729
rect 26936 22664 27298 22692
rect 26936 22652 26942 22664
rect 28902 22652 28908 22704
rect 28960 22692 28966 22704
rect 45373 22695 45431 22701
rect 28960 22664 29316 22692
rect 28960 22652 28966 22664
rect 24704 22624 24777 22627
rect 25498 22624 25504 22636
rect 24075 22621 24777 22624
rect 24075 22596 24732 22621
rect 25459 22596 25504 22624
rect 24075 22593 24087 22596
rect 24029 22587 24087 22593
rect 24688 22568 24716 22596
rect 25498 22584 25504 22596
rect 25556 22584 25562 22636
rect 25682 22624 25688 22636
rect 25643 22596 25688 22624
rect 25682 22584 25688 22596
rect 25740 22584 25746 22636
rect 26237 22627 26295 22633
rect 26237 22593 26249 22627
rect 26283 22624 26295 22627
rect 26510 22624 26516 22636
rect 26283 22596 26516 22624
rect 26283 22593 26295 22596
rect 26237 22587 26295 22593
rect 26510 22584 26516 22596
rect 26568 22624 26574 22636
rect 27154 22624 27160 22636
rect 26568 22596 27160 22624
rect 26568 22584 26574 22596
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 27270 22596 27353 22624
rect 16942 22556 16948 22568
rect 16903 22528 16948 22556
rect 16942 22516 16948 22528
rect 17000 22516 17006 22568
rect 17218 22556 17224 22568
rect 17179 22528 17224 22556
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 23661 22559 23719 22565
rect 23661 22525 23673 22559
rect 23707 22525 23719 22559
rect 23661 22519 23719 22525
rect 15194 22488 15200 22500
rect 13832 22460 15200 22488
rect 11388 22448 11394 22460
rect 15194 22448 15200 22460
rect 15252 22448 15258 22500
rect 15378 22448 15384 22500
rect 15436 22488 15442 22500
rect 19337 22491 19395 22497
rect 15436 22460 16574 22488
rect 15436 22448 15442 22460
rect 16546 22432 16574 22460
rect 19337 22457 19349 22491
rect 19383 22488 19395 22491
rect 21818 22488 21824 22500
rect 19383 22460 21824 22488
rect 19383 22457 19395 22460
rect 19337 22451 19395 22457
rect 21818 22448 21824 22460
rect 21876 22448 21882 22500
rect 22738 22448 22744 22500
rect 22796 22488 22802 22500
rect 23676 22488 23704 22519
rect 24670 22516 24676 22568
rect 24728 22516 24734 22568
rect 25774 22556 25780 22568
rect 25735 22528 25780 22556
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 27062 22516 27068 22568
rect 27120 22556 27126 22568
rect 27270 22556 27298 22596
rect 27341 22593 27353 22596
rect 27387 22593 27399 22627
rect 29086 22624 29092 22636
rect 29047 22596 29092 22624
rect 27341 22587 27399 22593
rect 29086 22584 29092 22596
rect 29144 22584 29150 22636
rect 29288 22633 29316 22664
rect 45373 22661 45385 22695
rect 45419 22692 45431 22695
rect 45554 22692 45560 22704
rect 45419 22664 45560 22692
rect 45419 22661 45431 22664
rect 45373 22655 45431 22661
rect 45554 22652 45560 22664
rect 45612 22652 45618 22704
rect 29273 22627 29331 22633
rect 29273 22593 29285 22627
rect 29319 22593 29331 22627
rect 29273 22587 29331 22593
rect 29822 22584 29828 22636
rect 29880 22624 29886 22636
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29880 22596 29929 22624
rect 29880 22584 29886 22596
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 39945 22627 40003 22633
rect 39945 22593 39957 22627
rect 39991 22624 40003 22627
rect 40218 22624 40224 22636
rect 39991 22596 40224 22624
rect 39991 22593 40003 22596
rect 39945 22587 40003 22593
rect 40218 22584 40224 22596
rect 40276 22584 40282 22636
rect 41049 22627 41107 22633
rect 41049 22624 41061 22627
rect 40420 22596 41061 22624
rect 27706 22556 27712 22568
rect 27120 22528 27298 22556
rect 27667 22528 27712 22556
rect 27120 22516 27126 22528
rect 27706 22516 27712 22528
rect 27764 22516 27770 22568
rect 40420 22565 40448 22596
rect 41049 22593 41061 22596
rect 41095 22593 41107 22627
rect 41049 22587 41107 22593
rect 42981 22627 43039 22633
rect 42981 22593 42993 22627
rect 43027 22593 43039 22627
rect 42981 22587 43039 22593
rect 43165 22627 43223 22633
rect 43165 22593 43177 22627
rect 43211 22624 43223 22627
rect 43438 22624 43444 22636
rect 43211 22596 43444 22624
rect 43211 22593 43223 22596
rect 43165 22587 43223 22593
rect 40405 22559 40463 22565
rect 40405 22525 40417 22559
rect 40451 22525 40463 22559
rect 42996 22556 43024 22587
rect 43438 22584 43444 22596
rect 43496 22584 43502 22636
rect 45094 22584 45100 22636
rect 45152 22624 45158 22636
rect 45189 22627 45247 22633
rect 45189 22624 45201 22627
rect 45152 22596 45201 22624
rect 45152 22584 45158 22596
rect 45189 22593 45201 22596
rect 45235 22593 45247 22627
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 45189 22587 45247 22593
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 43254 22556 43260 22568
rect 42996 22528 43260 22556
rect 40405 22519 40463 22525
rect 43254 22516 43260 22528
rect 43312 22556 43318 22568
rect 43714 22556 43720 22568
rect 43312 22528 43720 22556
rect 43312 22516 43318 22528
rect 43714 22516 43720 22528
rect 43772 22516 43778 22568
rect 43901 22559 43959 22565
rect 43901 22525 43913 22559
rect 43947 22525 43959 22559
rect 44174 22556 44180 22568
rect 44135 22528 44180 22556
rect 43901 22519 43959 22525
rect 25038 22488 25044 22500
rect 22796 22460 25044 22488
rect 22796 22448 22802 22460
rect 25038 22448 25044 22460
rect 25096 22448 25102 22500
rect 25317 22491 25375 22497
rect 25317 22457 25329 22491
rect 25363 22488 25375 22491
rect 25866 22488 25872 22500
rect 25363 22460 25872 22488
rect 25363 22457 25375 22460
rect 25317 22451 25375 22457
rect 25866 22448 25872 22460
rect 25924 22448 25930 22500
rect 26142 22448 26148 22500
rect 26200 22488 26206 22500
rect 41598 22488 41604 22500
rect 26200 22460 41604 22488
rect 26200 22448 26206 22460
rect 41598 22448 41604 22460
rect 41656 22448 41662 22500
rect 43916 22488 43944 22519
rect 44174 22516 44180 22528
rect 44232 22516 44238 22568
rect 46934 22556 46940 22568
rect 46895 22528 46940 22556
rect 46934 22516 46940 22528
rect 46992 22516 46998 22568
rect 47854 22556 47860 22568
rect 47815 22528 47860 22556
rect 47854 22516 47860 22528
rect 47912 22516 47918 22568
rect 46842 22488 46848 22500
rect 43916 22460 46848 22488
rect 46842 22448 46848 22460
rect 46900 22448 46906 22500
rect 16025 22423 16083 22429
rect 16025 22389 16037 22423
rect 16071 22420 16083 22423
rect 16298 22420 16304 22432
rect 16071 22392 16304 22420
rect 16071 22389 16083 22392
rect 16025 22383 16083 22389
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16482 22380 16488 22432
rect 16540 22420 16574 22432
rect 18693 22423 18751 22429
rect 18693 22420 18705 22423
rect 16540 22392 18705 22420
rect 16540 22380 16546 22392
rect 18693 22389 18705 22392
rect 18739 22389 18751 22423
rect 18693 22383 18751 22389
rect 20073 22423 20131 22429
rect 20073 22389 20085 22423
rect 20119 22420 20131 22423
rect 20162 22420 20168 22432
rect 20119 22392 20168 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20162 22380 20168 22392
rect 20220 22380 20226 22432
rect 24394 22380 24400 22432
rect 24452 22420 24458 22432
rect 24673 22423 24731 22429
rect 24673 22420 24685 22423
rect 24452 22392 24685 22420
rect 24452 22380 24458 22392
rect 24673 22389 24685 22392
rect 24719 22389 24731 22423
rect 24673 22383 24731 22389
rect 24762 22380 24768 22432
rect 24820 22420 24826 22432
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 24820 22392 24869 22420
rect 24820 22380 24826 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 26973 22423 27031 22429
rect 26973 22389 26985 22423
rect 27019 22420 27031 22423
rect 27246 22420 27252 22432
rect 27019 22392 27252 22420
rect 27019 22389 27031 22392
rect 26973 22383 27031 22389
rect 27246 22380 27252 22392
rect 27304 22380 27310 22432
rect 27338 22380 27344 22432
rect 27396 22420 27402 22432
rect 27617 22423 27675 22429
rect 27617 22420 27629 22423
rect 27396 22392 27629 22420
rect 27396 22380 27402 22392
rect 27617 22389 27629 22392
rect 27663 22389 27675 22423
rect 40034 22420 40040 22432
rect 39995 22392 40040 22420
rect 27617 22383 27675 22389
rect 40034 22380 40040 22392
rect 40092 22380 40098 22432
rect 41874 22380 41880 22432
rect 41932 22420 41938 22432
rect 46934 22420 46940 22432
rect 41932 22392 46940 22420
rect 41932 22380 41938 22392
rect 46934 22380 46940 22392
rect 46992 22380 46998 22432
rect 47670 22420 47676 22432
rect 47631 22392 47676 22420
rect 47670 22380 47676 22392
rect 47728 22380 47734 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 15473 22219 15531 22225
rect 15473 22185 15485 22219
rect 15519 22216 15531 22219
rect 15930 22216 15936 22228
rect 15519 22188 15936 22216
rect 15519 22185 15531 22188
rect 15473 22179 15531 22185
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 16853 22219 16911 22225
rect 16853 22185 16865 22219
rect 16899 22216 16911 22219
rect 17218 22216 17224 22228
rect 16899 22188 17224 22216
rect 16899 22185 16911 22188
rect 16853 22179 16911 22185
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 19886 22176 19892 22228
rect 19944 22216 19950 22228
rect 26142 22216 26148 22228
rect 19944 22188 26148 22216
rect 19944 22176 19950 22188
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 26329 22219 26387 22225
rect 26329 22216 26341 22219
rect 26292 22188 26341 22216
rect 26292 22176 26298 22188
rect 26329 22185 26341 22188
rect 26375 22185 26387 22219
rect 26329 22179 26387 22185
rect 27062 22176 27068 22228
rect 27120 22216 27126 22228
rect 27522 22216 27528 22228
rect 27120 22188 27528 22216
rect 27120 22176 27126 22188
rect 27522 22176 27528 22188
rect 27580 22176 27586 22228
rect 27709 22219 27767 22225
rect 27709 22185 27721 22219
rect 27755 22216 27767 22219
rect 28810 22216 28816 22228
rect 27755 22188 28816 22216
rect 27755 22185 27767 22188
rect 27709 22179 27767 22185
rect 28810 22176 28816 22188
rect 28868 22176 28874 22228
rect 29917 22219 29975 22225
rect 29917 22185 29929 22219
rect 29963 22216 29975 22219
rect 30006 22216 30012 22228
rect 29963 22188 30012 22216
rect 29963 22185 29975 22188
rect 29917 22179 29975 22185
rect 30006 22176 30012 22188
rect 30064 22176 30070 22228
rect 13078 22108 13084 22160
rect 13136 22108 13142 22160
rect 17494 22148 17500 22160
rect 17407 22120 17500 22148
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 11882 22080 11888 22092
rect 9631 22052 11888 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 13096 22080 13124 22108
rect 12452 22052 13124 22080
rect 13740 22052 14412 22080
rect 12452 22024 12480 22052
rect 12434 22012 12440 22024
rect 12347 21984 12440 22012
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12584 21984 13093 22012
rect 12584 21972 12590 21984
rect 13081 21981 13093 21984
rect 13127 22012 13139 22015
rect 13740 22012 13768 22052
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13127 21984 13768 22012
rect 13832 21984 14105 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 9769 21947 9827 21953
rect 9769 21913 9781 21947
rect 9815 21944 9827 21947
rect 9950 21944 9956 21956
rect 9815 21916 9956 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 9950 21904 9956 21916
rect 10008 21904 10014 21956
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 11425 21947 11483 21953
rect 11425 21944 11437 21947
rect 11112 21916 11437 21944
rect 11112 21904 11118 21916
rect 11425 21913 11437 21916
rect 11471 21913 11483 21947
rect 11425 21907 11483 21913
rect 13832 21888 13860 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 12526 21876 12532 21888
rect 12487 21848 12532 21876
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 13814 21876 13820 21888
rect 13311 21848 13820 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14274 21876 14280 21888
rect 14235 21848 14280 21876
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 14384 21876 14412 22052
rect 16574 22040 16580 22092
rect 16632 22080 16638 22092
rect 16632 22052 16677 22080
rect 16632 22040 16638 22052
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 15252 21984 15393 22012
rect 15252 21972 15258 21984
rect 15381 21981 15393 21984
rect 15427 21981 15439 22015
rect 16482 22012 16488 22024
rect 16443 21984 16488 22012
rect 15381 21975 15439 21981
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 17420 22021 17448 22120
rect 17494 22108 17500 22120
rect 17552 22148 17558 22160
rect 19904 22148 19932 22176
rect 26418 22148 26424 22160
rect 17552 22120 19932 22148
rect 21744 22120 26424 22148
rect 17552 22108 17558 22120
rect 18598 22080 18604 22092
rect 18559 22052 18604 22080
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 21744 22080 21772 22120
rect 26418 22108 26424 22120
rect 26476 22108 26482 22160
rect 27614 22108 27620 22160
rect 27672 22108 27678 22160
rect 19076 22052 21772 22080
rect 21821 22083 21879 22089
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 21981 17463 22015
rect 18509 22015 18567 22021
rect 18509 22012 18521 22015
rect 17405 21975 17463 21981
rect 17512 21984 18521 22012
rect 16298 21904 16304 21956
rect 16356 21944 16362 21956
rect 17512 21944 17540 21984
rect 18509 21981 18521 21984
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 16356 21916 17540 21944
rect 16356 21904 16362 21916
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 17865 21947 17923 21953
rect 17865 21944 17877 21947
rect 17736 21916 17877 21944
rect 17736 21904 17742 21916
rect 17865 21913 17877 21916
rect 17911 21944 17923 21947
rect 19076 21944 19104 22052
rect 21821 22049 21833 22083
rect 21867 22080 21879 22083
rect 27632 22080 27660 22108
rect 21867 22052 27660 22080
rect 28966 22052 29868 22080
rect 21867 22049 21879 22052
rect 21821 22043 21879 22049
rect 19150 21972 19156 22024
rect 19208 22012 19214 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19208 21984 19257 22012
rect 19208 21972 19214 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19978 22012 19984 22024
rect 19939 21984 19984 22012
rect 19245 21975 19303 21981
rect 17911 21916 19104 21944
rect 17911 21913 17923 21916
rect 17865 21907 17923 21913
rect 19260 21876 19288 21975
rect 19978 21972 19984 21984
rect 20036 21972 20042 22024
rect 23661 22015 23719 22021
rect 23661 21981 23673 22015
rect 23707 22012 23719 22015
rect 23750 22012 23756 22024
rect 23707 21984 23756 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 22012 23903 22015
rect 24670 22012 24676 22024
rect 23891 21984 24532 22012
rect 24631 21984 24676 22012
rect 23891 21981 23903 21984
rect 23845 21975 23903 21981
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21944 20223 21947
rect 20990 21944 20996 21956
rect 20211 21916 20996 21944
rect 20211 21913 20223 21916
rect 20165 21907 20223 21913
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 24210 21944 24216 21956
rect 23768 21916 24216 21944
rect 23768 21888 23796 21916
rect 24210 21904 24216 21916
rect 24268 21904 24274 21956
rect 24394 21944 24400 21956
rect 24355 21916 24400 21944
rect 24394 21904 24400 21916
rect 24452 21904 24458 21956
rect 24504 21944 24532 21984
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 26142 22012 26148 22024
rect 26103 21984 26148 22012
rect 26142 21972 26148 21984
rect 26200 21972 26206 22024
rect 26418 21972 26424 22024
rect 26476 22012 26482 22024
rect 28966 22012 28994 22052
rect 26476 21984 28994 22012
rect 26476 21972 26482 21984
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 29696 21984 29745 22012
rect 29696 21972 29702 21984
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 29840 22012 29868 22052
rect 31726 22052 41414 22080
rect 31726 22012 31754 22052
rect 29840 21984 31754 22012
rect 39945 22015 40003 22021
rect 29733 21975 29791 21981
rect 39945 21981 39957 22015
rect 39991 21981 40003 22015
rect 39945 21975 40003 21981
rect 24581 21947 24639 21953
rect 24581 21944 24593 21947
rect 24504 21916 24593 21944
rect 24581 21913 24593 21916
rect 24627 21944 24639 21947
rect 24854 21944 24860 21956
rect 24627 21916 24860 21944
rect 24627 21913 24639 21916
rect 24581 21907 24639 21913
rect 24854 21904 24860 21916
rect 24912 21904 24918 21956
rect 27430 21904 27436 21956
rect 27488 21944 27494 21956
rect 27525 21947 27583 21953
rect 27525 21944 27537 21947
rect 27488 21916 27537 21944
rect 27488 21904 27494 21916
rect 27525 21913 27537 21916
rect 27571 21913 27583 21947
rect 27525 21907 27583 21913
rect 27614 21904 27620 21956
rect 27672 21944 27678 21956
rect 37274 21944 37280 21956
rect 27672 21916 37280 21944
rect 27672 21904 27678 21916
rect 37274 21904 37280 21916
rect 37332 21904 37338 21956
rect 39960 21944 39988 21975
rect 40034 21972 40040 22024
rect 40092 22012 40098 22024
rect 40129 22015 40187 22021
rect 40129 22012 40141 22015
rect 40092 21984 40141 22012
rect 40092 21972 40098 21984
rect 40129 21981 40141 21984
rect 40175 21981 40187 22015
rect 40129 21975 40187 21981
rect 40218 21944 40224 21956
rect 39960 21916 40224 21944
rect 40218 21904 40224 21916
rect 40276 21904 40282 21956
rect 40313 21947 40371 21953
rect 40313 21913 40325 21947
rect 40359 21944 40371 21947
rect 40494 21944 40500 21956
rect 40359 21916 40500 21944
rect 40359 21913 40371 21916
rect 40313 21907 40371 21913
rect 40494 21904 40500 21916
rect 40552 21904 40558 21956
rect 41386 21944 41414 22052
rect 41690 22040 41696 22092
rect 41748 22080 41754 22092
rect 41748 22052 42656 22080
rect 41748 22040 41754 22052
rect 42518 22012 42524 22024
rect 42479 21984 42524 22012
rect 42518 21972 42524 21984
rect 42576 21972 42582 22024
rect 42628 22006 42656 22052
rect 45554 22040 45560 22092
rect 45612 22080 45618 22092
rect 47121 22083 47179 22089
rect 47121 22080 47133 22083
rect 45612 22052 47133 22080
rect 45612 22040 45618 22052
rect 47121 22049 47133 22052
rect 47167 22049 47179 22083
rect 47121 22043 47179 22049
rect 42705 22015 42763 22021
rect 42705 22006 42717 22015
rect 42628 21981 42717 22006
rect 42751 21981 42763 22015
rect 42628 21978 42763 21981
rect 42705 21975 42763 21978
rect 43809 22015 43867 22021
rect 43809 21981 43821 22015
rect 43855 22012 43867 22015
rect 44542 22012 44548 22024
rect 43855 21984 44548 22012
rect 43855 21981 43867 21984
rect 43809 21975 43867 21981
rect 44542 21972 44548 21984
rect 44600 22012 44606 22024
rect 45278 22012 45284 22024
rect 44600 21984 45284 22012
rect 44600 21972 44606 21984
rect 45278 21972 45284 21984
rect 45336 22012 45342 22024
rect 45373 22015 45431 22021
rect 45373 22012 45385 22015
rect 45336 21984 45385 22012
rect 45336 21972 45342 21984
rect 45373 21981 45385 21984
rect 45419 21981 45431 22015
rect 45373 21975 45431 21981
rect 46845 22015 46903 22021
rect 46845 21981 46857 22015
rect 46891 22012 46903 22015
rect 47026 22012 47032 22024
rect 46891 21984 47032 22012
rect 46891 21981 46903 21984
rect 46845 21975 46903 21981
rect 47026 21972 47032 21984
rect 47084 21972 47090 22024
rect 42242 21944 42248 21956
rect 41386 21916 42248 21944
rect 42242 21904 42248 21916
rect 42300 21904 42306 21956
rect 42426 21904 42432 21956
rect 42484 21944 42490 21956
rect 44174 21944 44180 21956
rect 42484 21916 44180 21944
rect 42484 21904 42490 21916
rect 44174 21904 44180 21916
rect 44232 21904 44238 21956
rect 44266 21904 44272 21956
rect 44324 21944 44330 21956
rect 45922 21944 45928 21956
rect 44324 21916 45928 21944
rect 44324 21904 44330 21916
rect 45922 21904 45928 21916
rect 45980 21904 45986 21956
rect 46014 21904 46020 21956
rect 46072 21944 46078 21956
rect 46201 21947 46259 21953
rect 46201 21944 46213 21947
rect 46072 21916 46213 21944
rect 46072 21904 46078 21916
rect 46201 21913 46213 21916
rect 46247 21913 46259 21947
rect 46201 21907 46259 21913
rect 14384 21848 19288 21876
rect 19429 21879 19487 21885
rect 19429 21845 19441 21879
rect 19475 21876 19487 21879
rect 20070 21876 20076 21888
rect 19475 21848 20076 21876
rect 19475 21845 19487 21848
rect 19429 21839 19487 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 23750 21876 23756 21888
rect 23711 21848 23756 21876
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 23842 21836 23848 21888
rect 23900 21876 23906 21888
rect 24495 21879 24553 21885
rect 24495 21876 24507 21879
rect 23900 21848 24507 21876
rect 23900 21836 23906 21848
rect 24495 21845 24507 21848
rect 24541 21845 24553 21879
rect 24495 21839 24553 21845
rect 27706 21836 27712 21888
rect 27764 21885 27770 21888
rect 27764 21879 27783 21885
rect 27771 21845 27783 21879
rect 27890 21876 27896 21888
rect 27851 21848 27896 21876
rect 27764 21839 27783 21845
rect 27764 21836 27770 21839
rect 27890 21836 27896 21848
rect 27948 21836 27954 21888
rect 42334 21836 42340 21888
rect 42392 21876 42398 21888
rect 42889 21879 42947 21885
rect 42889 21876 42901 21879
rect 42392 21848 42901 21876
rect 42392 21836 42398 21848
rect 42889 21845 42901 21848
rect 42935 21845 42947 21879
rect 42889 21839 42947 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 9950 21672 9956 21684
rect 9911 21644 9956 21672
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 11440 21644 27476 21672
rect 11330 21604 11336 21616
rect 9876 21576 11336 21604
rect 9876 21545 9904 21576
rect 11330 21564 11336 21576
rect 11388 21564 11394 21616
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 9263 21508 9873 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 10410 21496 10416 21548
rect 10468 21536 10474 21548
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 10468 21508 10701 21536
rect 10468 21496 10474 21508
rect 10689 21505 10701 21508
rect 10735 21505 10747 21539
rect 11440 21536 11468 21644
rect 12526 21564 12532 21616
rect 12584 21564 12590 21616
rect 16942 21564 16948 21616
rect 17000 21604 17006 21616
rect 17497 21607 17555 21613
rect 17497 21604 17509 21607
rect 17000 21576 17509 21604
rect 17000 21564 17006 21576
rect 17497 21573 17509 21576
rect 17543 21573 17555 21607
rect 20990 21604 20996 21616
rect 20951 21576 20996 21604
rect 17497 21567 17555 21573
rect 20990 21564 20996 21576
rect 21048 21564 21054 21616
rect 23842 21604 23848 21616
rect 23584 21576 23848 21604
rect 14274 21536 14280 21548
rect 10689 21499 10747 21505
rect 10796 21508 11468 21536
rect 14235 21508 14280 21536
rect 2866 21428 2872 21480
rect 2924 21468 2930 21480
rect 10796 21468 10824 21508
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 15654 21496 15660 21548
rect 15712 21496 15718 21548
rect 17405 21539 17463 21545
rect 17405 21505 17417 21539
rect 17451 21536 17463 21539
rect 20070 21536 20076 21548
rect 17451 21508 20076 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21505 20959 21539
rect 21818 21536 21824 21548
rect 21779 21508 21824 21536
rect 20901 21499 20959 21505
rect 2924 21440 10824 21468
rect 10965 21471 11023 21477
rect 2924 21428 2930 21440
rect 10965 21437 10977 21471
rect 11011 21468 11023 21471
rect 11609 21471 11667 21477
rect 11609 21468 11621 21471
rect 11011 21440 11621 21468
rect 11011 21437 11023 21440
rect 10965 21431 11023 21437
rect 11609 21437 11621 21440
rect 11655 21437 11667 21471
rect 11882 21468 11888 21480
rect 11843 21440 11888 21468
rect 11609 21431 11667 21437
rect 11882 21428 11888 21440
rect 11940 21428 11946 21480
rect 11974 21428 11980 21480
rect 12032 21468 12038 21480
rect 14550 21468 14556 21480
rect 12032 21440 13400 21468
rect 14511 21440 14556 21468
rect 12032 21428 12038 21440
rect 9306 21332 9312 21344
rect 9267 21304 9312 21332
rect 9306 21292 9312 21304
rect 9364 21292 9370 21344
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 12526 21332 12532 21344
rect 9640 21304 12532 21332
rect 9640 21292 9646 21304
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13372 21341 13400 21440
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 20162 21468 20168 21480
rect 19484 21440 20168 21468
rect 19484 21428 19490 21440
rect 20162 21428 20168 21440
rect 20220 21468 20226 21480
rect 20916 21468 20944 21499
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22738 21536 22744 21548
rect 22699 21508 22744 21536
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23584 21545 23612 21576
rect 23842 21564 23848 21576
rect 23900 21564 23906 21616
rect 26970 21564 26976 21616
rect 27028 21604 27034 21616
rect 27341 21607 27399 21613
rect 27341 21604 27353 21607
rect 27028 21576 27353 21604
rect 27028 21564 27034 21576
rect 27341 21573 27353 21576
rect 27387 21573 27399 21607
rect 27448 21604 27476 21644
rect 27522 21632 27528 21684
rect 27580 21681 27586 21684
rect 27580 21675 27599 21681
rect 27587 21641 27599 21675
rect 27706 21672 27712 21684
rect 27667 21644 27712 21672
rect 27580 21635 27599 21641
rect 27580 21632 27586 21635
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 42426 21672 42432 21684
rect 30944 21644 42432 21672
rect 30944 21613 30972 21644
rect 42426 21632 42432 21644
rect 42484 21632 42490 21684
rect 42797 21675 42855 21681
rect 42797 21641 42809 21675
rect 42843 21672 42855 21675
rect 43162 21672 43168 21684
rect 42843 21644 43168 21672
rect 42843 21641 42855 21644
rect 42797 21635 42855 21641
rect 43162 21632 43168 21644
rect 43220 21632 43226 21684
rect 47486 21632 47492 21684
rect 47544 21672 47550 21684
rect 47765 21675 47823 21681
rect 47765 21672 47777 21675
rect 47544 21644 47777 21672
rect 47544 21632 47550 21644
rect 47765 21641 47777 21644
rect 47811 21641 47823 21675
rect 47765 21635 47823 21641
rect 30929 21607 30987 21613
rect 27448 21576 30144 21604
rect 27341 21567 27399 21573
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21505 23627 21539
rect 23569 21499 23627 21505
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21536 23811 21539
rect 24762 21536 24768 21548
rect 23799 21508 24768 21536
rect 23799 21505 23811 21508
rect 23753 21499 23811 21505
rect 20220 21440 20944 21468
rect 22833 21471 22891 21477
rect 20220 21428 20226 21440
rect 22833 21437 22845 21471
rect 22879 21468 22891 21471
rect 23768 21468 23796 21499
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 26142 21536 26148 21548
rect 25976 21508 26148 21536
rect 22879 21440 23796 21468
rect 22879 21437 22891 21440
rect 22833 21431 22891 21437
rect 20346 21400 20352 21412
rect 20259 21372 20352 21400
rect 20346 21360 20352 21372
rect 20404 21400 20410 21412
rect 25976 21400 26004 21508
rect 26142 21496 26148 21508
rect 26200 21536 26206 21548
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 26200 21508 26249 21536
rect 26200 21496 26206 21508
rect 26237 21505 26249 21508
rect 26283 21536 26295 21539
rect 29638 21536 29644 21548
rect 26283 21508 29644 21536
rect 26283 21505 26295 21508
rect 26237 21499 26295 21505
rect 29638 21496 29644 21508
rect 29696 21536 29702 21548
rect 29822 21536 29828 21548
rect 29696 21508 29828 21536
rect 29696 21496 29702 21508
rect 29822 21496 29828 21508
rect 29880 21496 29886 21548
rect 20404 21372 26004 21400
rect 20404 21360 20410 21372
rect 26050 21360 26056 21412
rect 26108 21400 26114 21412
rect 29822 21400 29828 21412
rect 26108 21372 29828 21400
rect 26108 21360 26114 21372
rect 29822 21360 29828 21372
rect 29880 21360 29886 21412
rect 13357 21335 13415 21341
rect 13357 21301 13369 21335
rect 13403 21332 13415 21335
rect 14734 21332 14740 21344
rect 13403 21304 14740 21332
rect 13403 21301 13415 21304
rect 13357 21295 13415 21301
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 16022 21332 16028 21344
rect 15935 21304 16028 21332
rect 16022 21292 16028 21304
rect 16080 21332 16086 21344
rect 19978 21332 19984 21344
rect 16080 21304 19984 21332
rect 16080 21292 16086 21304
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 21082 21292 21088 21344
rect 21140 21332 21146 21344
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21140 21304 21925 21332
rect 21140 21292 21146 21304
rect 21913 21301 21925 21304
rect 21959 21301 21971 21335
rect 23106 21332 23112 21344
rect 23067 21304 23112 21332
rect 21913 21295 21971 21301
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 23569 21335 23627 21341
rect 23569 21332 23581 21335
rect 23532 21304 23581 21332
rect 23532 21292 23538 21304
rect 23569 21301 23581 21304
rect 23615 21301 23627 21335
rect 23569 21295 23627 21301
rect 26329 21335 26387 21341
rect 26329 21301 26341 21335
rect 26375 21332 26387 21335
rect 26878 21332 26884 21344
rect 26375 21304 26884 21332
rect 26375 21301 26387 21304
rect 26329 21295 26387 21301
rect 26878 21292 26884 21304
rect 26936 21292 26942 21344
rect 27522 21332 27528 21344
rect 27483 21304 27528 21332
rect 27522 21292 27528 21304
rect 27580 21292 27586 21344
rect 30116 21332 30144 21576
rect 30929 21573 30941 21607
rect 30975 21573 30987 21607
rect 30929 21567 30987 21573
rect 31021 21607 31079 21613
rect 31021 21573 31033 21607
rect 31067 21604 31079 21607
rect 32030 21604 32036 21616
rect 31067 21576 32036 21604
rect 31067 21573 31079 21576
rect 31021 21567 31079 21573
rect 32030 21564 32036 21576
rect 32088 21564 32094 21616
rect 41785 21607 41843 21613
rect 41785 21573 41797 21607
rect 41831 21604 41843 21607
rect 45738 21604 45744 21616
rect 41831 21576 43208 21604
rect 41831 21573 41843 21576
rect 41785 21567 41843 21573
rect 41690 21536 41696 21548
rect 41651 21508 41696 21536
rect 41690 21496 41696 21508
rect 41748 21496 41754 21548
rect 41877 21539 41935 21545
rect 41877 21505 41889 21539
rect 41923 21536 41935 21539
rect 42518 21536 42524 21548
rect 41923 21508 42524 21536
rect 41923 21505 41935 21508
rect 41877 21499 41935 21505
rect 42518 21496 42524 21508
rect 42576 21496 42582 21548
rect 42702 21496 42708 21548
rect 42760 21536 42766 21548
rect 43180 21545 43208 21576
rect 44008 21576 45744 21604
rect 42981 21539 43039 21545
rect 42981 21536 42993 21539
rect 42760 21508 42993 21536
rect 42760 21496 42766 21508
rect 42981 21505 42993 21508
rect 43027 21505 43039 21539
rect 42981 21499 43039 21505
rect 43165 21539 43223 21545
rect 43165 21505 43177 21539
rect 43211 21505 43223 21539
rect 43165 21499 43223 21505
rect 43254 21496 43260 21548
rect 43312 21536 43318 21548
rect 44008 21545 44036 21576
rect 45738 21564 45744 21576
rect 45796 21564 45802 21616
rect 47210 21564 47216 21616
rect 47268 21604 47274 21616
rect 47581 21607 47639 21613
rect 47581 21604 47593 21607
rect 47268 21576 47593 21604
rect 47268 21564 47274 21576
rect 47581 21573 47593 21576
rect 47627 21573 47639 21607
rect 47581 21567 47639 21573
rect 43993 21539 44051 21545
rect 43312 21508 43357 21536
rect 43312 21496 43318 21508
rect 43993 21505 44005 21539
rect 44039 21505 44051 21539
rect 44542 21536 44548 21548
rect 44503 21508 44548 21536
rect 43993 21499 44051 21505
rect 44542 21496 44548 21508
rect 44600 21536 44606 21548
rect 45370 21536 45376 21548
rect 44600 21508 45376 21536
rect 44600 21496 44606 21508
rect 45370 21496 45376 21508
rect 45428 21536 45434 21548
rect 45465 21539 45523 21545
rect 45465 21536 45477 21539
rect 45428 21508 45477 21536
rect 45428 21496 45434 21508
rect 45465 21505 45477 21508
rect 45511 21505 45523 21539
rect 47854 21536 47860 21548
rect 47815 21508 47860 21536
rect 45465 21499 45523 21505
rect 47854 21496 47860 21508
rect 47912 21496 47918 21548
rect 47949 21539 48007 21545
rect 47949 21505 47961 21539
rect 47995 21536 48007 21539
rect 48038 21536 48044 21548
rect 47995 21508 48044 21536
rect 47995 21505 48007 21508
rect 47949 21499 48007 21505
rect 48038 21496 48044 21508
rect 48096 21496 48102 21548
rect 32122 21468 32128 21480
rect 32083 21440 32128 21468
rect 32122 21428 32128 21440
rect 32180 21428 32186 21480
rect 32309 21471 32367 21477
rect 32309 21437 32321 21471
rect 32355 21437 32367 21471
rect 32582 21468 32588 21480
rect 32543 21440 32588 21468
rect 32309 21431 32367 21437
rect 30190 21360 30196 21412
rect 30248 21400 30254 21412
rect 31481 21403 31539 21409
rect 31481 21400 31493 21403
rect 30248 21372 31493 21400
rect 30248 21360 30254 21372
rect 31481 21369 31493 21372
rect 31527 21369 31539 21403
rect 32324 21400 32352 21431
rect 32582 21428 32588 21440
rect 32640 21428 32646 21480
rect 44085 21471 44143 21477
rect 44085 21468 44097 21471
rect 41386 21440 44097 21468
rect 41386 21400 41414 21440
rect 44085 21437 44097 21440
rect 44131 21437 44143 21471
rect 44085 21431 44143 21437
rect 44821 21471 44879 21477
rect 44821 21437 44833 21471
rect 44867 21468 44879 21471
rect 45002 21468 45008 21480
rect 44867 21440 45008 21468
rect 44867 21437 44879 21440
rect 44821 21431 44879 21437
rect 45002 21428 45008 21440
rect 45060 21428 45066 21480
rect 46198 21468 46204 21480
rect 46159 21440 46204 21468
rect 46198 21428 46204 21440
rect 46256 21428 46262 21480
rect 48133 21403 48191 21409
rect 48133 21400 48145 21403
rect 32324 21372 41414 21400
rect 41708 21372 48145 21400
rect 31481 21363 31539 21369
rect 34790 21332 34796 21344
rect 30116 21304 34796 21332
rect 34790 21292 34796 21304
rect 34848 21292 34854 21344
rect 40218 21292 40224 21344
rect 40276 21332 40282 21344
rect 41708 21332 41736 21372
rect 48133 21369 48145 21372
rect 48179 21369 48191 21403
rect 48133 21363 48191 21369
rect 40276 21304 41736 21332
rect 40276 21292 40282 21304
rect 42242 21292 42248 21344
rect 42300 21332 42306 21344
rect 46750 21332 46756 21344
rect 42300 21304 46756 21332
rect 42300 21292 42306 21304
rect 46750 21292 46756 21304
rect 46808 21292 46814 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 11882 21128 11888 21140
rect 11471 21100 11888 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 11882 21088 11888 21100
rect 11940 21088 11946 21140
rect 26050 21128 26056 21140
rect 11992 21100 26056 21128
rect 3510 21020 3516 21072
rect 3568 21060 3574 21072
rect 11992 21060 12020 21100
rect 26050 21088 26056 21100
rect 26108 21088 26114 21140
rect 27246 21128 27252 21140
rect 26160 21100 27252 21128
rect 3568 21032 12020 21060
rect 12069 21063 12127 21069
rect 3568 21020 3574 21032
rect 12069 21029 12081 21063
rect 12115 21029 12127 21063
rect 12069 21023 12127 21029
rect 13357 21063 13415 21069
rect 13357 21029 13369 21063
rect 13403 21060 13415 21063
rect 14550 21060 14556 21072
rect 13403 21032 14556 21060
rect 13403 21029 13415 21032
rect 13357 21023 13415 21029
rect 9582 20992 9588 21004
rect 9543 20964 9588 20992
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9861 20995 9919 21001
rect 9861 20961 9873 20995
rect 9907 20992 9919 20995
rect 10134 20992 10140 21004
rect 9907 20964 10140 20992
rect 9907 20961 9919 20964
rect 9861 20955 9919 20961
rect 10134 20952 10140 20964
rect 10192 20952 10198 21004
rect 12084 20992 12112 21023
rect 14550 21020 14556 21032
rect 14608 21020 14614 21072
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 15749 21063 15807 21069
rect 15749 21060 15761 21063
rect 15712 21032 15761 21060
rect 15712 21020 15718 21032
rect 15749 21029 15761 21032
rect 15795 21029 15807 21063
rect 15749 21023 15807 21029
rect 14645 20995 14703 21001
rect 14645 20992 14657 20995
rect 11440 20964 12112 20992
rect 13556 20964 14657 20992
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 11440 20933 11468 20964
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 9180 20896 9505 20924
rect 9180 20884 9186 20896
rect 9493 20893 9505 20896
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20924 11667 20927
rect 12345 20927 12403 20933
rect 11655 20896 12204 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 12069 20859 12127 20865
rect 12069 20856 12081 20859
rect 12032 20828 12081 20856
rect 12032 20816 12038 20828
rect 12069 20825 12081 20828
rect 12115 20825 12127 20859
rect 12176 20856 12204 20896
rect 12345 20893 12357 20927
rect 12391 20924 12403 20927
rect 12526 20924 12532 20936
rect 12391 20896 12532 20924
rect 12391 20893 12403 20896
rect 12345 20887 12403 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 13556 20933 13584 20964
rect 14645 20961 14657 20964
rect 14691 20961 14703 20995
rect 21082 20992 21088 21004
rect 21043 20964 21088 20992
rect 14645 20955 14703 20961
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 21361 20995 21419 21001
rect 21361 20961 21373 20995
rect 21407 20992 21419 20995
rect 23106 20992 23112 21004
rect 21407 20964 23112 20992
rect 21407 20961 21419 20964
rect 21361 20955 21419 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 26160 21001 26188 21100
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 29546 21088 29552 21140
rect 29604 21128 29610 21140
rect 30929 21131 30987 21137
rect 30929 21128 30941 21131
rect 29604 21100 30941 21128
rect 29604 21088 29610 21100
rect 30116 21004 30144 21100
rect 26145 20995 26203 21001
rect 26145 20961 26157 20995
rect 26191 20961 26203 20995
rect 26145 20955 26203 20961
rect 26421 20995 26479 21001
rect 26421 20961 26433 20995
rect 26467 20992 26479 20995
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 26467 20964 27169 20992
rect 26467 20961 26479 20964
rect 26421 20955 26479 20961
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 30009 20995 30067 21001
rect 30009 20961 30021 20995
rect 30055 20992 30067 20995
rect 30098 20992 30104 21004
rect 30055 20964 30104 20992
rect 30055 20961 30067 20964
rect 30009 20955 30067 20961
rect 30098 20952 30104 20964
rect 30156 20952 30162 21004
rect 30190 20952 30196 21004
rect 30248 20992 30254 21004
rect 30377 20995 30435 21001
rect 30377 20992 30389 20995
rect 30248 20964 30389 20992
rect 30248 20952 30254 20964
rect 30377 20961 30389 20964
rect 30423 20961 30435 20995
rect 30852 20992 30880 21100
rect 30929 21097 30941 21100
rect 30975 21097 30987 21131
rect 31202 21128 31208 21140
rect 31163 21100 31208 21128
rect 30929 21091 30987 21097
rect 31202 21088 31208 21100
rect 31260 21088 31266 21140
rect 32030 21128 32036 21140
rect 31991 21100 32036 21128
rect 32030 21088 32036 21100
rect 32088 21088 32094 21140
rect 34790 21128 34796 21140
rect 34751 21100 34796 21128
rect 34790 21088 34796 21100
rect 34848 21128 34854 21140
rect 35437 21131 35495 21137
rect 35437 21128 35449 21131
rect 34848 21100 35449 21128
rect 34848 21088 34854 21100
rect 35437 21097 35449 21100
rect 35483 21097 35495 21131
rect 35437 21091 35495 21097
rect 41693 21063 41751 21069
rect 41693 21029 41705 21063
rect 41739 21060 41751 21063
rect 41739 21032 46336 21060
rect 41739 21029 41751 21032
rect 41693 21023 41751 21029
rect 31573 20995 31631 21001
rect 30852 20964 31248 20992
rect 30377 20955 30435 20961
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20893 14335 20927
rect 14458 20924 14464 20936
rect 14419 20896 14464 20924
rect 14277 20887 14335 20893
rect 12710 20856 12716 20868
rect 12176 20828 12716 20856
rect 12069 20819 12127 20825
rect 12710 20816 12716 20828
rect 12768 20816 12774 20868
rect 14292 20856 14320 20887
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20924 15715 20927
rect 16298 20924 16304 20936
rect 15703 20896 16304 20924
rect 15703 20893 15715 20896
rect 15657 20887 15715 20893
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19426 20924 19432 20936
rect 19291 20896 19432 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 26053 20927 26111 20933
rect 26053 20893 26065 20927
rect 26099 20924 26111 20927
rect 26234 20924 26240 20936
rect 26099 20896 26240 20924
rect 26099 20893 26111 20896
rect 26053 20887 26111 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26878 20924 26884 20936
rect 26839 20896 26884 20924
rect 26878 20884 26884 20896
rect 26936 20884 26942 20936
rect 31113 20927 31171 20933
rect 31113 20924 31125 20927
rect 30760 20896 31125 20924
rect 14366 20856 14372 20868
rect 14292 20828 14372 20856
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 22094 20816 22100 20868
rect 22152 20816 22158 20868
rect 27798 20816 27804 20868
rect 27856 20816 27862 20868
rect 30101 20859 30159 20865
rect 30101 20825 30113 20859
rect 30147 20825 30159 20859
rect 30101 20819 30159 20825
rect 12250 20788 12256 20800
rect 12211 20760 12256 20788
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 19334 20788 19340 20800
rect 19295 20760 19340 20788
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 22738 20748 22744 20800
rect 22796 20788 22802 20800
rect 22833 20791 22891 20797
rect 22833 20788 22845 20791
rect 22796 20760 22845 20788
rect 22796 20748 22802 20760
rect 22833 20757 22845 20760
rect 22879 20757 22891 20791
rect 22833 20751 22891 20757
rect 27522 20748 27528 20800
rect 27580 20788 27586 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 27580 20760 28641 20788
rect 27580 20748 27586 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 30116 20788 30144 20819
rect 30760 20788 30788 20896
rect 31113 20893 31125 20896
rect 31159 20893 31171 20927
rect 31113 20887 31171 20893
rect 31220 20856 31248 20964
rect 31573 20961 31585 20995
rect 31619 20992 31631 20995
rect 35161 20995 35219 21001
rect 31619 20964 31754 20992
rect 31619 20961 31631 20964
rect 31573 20955 31631 20961
rect 31726 20924 31754 20964
rect 35161 20961 35173 20995
rect 35207 20992 35219 20995
rect 36354 20992 36360 21004
rect 35207 20964 36360 20992
rect 35207 20961 35219 20964
rect 35161 20955 35219 20961
rect 36354 20952 36360 20964
rect 36412 20952 36418 21004
rect 46308 21001 46336 21032
rect 42245 20995 42303 21001
rect 42245 20961 42257 20995
rect 42291 20992 42303 20995
rect 42981 20995 43039 21001
rect 42981 20992 42993 20995
rect 42291 20964 42993 20992
rect 42291 20961 42303 20964
rect 42245 20955 42303 20961
rect 42981 20961 42993 20964
rect 43027 20961 43039 20995
rect 42981 20955 43039 20961
rect 46293 20995 46351 21001
rect 46293 20961 46305 20995
rect 46339 20961 46351 20995
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 46293 20955 46351 20961
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 32217 20927 32275 20933
rect 32217 20924 32229 20927
rect 31726 20896 32229 20924
rect 32217 20893 32229 20896
rect 32263 20893 32275 20927
rect 32217 20887 32275 20893
rect 34701 20927 34759 20933
rect 34701 20893 34713 20927
rect 34747 20924 34759 20927
rect 35618 20924 35624 20936
rect 34747 20896 35624 20924
rect 34747 20893 34759 20896
rect 34701 20887 34759 20893
rect 35618 20884 35624 20896
rect 35676 20884 35682 20936
rect 42153 20927 42211 20933
rect 42153 20893 42165 20927
rect 42199 20893 42211 20927
rect 42334 20924 42340 20936
rect 42295 20896 42340 20924
rect 42153 20887 42211 20893
rect 34790 20856 34796 20868
rect 31220 20828 34796 20856
rect 34790 20816 34796 20828
rect 34848 20816 34854 20868
rect 42168 20856 42196 20887
rect 42334 20884 42340 20896
rect 42392 20884 42398 20936
rect 43254 20924 43260 20936
rect 43167 20896 43260 20924
rect 43254 20884 43260 20896
rect 43312 20924 43318 20936
rect 43622 20924 43628 20936
rect 43312 20896 43628 20924
rect 43312 20884 43318 20896
rect 43622 20884 43628 20896
rect 43680 20884 43686 20936
rect 45370 20924 45376 20936
rect 45331 20896 45376 20924
rect 45370 20884 45376 20896
rect 45428 20884 45434 20936
rect 42702 20856 42708 20868
rect 42168 20828 42708 20856
rect 42702 20816 42708 20828
rect 42760 20816 42766 20868
rect 45649 20859 45707 20865
rect 45649 20825 45661 20859
rect 45695 20856 45707 20859
rect 45738 20856 45744 20868
rect 45695 20828 45744 20856
rect 45695 20825 45707 20828
rect 45649 20819 45707 20825
rect 45738 20816 45744 20828
rect 45796 20816 45802 20868
rect 46474 20856 46480 20868
rect 46435 20828 46480 20856
rect 46474 20816 46480 20828
rect 46532 20816 46538 20868
rect 43898 20788 43904 20800
rect 29420 20760 30788 20788
rect 43859 20760 43904 20788
rect 29420 20748 29426 20760
rect 43898 20748 43904 20760
rect 43956 20748 43962 20800
rect 47210 20748 47216 20800
rect 47268 20788 47274 20800
rect 47854 20788 47860 20800
rect 47268 20760 47860 20788
rect 47268 20748 47274 20760
rect 47854 20748 47860 20760
rect 47912 20748 47918 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3418 20544 3424 20596
rect 3476 20584 3482 20596
rect 3476 20556 12664 20584
rect 3476 20544 3482 20556
rect 9306 20516 9312 20528
rect 9267 20488 9312 20516
rect 9306 20476 9312 20488
rect 9364 20476 9370 20528
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 12345 20519 12403 20525
rect 12345 20516 12357 20519
rect 12032 20488 12357 20516
rect 12032 20476 12038 20488
rect 12345 20485 12357 20488
rect 12391 20485 12403 20519
rect 12345 20479 12403 20485
rect 12526 20476 12532 20528
rect 12584 20525 12590 20528
rect 12584 20519 12603 20525
rect 12591 20485 12603 20519
rect 12636 20516 12664 20556
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 14277 20587 14335 20593
rect 12768 20556 12813 20584
rect 12768 20544 12774 20556
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14458 20584 14464 20596
rect 14323 20556 14464 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 14734 20584 14740 20596
rect 14695 20556 14740 20584
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 16632 20556 17325 20584
rect 16632 20544 16638 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22152 20556 22197 20584
rect 22152 20544 22158 20556
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 26292 20556 27169 20584
rect 26292 20544 26298 20556
rect 27157 20553 27169 20556
rect 27203 20584 27215 20587
rect 27522 20584 27528 20596
rect 27203 20556 27528 20584
rect 27203 20553 27215 20556
rect 27157 20547 27215 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 27798 20584 27804 20596
rect 27759 20556 27804 20584
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 36173 20587 36231 20593
rect 36173 20584 36185 20587
rect 34808 20556 36185 20584
rect 18877 20519 18935 20525
rect 12636 20488 18552 20516
rect 12584 20479 12603 20485
rect 12584 20476 12590 20479
rect 9122 20448 9128 20460
rect 9083 20420 9128 20448
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 12434 20448 12440 20460
rect 11563 20420 12440 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 12544 20448 12572 20476
rect 13630 20448 13636 20460
rect 12544 20420 13636 20448
rect 13630 20408 13636 20420
rect 13688 20408 13694 20460
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 15010 20448 15016 20460
rect 13863 20420 15016 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 16114 20408 16120 20460
rect 16172 20448 16178 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16172 20420 16957 20448
rect 16172 20408 16178 20420
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 17037 20451 17095 20457
rect 17037 20426 17049 20451
rect 17083 20426 17095 20451
rect 17129 20451 17187 20457
rect 16945 20411 17003 20417
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20349 9643 20383
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 9585 20343 9643 20349
rect 14384 20352 14473 20380
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 9600 20312 9628 20343
rect 4028 20284 9628 20312
rect 14384 20312 14412 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 14826 20380 14832 20392
rect 14608 20352 14653 20380
rect 14787 20352 14832 20380
rect 14608 20340 14614 20352
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20380 14979 20383
rect 16666 20380 16672 20392
rect 14967 20352 16672 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 16724 20352 16988 20380
rect 17034 20374 17040 20426
rect 17092 20374 17098 20426
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 16724 20340 16730 20352
rect 15194 20312 15200 20324
rect 14384 20284 15200 20312
rect 4028 20272 4034 20284
rect 15194 20272 15200 20284
rect 15252 20312 15258 20324
rect 16022 20312 16028 20324
rect 15252 20284 16028 20312
rect 15252 20272 15258 20284
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 16758 20312 16764 20324
rect 16719 20284 16764 20312
rect 16758 20272 16764 20284
rect 16816 20272 16822 20324
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11480 20216 11621 20244
rect 11480 20204 11486 20216
rect 11609 20213 11621 20216
rect 11655 20213 11667 20247
rect 11609 20207 11667 20213
rect 12250 20204 12256 20256
rect 12308 20244 12314 20256
rect 12529 20247 12587 20253
rect 12529 20244 12541 20247
rect 12308 20216 12541 20244
rect 12308 20204 12314 20216
rect 12529 20213 12541 20216
rect 12575 20213 12587 20247
rect 12529 20207 12587 20213
rect 13725 20247 13783 20253
rect 13725 20213 13737 20247
rect 13771 20244 13783 20247
rect 14366 20244 14372 20256
rect 13771 20216 14372 20244
rect 13771 20213 13783 20216
rect 13725 20207 13783 20213
rect 14366 20204 14372 20216
rect 14424 20204 14430 20256
rect 16960 20244 16988 20352
rect 17144 20244 17172 20411
rect 18524 20312 18552 20488
rect 18877 20485 18889 20519
rect 18923 20516 18935 20519
rect 19334 20516 19340 20528
rect 18923 20488 19340 20516
rect 18923 20485 18935 20488
rect 18877 20479 18935 20485
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 23201 20519 23259 20525
rect 23201 20485 23213 20519
rect 23247 20516 23259 20519
rect 23474 20516 23480 20528
rect 23247 20488 23480 20516
rect 23247 20485 23259 20488
rect 23201 20479 23259 20485
rect 23474 20476 23480 20488
rect 23532 20476 23538 20528
rect 23658 20476 23664 20528
rect 23716 20476 23722 20528
rect 26510 20476 26516 20528
rect 26568 20516 26574 20528
rect 26878 20516 26884 20528
rect 26568 20488 26884 20516
rect 26568 20476 26574 20488
rect 26878 20476 26884 20488
rect 26936 20516 26942 20528
rect 26936 20488 27752 20516
rect 26936 20476 26942 20488
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20448 22063 20451
rect 22830 20448 22836 20460
rect 22051 20420 22836 20448
rect 22051 20417 22063 20420
rect 22005 20411 22063 20417
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25866 20448 25872 20460
rect 25827 20420 25872 20448
rect 25685 20411 25743 20417
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 19242 20380 19248 20392
rect 18739 20352 19248 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 19337 20383 19395 20389
rect 19337 20349 19349 20383
rect 19383 20349 19395 20383
rect 22922 20380 22928 20392
rect 22883 20352 22928 20380
rect 19337 20343 19395 20349
rect 19352 20312 19380 20343
rect 22922 20340 22928 20352
rect 22980 20340 22986 20392
rect 24394 20340 24400 20392
rect 24452 20380 24458 20392
rect 24949 20383 25007 20389
rect 24949 20380 24961 20383
rect 24452 20352 24961 20380
rect 24452 20340 24458 20352
rect 24949 20349 24961 20352
rect 24995 20349 25007 20383
rect 25700 20380 25728 20411
rect 25866 20408 25872 20420
rect 25924 20408 25930 20460
rect 26970 20448 26976 20460
rect 26931 20420 26976 20448
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 27246 20408 27252 20460
rect 27304 20448 27310 20460
rect 27724 20457 27752 20488
rect 28350 20476 28356 20528
rect 28408 20516 28414 20528
rect 34808 20525 34836 20556
rect 36173 20553 36185 20556
rect 36219 20553 36231 20587
rect 36173 20547 36231 20553
rect 44652 20556 45692 20584
rect 34701 20519 34759 20525
rect 34701 20516 34713 20519
rect 28408 20488 34713 20516
rect 28408 20476 28414 20488
rect 34701 20485 34713 20488
rect 34747 20485 34759 20519
rect 34701 20479 34759 20485
rect 34793 20519 34851 20525
rect 34793 20485 34805 20519
rect 34839 20485 34851 20519
rect 44652 20516 44680 20556
rect 34793 20479 34851 20485
rect 43640 20488 44680 20516
rect 27709 20451 27767 20457
rect 27304 20420 27349 20448
rect 27304 20408 27310 20420
rect 27709 20417 27721 20451
rect 27755 20417 27767 20451
rect 27709 20411 27767 20417
rect 30926 20408 30932 20460
rect 30984 20448 30990 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 30984 20420 31493 20448
rect 30984 20408 30990 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 32122 20448 32128 20460
rect 31481 20411 31539 20417
rect 31726 20420 32128 20448
rect 25700 20352 27016 20380
rect 24949 20343 25007 20349
rect 18524 20284 19380 20312
rect 24964 20312 24992 20343
rect 26988 20321 27016 20352
rect 26973 20315 27031 20321
rect 24964 20284 25820 20312
rect 25682 20244 25688 20256
rect 16960 20216 17172 20244
rect 25643 20216 25688 20244
rect 25682 20204 25688 20216
rect 25740 20204 25746 20256
rect 25792 20244 25820 20284
rect 26973 20281 26985 20315
rect 27019 20281 27031 20315
rect 26973 20275 27031 20281
rect 31297 20315 31355 20321
rect 31297 20281 31309 20315
rect 31343 20312 31355 20315
rect 31726 20312 31754 20420
rect 32122 20408 32128 20420
rect 32180 20448 32186 20460
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 32180 20420 32321 20448
rect 32180 20408 32186 20420
rect 32309 20417 32321 20420
rect 32355 20417 32367 20451
rect 36354 20448 36360 20460
rect 36315 20420 36360 20448
rect 32309 20411 32367 20417
rect 36354 20408 36360 20420
rect 36412 20408 36418 20460
rect 41690 20408 41696 20460
rect 41748 20448 41754 20460
rect 42705 20451 42763 20457
rect 42705 20448 42717 20451
rect 41748 20420 42717 20448
rect 41748 20408 41754 20420
rect 42705 20417 42717 20420
rect 42751 20417 42763 20451
rect 42705 20411 42763 20417
rect 42794 20408 42800 20460
rect 42852 20448 42858 20460
rect 42889 20451 42947 20457
rect 42889 20448 42901 20451
rect 42852 20420 42901 20448
rect 42852 20408 42858 20420
rect 42889 20417 42901 20420
rect 42935 20448 42947 20451
rect 43070 20448 43076 20460
rect 42935 20420 43076 20448
rect 42935 20417 42947 20420
rect 42889 20411 42947 20417
rect 43070 20408 43076 20420
rect 43128 20408 43134 20460
rect 32493 20383 32551 20389
rect 32493 20349 32505 20383
rect 32539 20380 32551 20383
rect 33134 20380 33140 20392
rect 32539 20352 33140 20380
rect 32539 20349 32551 20352
rect 32493 20343 32551 20349
rect 33134 20340 33140 20352
rect 33192 20340 33198 20392
rect 34146 20380 34152 20392
rect 34107 20352 34152 20380
rect 34146 20340 34152 20352
rect 34204 20340 34210 20392
rect 35710 20380 35716 20392
rect 35671 20352 35716 20380
rect 35710 20340 35716 20352
rect 35768 20340 35774 20392
rect 43162 20340 43168 20392
rect 43220 20380 43226 20392
rect 43640 20389 43668 20488
rect 44652 20457 44680 20488
rect 45373 20519 45431 20525
rect 45373 20485 45385 20519
rect 45419 20516 45431 20519
rect 45554 20516 45560 20528
rect 45419 20488 45560 20516
rect 45419 20485 45431 20488
rect 45373 20479 45431 20485
rect 45554 20476 45560 20488
rect 45612 20476 45618 20528
rect 45664 20516 45692 20556
rect 47026 20544 47032 20596
rect 47084 20584 47090 20596
rect 47949 20587 48007 20593
rect 47949 20584 47961 20587
rect 47084 20556 47961 20584
rect 47084 20544 47090 20556
rect 47949 20553 47961 20556
rect 47995 20553 48007 20587
rect 47949 20547 48007 20553
rect 47581 20519 47639 20525
rect 45664 20488 47164 20516
rect 43809 20451 43867 20457
rect 43809 20448 43821 20451
rect 43732 20420 43821 20448
rect 43625 20383 43683 20389
rect 43625 20380 43637 20383
rect 43220 20352 43637 20380
rect 43220 20340 43226 20352
rect 43625 20349 43637 20352
rect 43671 20349 43683 20383
rect 43625 20343 43683 20349
rect 42702 20312 42708 20324
rect 31343 20284 31754 20312
rect 42663 20284 42708 20312
rect 31343 20281 31355 20284
rect 31297 20275 31355 20281
rect 42702 20272 42708 20284
rect 42760 20272 42766 20324
rect 42978 20272 42984 20324
rect 43036 20312 43042 20324
rect 43732 20312 43760 20420
rect 43809 20417 43821 20420
rect 43855 20448 43867 20451
rect 44453 20451 44511 20457
rect 44453 20448 44465 20451
rect 43855 20420 44465 20448
rect 43855 20417 43867 20420
rect 43809 20411 43867 20417
rect 44453 20417 44465 20420
rect 44499 20417 44511 20451
rect 44453 20411 44511 20417
rect 44637 20451 44695 20457
rect 44637 20417 44649 20451
rect 44683 20417 44695 20451
rect 44637 20411 44695 20417
rect 43898 20340 43904 20392
rect 43956 20380 43962 20392
rect 45189 20383 45247 20389
rect 45189 20380 45201 20383
rect 43956 20352 45201 20380
rect 43956 20340 43962 20352
rect 45189 20349 45201 20352
rect 45235 20349 45247 20383
rect 47026 20380 47032 20392
rect 46987 20352 47032 20380
rect 45189 20343 45247 20349
rect 47026 20340 47032 20352
rect 47084 20340 47090 20392
rect 47136 20380 47164 20488
rect 47581 20485 47593 20519
rect 47627 20516 47639 20519
rect 47670 20516 47676 20528
rect 47627 20488 47676 20516
rect 47627 20485 47639 20488
rect 47581 20479 47639 20485
rect 47670 20476 47676 20488
rect 47728 20476 47734 20528
rect 47486 20408 47492 20460
rect 47544 20448 47550 20460
rect 47765 20451 47823 20457
rect 47765 20448 47777 20451
rect 47544 20420 47777 20448
rect 47544 20408 47550 20420
rect 47765 20417 47777 20420
rect 47811 20417 47823 20451
rect 47765 20411 47823 20417
rect 47946 20380 47952 20392
rect 47136 20352 47952 20380
rect 47946 20340 47952 20352
rect 48004 20340 48010 20392
rect 43036 20284 43760 20312
rect 43036 20272 43042 20284
rect 43806 20272 43812 20324
rect 43864 20312 43870 20324
rect 44453 20315 44511 20321
rect 44453 20312 44465 20315
rect 43864 20284 44465 20312
rect 43864 20272 43870 20284
rect 44453 20281 44465 20284
rect 44499 20281 44511 20315
rect 44453 20275 44511 20281
rect 37274 20244 37280 20256
rect 25792 20216 37280 20244
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 43993 20247 44051 20253
rect 43993 20213 44005 20247
rect 44039 20244 44051 20247
rect 44174 20244 44180 20256
rect 44039 20216 44180 20244
rect 44039 20213 44051 20216
rect 43993 20207 44051 20213
rect 44174 20204 44180 20216
rect 44232 20204 44238 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 9180 20012 11621 20040
rect 9180 20000 9186 20012
rect 11609 20009 11621 20012
rect 11655 20040 11667 20043
rect 12250 20040 12256 20052
rect 11655 20012 12256 20040
rect 11655 20009 11667 20012
rect 11609 20003 11667 20009
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 15010 20040 15016 20052
rect 14971 20012 15016 20040
rect 15010 20000 15016 20012
rect 15068 20040 15074 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 15068 20012 16313 20040
rect 15068 20000 15074 20012
rect 16301 20009 16313 20012
rect 16347 20040 16359 20043
rect 17034 20040 17040 20052
rect 16347 20012 17040 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 22922 20040 22928 20052
rect 22883 20012 22928 20040
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 23569 20043 23627 20049
rect 23569 20009 23581 20043
rect 23615 20040 23627 20043
rect 23658 20040 23664 20052
rect 23615 20012 23664 20040
rect 23615 20009 23627 20012
rect 23569 20003 23627 20009
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 43622 20040 43628 20052
rect 25516 20012 31754 20040
rect 43583 20012 43628 20040
rect 14461 19975 14519 19981
rect 14461 19941 14473 19975
rect 14507 19972 14519 19975
rect 15194 19972 15200 19984
rect 14507 19944 15200 19972
rect 14507 19941 14519 19944
rect 14461 19935 14519 19941
rect 15194 19932 15200 19944
rect 15252 19932 15258 19984
rect 16485 19975 16543 19981
rect 16485 19941 16497 19975
rect 16531 19941 16543 19975
rect 16485 19935 16543 19941
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 16500 19904 16528 19935
rect 18690 19932 18696 19984
rect 18748 19972 18754 19984
rect 25516 19972 25544 20012
rect 30190 19972 30196 19984
rect 18748 19944 25544 19972
rect 29748 19944 30196 19972
rect 18748 19932 18754 19944
rect 17218 19904 17224 19916
rect 16500 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19904 17555 19907
rect 18046 19904 18052 19916
rect 17543 19876 18052 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 20990 19904 20996 19916
rect 18564 19876 20996 19904
rect 18564 19864 18570 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 9858 19836 9864 19848
rect 9819 19808 9864 19836
rect 2041 19799 2099 19805
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11532 19808 12173 19836
rect 11422 19768 11428 19780
rect 11362 19740 11428 19768
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 11532 19700 11560 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12176 19768 12204 19799
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 14826 19836 14832 19848
rect 12308 19808 14832 19836
rect 12308 19796 12314 19808
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 16758 19796 16764 19848
rect 16816 19836 16822 19848
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 16816 19808 17141 19836
rect 16816 19796 16822 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 18322 19836 18328 19848
rect 18187 19808 18328 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 13814 19768 13820 19780
rect 12176 19740 13820 19768
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 14734 19768 14740 19780
rect 14695 19740 14740 19768
rect 14734 19728 14740 19740
rect 14792 19728 14798 19780
rect 16114 19768 16120 19780
rect 16075 19740 16120 19768
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 16333 19771 16391 19777
rect 16333 19737 16345 19771
rect 16379 19768 16391 19771
rect 16666 19768 16672 19780
rect 16379 19740 16672 19768
rect 16379 19737 16391 19740
rect 16333 19731 16391 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 17144 19768 17172 19799
rect 18322 19796 18328 19808
rect 18380 19836 18386 19848
rect 20070 19836 20076 19848
rect 18380 19808 20076 19836
rect 18380 19796 18386 19808
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 20732 19845 20760 19876
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 25682 19904 25688 19916
rect 22756 19876 24808 19904
rect 25643 19876 25688 19904
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 22756 19845 22784 19876
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 20956 19808 22753 19836
rect 20956 19796 20962 19808
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 24780 19845 24808 19876
rect 25682 19864 25688 19876
rect 25740 19864 25746 19916
rect 23477 19839 23535 19845
rect 23477 19836 23489 19839
rect 22888 19808 23489 19836
rect 22888 19796 22894 19808
rect 23477 19805 23489 19808
rect 23523 19805 23535 19839
rect 23477 19799 23535 19805
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 24854 19836 24860 19848
rect 24811 19808 24860 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 24995 19808 25421 19836
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 29748 19845 29776 19944
rect 30190 19932 30196 19944
rect 30248 19932 30254 19984
rect 30926 19972 30932 19984
rect 30887 19944 30932 19972
rect 30926 19932 30932 19944
rect 30984 19932 30990 19984
rect 31726 19972 31754 20012
rect 43622 20000 43628 20012
rect 43680 20000 43686 20052
rect 45373 20043 45431 20049
rect 45373 20009 45385 20043
rect 45419 20040 45431 20043
rect 46474 20040 46480 20052
rect 45419 20012 46480 20040
rect 45419 20009 45431 20012
rect 45373 20003 45431 20009
rect 46474 20000 46480 20012
rect 46532 20000 46538 20052
rect 34146 19972 34152 19984
rect 31726 19944 34152 19972
rect 34146 19932 34152 19944
rect 34204 19932 34210 19984
rect 34790 19932 34796 19984
rect 34848 19972 34854 19984
rect 46658 19972 46664 19984
rect 34848 19944 46664 19972
rect 34848 19932 34854 19944
rect 35176 19913 35204 19944
rect 46658 19932 46664 19944
rect 46716 19932 46722 19984
rect 30101 19907 30159 19913
rect 30101 19873 30113 19907
rect 30147 19904 30159 19907
rect 35161 19907 35219 19913
rect 30147 19876 30788 19904
rect 30147 19873 30159 19876
rect 30101 19867 30159 19873
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29696 19808 29745 19836
rect 29696 19796 29702 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 30006 19796 30012 19848
rect 30064 19836 30070 19848
rect 30760 19845 30788 19876
rect 35161 19873 35173 19907
rect 35207 19873 35219 19907
rect 35161 19867 35219 19873
rect 35710 19864 35716 19916
rect 35768 19904 35774 19916
rect 36173 19907 36231 19913
rect 36173 19904 36185 19907
rect 35768 19876 36185 19904
rect 35768 19864 35774 19876
rect 36173 19873 36185 19876
rect 36219 19904 36231 19907
rect 47026 19904 47032 19916
rect 36219 19876 41414 19904
rect 46987 19876 47032 19904
rect 36219 19873 36231 19876
rect 36173 19867 36231 19873
rect 30561 19839 30619 19845
rect 30561 19836 30573 19839
rect 30064 19808 30573 19836
rect 30064 19796 30070 19808
rect 30561 19805 30573 19808
rect 30607 19805 30619 19839
rect 30561 19799 30619 19805
rect 30745 19839 30803 19845
rect 30745 19805 30757 19839
rect 30791 19805 30803 19839
rect 30745 19799 30803 19805
rect 33594 19796 33600 19848
rect 33652 19836 33658 19848
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 33652 19808 33793 19836
rect 33652 19796 33658 19808
rect 33781 19805 33793 19808
rect 33827 19805 33839 19839
rect 41386 19836 41414 19876
rect 47026 19864 47032 19876
rect 47084 19864 47090 19916
rect 42978 19836 42984 19848
rect 41386 19808 42984 19836
rect 33781 19799 33839 19805
rect 42978 19796 42984 19808
rect 43036 19796 43042 19848
rect 43162 19836 43168 19848
rect 43123 19808 43168 19836
rect 43162 19796 43168 19808
rect 43220 19796 43226 19848
rect 43806 19836 43812 19848
rect 43767 19808 43812 19836
rect 43806 19796 43812 19808
rect 43864 19796 43870 19848
rect 44085 19839 44143 19845
rect 44085 19805 44097 19839
rect 44131 19836 44143 19839
rect 44542 19836 44548 19848
rect 44131 19808 44548 19836
rect 44131 19805 44143 19808
rect 44085 19799 44143 19805
rect 44542 19796 44548 19808
rect 44600 19796 44606 19848
rect 45002 19796 45008 19848
rect 45060 19836 45066 19848
rect 45281 19839 45339 19845
rect 45281 19836 45293 19839
rect 45060 19808 45293 19836
rect 45060 19796 45066 19808
rect 45281 19805 45293 19808
rect 45327 19805 45339 19839
rect 45281 19799 45339 19805
rect 45646 19796 45652 19848
rect 45704 19836 45710 19848
rect 45925 19839 45983 19845
rect 45925 19836 45937 19839
rect 45704 19808 45937 19836
rect 45704 19796 45710 19808
rect 45925 19805 45937 19808
rect 45971 19805 45983 19839
rect 45925 19799 45983 19805
rect 19242 19768 19248 19780
rect 17144 19740 19248 19768
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 27062 19768 27068 19780
rect 26910 19740 27068 19768
rect 27062 19728 27068 19740
rect 27120 19728 27126 19780
rect 29822 19728 29828 19780
rect 29880 19768 29886 19780
rect 29917 19771 29975 19777
rect 29917 19768 29929 19771
rect 29880 19740 29929 19768
rect 29880 19728 29886 19740
rect 29917 19737 29929 19740
rect 29963 19737 29975 19771
rect 29917 19731 29975 19737
rect 35253 19771 35311 19777
rect 35253 19737 35265 19771
rect 35299 19768 35311 19771
rect 35618 19768 35624 19780
rect 35299 19740 35624 19768
rect 35299 19737 35311 19740
rect 35253 19731 35311 19737
rect 35618 19728 35624 19740
rect 35676 19728 35682 19780
rect 43073 19771 43131 19777
rect 43073 19737 43085 19771
rect 43119 19768 43131 19771
rect 43993 19771 44051 19777
rect 43993 19768 44005 19771
rect 43119 19740 44005 19768
rect 43119 19737 43131 19740
rect 43073 19731 43131 19737
rect 43993 19737 44005 19740
rect 44039 19737 44051 19771
rect 46106 19768 46112 19780
rect 46067 19740 46112 19768
rect 43993 19731 44051 19737
rect 46106 19728 46112 19740
rect 46164 19728 46170 19780
rect 10468 19672 11560 19700
rect 10468 19660 10474 19672
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 11756 19672 12357 19700
rect 11756 19660 11762 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 13446 19660 13452 19712
rect 13504 19700 13510 19712
rect 14550 19700 14556 19712
rect 13504 19672 14556 19700
rect 13504 19660 13510 19672
rect 14550 19660 14556 19672
rect 14608 19700 14614 19712
rect 14645 19703 14703 19709
rect 14645 19700 14657 19703
rect 14608 19672 14657 19700
rect 14608 19660 14614 19672
rect 14645 19669 14657 19672
rect 14691 19669 14703 19703
rect 14645 19663 14703 19669
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17828 19672 18153 19700
rect 17828 19660 17834 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 20806 19700 20812 19712
rect 20767 19672 20812 19700
rect 18141 19663 18199 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 26510 19660 26516 19712
rect 26568 19700 26574 19712
rect 26970 19700 26976 19712
rect 26568 19672 26976 19700
rect 26568 19660 26574 19672
rect 26970 19660 26976 19672
rect 27028 19700 27034 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27028 19672 27169 19700
rect 27028 19660 27034 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 33870 19700 33876 19712
rect 33831 19672 33876 19700
rect 27157 19663 27215 19669
rect 33870 19660 33876 19672
rect 33928 19660 33934 19712
rect 33962 19660 33968 19712
rect 34020 19700 34026 19712
rect 38286 19700 38292 19712
rect 34020 19672 38292 19700
rect 34020 19660 34026 19672
rect 38286 19660 38292 19672
rect 38344 19660 38350 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 9916 19468 10517 19496
rect 9916 19456 9922 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 27062 19496 27068 19508
rect 10505 19459 10563 19465
rect 10612 19468 23428 19496
rect 27023 19468 27068 19496
rect 4890 19388 4896 19440
rect 4948 19428 4954 19440
rect 10612 19428 10640 19468
rect 4948 19400 10640 19428
rect 4948 19388 4954 19400
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 12492 19400 13032 19428
rect 12492 19388 12498 19400
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 10410 19360 10416 19372
rect 10371 19332 10416 19360
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 13004 19369 13032 19400
rect 15746 19388 15752 19440
rect 15804 19428 15810 19440
rect 16114 19428 16120 19440
rect 15804 19400 15976 19428
rect 16075 19400 16120 19428
rect 15804 19388 15810 19400
rect 15948 19369 15976 19400
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 19334 19428 19340 19440
rect 19274 19400 19340 19428
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 23106 19388 23112 19440
rect 23164 19388 23170 19440
rect 23400 19428 23428 19468
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 29917 19499 29975 19505
rect 29917 19465 29929 19499
rect 29963 19496 29975 19499
rect 30006 19496 30012 19508
rect 29963 19468 30012 19496
rect 29963 19465 29975 19468
rect 29917 19459 29975 19465
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 33229 19499 33287 19505
rect 33229 19465 33241 19499
rect 33275 19465 33287 19499
rect 33229 19459 33287 19465
rect 33704 19468 38240 19496
rect 28994 19428 29000 19440
rect 23400 19400 29000 19428
rect 28994 19388 29000 19400
rect 29052 19428 29058 19440
rect 29822 19428 29828 19440
rect 29052 19400 29828 19428
rect 29052 19388 29058 19400
rect 29822 19388 29828 19400
rect 29880 19428 29886 19440
rect 33244 19428 33272 19459
rect 29880 19400 29960 19428
rect 29880 19388 29886 19400
rect 12161 19363 12219 19369
rect 12161 19329 12173 19363
rect 12207 19360 12219 19363
rect 12989 19363 13047 19369
rect 12207 19332 12940 19360
rect 12207 19329 12219 19332
rect 12161 19323 12219 19329
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12710 19292 12716 19304
rect 12299 19264 12716 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 12912 19292 12940 19332
rect 12989 19329 13001 19363
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 14507 19332 15945 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 16724 19332 16896 19360
rect 16724 19320 16730 19332
rect 13446 19292 13452 19304
rect 12912 19264 13452 19292
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 14366 19292 14372 19304
rect 14327 19264 14372 19292
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19292 15807 19295
rect 16758 19292 16764 19304
rect 15795 19264 16764 19292
rect 15795 19261 15807 19264
rect 15749 19255 15807 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 16868 19301 16896 19332
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17770 19360 17776 19372
rect 17000 19332 17045 19360
rect 17731 19332 17776 19360
rect 17000 19320 17006 19332
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20128 19332 20729 19360
rect 20128 19320 20134 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 24394 19360 24400 19372
rect 24351 19332 24400 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 24489 19363 24547 19369
rect 24489 19329 24501 19363
rect 24535 19360 24547 19363
rect 24762 19360 24768 19372
rect 24535 19332 24768 19360
rect 24535 19329 24547 19332
rect 24489 19323 24547 19329
rect 24762 19320 24768 19332
rect 24820 19320 24826 19372
rect 26878 19320 26884 19372
rect 26936 19360 26942 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26936 19332 26985 19360
rect 26936 19320 26942 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 29932 19369 29960 19400
rect 32324 19400 33272 19428
rect 32324 19369 32352 19400
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29696 19332 29745 19360
rect 29696 19320 29702 19332
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29917 19363 29975 19369
rect 29917 19329 29929 19363
rect 29963 19329 29975 19363
rect 29917 19323 29975 19329
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 32769 19363 32827 19369
rect 32769 19329 32781 19363
rect 32815 19360 32827 19363
rect 33134 19360 33140 19372
rect 32815 19332 33140 19360
rect 32815 19329 32827 19332
rect 32769 19323 32827 19329
rect 33134 19320 33140 19332
rect 33192 19360 33198 19372
rect 33704 19369 33732 19468
rect 33870 19428 33876 19440
rect 33831 19400 33876 19428
rect 33870 19388 33876 19400
rect 33928 19388 33934 19440
rect 38212 19428 38240 19468
rect 38286 19456 38292 19508
rect 38344 19496 38350 19508
rect 45922 19496 45928 19508
rect 38344 19468 45928 19496
rect 38344 19456 38350 19468
rect 45922 19456 45928 19468
rect 45980 19456 45986 19508
rect 47118 19496 47124 19508
rect 46032 19468 47124 19496
rect 43898 19428 43904 19440
rect 38212 19400 43904 19428
rect 43898 19388 43904 19400
rect 43956 19388 43962 19440
rect 33689 19363 33747 19369
rect 33192 19332 33640 19360
rect 33192 19320 33198 19332
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 16853 19255 16911 19261
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 18046 19292 18052 19304
rect 17184 19264 17229 19292
rect 18007 19264 18052 19292
rect 17184 19252 17190 19264
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19300 19264 19533 19292
rect 19300 19252 19306 19264
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 21818 19292 21824 19304
rect 21779 19264 21824 19292
rect 19521 19255 19579 19261
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 33612 19292 33640 19332
rect 33689 19329 33701 19363
rect 33735 19329 33747 19363
rect 35526 19360 35532 19372
rect 35487 19332 35532 19360
rect 33689 19323 33747 19329
rect 35526 19320 35532 19332
rect 35584 19320 35590 19372
rect 37274 19360 37280 19372
rect 37235 19332 37280 19360
rect 37274 19320 37280 19332
rect 37332 19320 37338 19372
rect 39114 19360 39120 19372
rect 39075 19332 39120 19360
rect 39114 19320 39120 19332
rect 39172 19320 39178 19372
rect 44542 19360 44548 19372
rect 44503 19332 44548 19360
rect 44542 19320 44548 19332
rect 44600 19320 44606 19372
rect 33962 19292 33968 19304
rect 22152 19264 22197 19292
rect 33612 19264 33968 19292
rect 22152 19252 22158 19264
rect 33962 19252 33968 19264
rect 34020 19252 34026 19304
rect 37458 19292 37464 19304
rect 37419 19264 37464 19292
rect 37458 19252 37464 19264
rect 37516 19252 37522 19304
rect 44082 19252 44088 19304
rect 44140 19292 44146 19304
rect 44269 19295 44327 19301
rect 44269 19292 44281 19295
rect 44140 19264 44281 19292
rect 44140 19252 44146 19264
rect 44269 19261 44281 19264
rect 44315 19261 44327 19295
rect 45094 19292 45100 19304
rect 45055 19264 45100 19292
rect 44269 19255 44327 19261
rect 45094 19252 45100 19264
rect 45152 19252 45158 19304
rect 46032 19301 46060 19468
rect 47118 19456 47124 19468
rect 47176 19496 47182 19508
rect 47949 19499 48007 19505
rect 47949 19496 47961 19499
rect 47176 19468 47961 19496
rect 47176 19456 47182 19468
rect 47949 19465 47961 19468
rect 47995 19465 48007 19499
rect 47949 19459 48007 19465
rect 46106 19388 46112 19440
rect 46164 19428 46170 19440
rect 46293 19431 46351 19437
rect 46293 19428 46305 19431
rect 46164 19400 46305 19428
rect 46164 19388 46170 19400
rect 46293 19397 46305 19400
rect 46339 19397 46351 19431
rect 47857 19431 47915 19437
rect 47857 19428 47869 19431
rect 46293 19391 46351 19397
rect 46400 19400 47869 19428
rect 46400 19372 46428 19400
rect 47857 19397 47869 19400
rect 47903 19397 47915 19431
rect 47857 19391 47915 19397
rect 46382 19360 46388 19372
rect 46343 19332 46388 19360
rect 46382 19320 46388 19332
rect 46440 19320 46446 19372
rect 46753 19363 46811 19369
rect 46753 19360 46765 19363
rect 46492 19332 46765 19360
rect 46017 19295 46075 19301
rect 46017 19261 46029 19295
rect 46063 19261 46075 19295
rect 46017 19255 46075 19261
rect 3970 19184 3976 19236
rect 4028 19224 4034 19236
rect 4028 19196 17908 19224
rect 4028 19184 4034 19196
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12529 19159 12587 19165
rect 12529 19156 12541 19159
rect 12032 19128 12541 19156
rect 12032 19116 12038 19128
rect 12529 19125 12541 19128
rect 12575 19125 12587 19159
rect 13078 19156 13084 19168
rect 13039 19128 13084 19156
rect 12529 19119 12587 19125
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 14734 19156 14740 19168
rect 14695 19128 14740 19156
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 16669 19159 16727 19165
rect 16669 19125 16681 19159
rect 16715 19156 16727 19159
rect 17310 19156 17316 19168
rect 16715 19128 17316 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17880 19156 17908 19196
rect 19076 19196 21404 19224
rect 19076 19156 19104 19196
rect 20898 19156 20904 19168
rect 17880 19128 19104 19156
rect 20859 19128 20904 19156
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 21376 19156 21404 19196
rect 23382 19184 23388 19236
rect 23440 19224 23446 19236
rect 23569 19227 23627 19233
rect 23569 19224 23581 19227
rect 23440 19196 23581 19224
rect 23440 19184 23446 19196
rect 23569 19193 23581 19196
rect 23615 19193 23627 19227
rect 31018 19224 31024 19236
rect 23569 19187 23627 19193
rect 24136 19196 31024 19224
rect 24136 19156 24164 19196
rect 31018 19184 31024 19196
rect 31076 19184 31082 19236
rect 33134 19184 33140 19236
rect 33192 19224 33198 19236
rect 33192 19196 45876 19224
rect 33192 19184 33198 19196
rect 24302 19156 24308 19168
rect 21376 19128 24164 19156
rect 24263 19128 24308 19156
rect 24302 19116 24308 19128
rect 24360 19116 24366 19168
rect 32125 19159 32183 19165
rect 32125 19125 32137 19159
rect 32171 19156 32183 19159
rect 32306 19156 32312 19168
rect 32171 19128 32312 19156
rect 32171 19125 32183 19128
rect 32125 19119 32183 19125
rect 32306 19116 32312 19128
rect 32364 19116 32370 19168
rect 33042 19156 33048 19168
rect 33003 19128 33048 19156
rect 33042 19116 33048 19128
rect 33100 19116 33106 19168
rect 43622 19156 43628 19168
rect 43583 19128 43628 19156
rect 43622 19116 43628 19128
rect 43680 19116 43686 19168
rect 45848 19156 45876 19196
rect 45922 19184 45928 19236
rect 45980 19224 45986 19236
rect 46492 19224 46520 19332
rect 46753 19329 46765 19332
rect 46799 19360 46811 19363
rect 47029 19363 47087 19369
rect 46799 19332 46980 19360
rect 46799 19329 46811 19332
rect 46753 19323 46811 19329
rect 46952 19292 46980 19332
rect 47029 19329 47041 19363
rect 47075 19360 47087 19363
rect 47075 19332 47624 19360
rect 47075 19329 47087 19332
rect 47029 19323 47087 19329
rect 46952 19264 47440 19292
rect 45980 19196 46520 19224
rect 45980 19184 45986 19196
rect 47412 19168 47440 19264
rect 47596 19233 47624 19332
rect 47670 19320 47676 19372
rect 47728 19360 47734 19372
rect 47765 19363 47823 19369
rect 47765 19360 47777 19363
rect 47728 19332 47777 19360
rect 47728 19320 47734 19332
rect 47765 19329 47777 19332
rect 47811 19329 47823 19363
rect 47765 19323 47823 19329
rect 48038 19252 48044 19304
rect 48096 19292 48102 19304
rect 48133 19295 48191 19301
rect 48133 19292 48145 19295
rect 48096 19264 48145 19292
rect 48096 19252 48102 19264
rect 48133 19261 48145 19264
rect 48179 19261 48191 19295
rect 48133 19255 48191 19261
rect 47581 19227 47639 19233
rect 47581 19193 47593 19227
rect 47627 19224 47639 19227
rect 47762 19224 47768 19236
rect 47627 19196 47768 19224
rect 47627 19193 47639 19196
rect 47581 19187 47639 19193
rect 47762 19184 47768 19196
rect 47820 19184 47826 19236
rect 46382 19156 46388 19168
rect 45848 19128 46388 19156
rect 46382 19116 46388 19128
rect 46440 19116 46446 19168
rect 47394 19116 47400 19168
rect 47452 19156 47458 19168
rect 47670 19156 47676 19168
rect 47452 19128 47676 19156
rect 47452 19116 47458 19128
rect 47670 19116 47676 19128
rect 47728 19116 47734 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 6638 18952 6644 18964
rect 2225 18915 2283 18921
rect 2746 18924 6644 18952
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 2746 18884 2774 18924
rect 6638 18912 6644 18924
rect 6696 18952 6702 18964
rect 46014 18952 46020 18964
rect 6696 18924 46020 18952
rect 6696 18912 6702 18924
rect 46014 18912 46020 18924
rect 46072 18912 46078 18964
rect 2188 18856 2774 18884
rect 2188 18844 2194 18856
rect 15746 18844 15752 18896
rect 15804 18884 15810 18896
rect 16209 18887 16267 18893
rect 16209 18884 16221 18887
rect 15804 18856 16221 18884
rect 15804 18844 15810 18856
rect 16209 18853 16221 18856
rect 16255 18884 16267 18887
rect 17034 18884 17040 18896
rect 16255 18856 17040 18884
rect 16255 18853 16267 18856
rect 16209 18847 16267 18853
rect 17034 18844 17040 18856
rect 17092 18844 17098 18896
rect 17310 18884 17316 18896
rect 17271 18856 17316 18884
rect 17310 18844 17316 18856
rect 17368 18844 17374 18896
rect 17678 18844 17684 18896
rect 17736 18884 17742 18896
rect 17862 18884 17868 18896
rect 17736 18856 17868 18884
rect 17736 18844 17742 18856
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 19334 18884 19340 18896
rect 19295 18856 19340 18884
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 23017 18887 23075 18893
rect 20640 18856 22094 18884
rect 11698 18816 11704 18828
rect 11659 18788 11704 18816
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11974 18816 11980 18828
rect 11935 18788 11980 18816
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 14734 18816 14740 18828
rect 14695 18788 14740 18816
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17126 18816 17132 18828
rect 16816 18788 17132 18816
rect 16816 18776 16822 18788
rect 17126 18776 17132 18788
rect 17184 18816 17190 18828
rect 20070 18816 20076 18828
rect 17184 18788 20076 18816
rect 17184 18776 17190 18788
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 20640 18825 20668 18856
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18785 20683 18819
rect 20806 18816 20812 18828
rect 20767 18788 20812 18816
rect 20625 18779 20683 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 22066 18816 22094 18856
rect 23017 18853 23029 18887
rect 23063 18884 23075 18887
rect 23106 18884 23112 18896
rect 23063 18856 23112 18884
rect 23063 18853 23075 18856
rect 23017 18847 23075 18853
rect 23106 18844 23112 18856
rect 23164 18844 23170 18896
rect 24394 18844 24400 18896
rect 24452 18884 24458 18896
rect 24489 18887 24547 18893
rect 24489 18884 24501 18887
rect 24452 18856 24501 18884
rect 24452 18844 24458 18856
rect 24489 18853 24501 18856
rect 24535 18853 24547 18887
rect 24489 18847 24547 18853
rect 37185 18887 37243 18893
rect 37185 18853 37197 18887
rect 37231 18884 37243 18887
rect 37458 18884 37464 18896
rect 37231 18856 37464 18884
rect 37231 18853 37243 18856
rect 37185 18847 37243 18853
rect 37458 18844 37464 18856
rect 37516 18844 37522 18896
rect 47762 18884 47768 18896
rect 41386 18856 47768 18884
rect 25038 18816 25044 18828
rect 22066 18788 23612 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 13078 18708 13084 18760
rect 13136 18708 13142 18760
rect 14090 18708 14096 18760
rect 14148 18748 14154 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14148 18720 14473 18748
rect 14148 18708 14154 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 15838 18708 15844 18760
rect 15896 18708 15902 18760
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17218 18748 17224 18760
rect 17083 18720 17224 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18748 19303 18751
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 19291 18720 19901 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 19889 18717 19901 18720
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 19260 18680 19288 18711
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22888 18720 22937 18748
rect 22888 18708 22894 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 17420 18652 19288 18680
rect 13446 18612 13452 18624
rect 13407 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 17420 18612 17448 18652
rect 22370 18640 22376 18692
rect 22428 18680 22434 18692
rect 22465 18683 22523 18689
rect 22465 18680 22477 18683
rect 22428 18652 22477 18680
rect 22428 18640 22434 18652
rect 22465 18649 22477 18652
rect 22511 18649 22523 18683
rect 23584 18680 23612 18788
rect 23676 18788 25044 18816
rect 23676 18757 23704 18788
rect 25038 18776 25044 18788
rect 25096 18816 25102 18828
rect 26510 18816 26516 18828
rect 25096 18788 25912 18816
rect 26471 18788 26516 18816
rect 25096 18776 25102 18788
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 24765 18751 24823 18757
rect 23661 18711 23719 18717
rect 24320 18720 24716 18748
rect 24320 18680 24348 18720
rect 23584 18652 24348 18680
rect 22465 18643 22523 18649
rect 24394 18640 24400 18692
rect 24452 18680 24458 18692
rect 24489 18683 24547 18689
rect 24489 18680 24501 18683
rect 24452 18652 24501 18680
rect 24452 18640 24458 18652
rect 24489 18649 24501 18652
rect 24535 18649 24547 18683
rect 24688 18680 24716 18720
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 25774 18748 25780 18760
rect 24811 18720 25780 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 25884 18757 25912 18788
rect 26510 18776 26516 18788
rect 26568 18776 26574 18828
rect 28905 18819 28963 18825
rect 28905 18785 28917 18819
rect 28951 18816 28963 18819
rect 29825 18819 29883 18825
rect 29825 18816 29837 18819
rect 28951 18788 29837 18816
rect 28951 18785 28963 18788
rect 28905 18779 28963 18785
rect 29825 18785 29837 18788
rect 29871 18785 29883 18819
rect 29825 18779 29883 18785
rect 30285 18819 30343 18825
rect 30285 18785 30297 18819
rect 30331 18785 30343 18819
rect 31018 18816 31024 18828
rect 30979 18788 31024 18816
rect 30285 18779 30343 18785
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 28810 18748 28816 18760
rect 28771 18720 28816 18748
rect 25869 18711 25927 18717
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 28994 18748 29000 18760
rect 28955 18720 29000 18748
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18748 29975 18751
rect 30006 18748 30012 18760
rect 29963 18720 30012 18748
rect 29963 18717 29975 18720
rect 29917 18711 29975 18717
rect 30006 18708 30012 18720
rect 30064 18708 30070 18760
rect 30300 18748 30328 18779
rect 31018 18776 31024 18788
rect 31076 18776 31082 18828
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 41386 18816 41414 18856
rect 47762 18844 47768 18856
rect 47820 18844 47826 18896
rect 33100 18788 41414 18816
rect 33100 18776 33106 18788
rect 30558 18748 30564 18760
rect 30300 18720 30564 18748
rect 30558 18708 30564 18720
rect 30616 18708 30622 18760
rect 32769 18751 32827 18757
rect 32769 18717 32781 18751
rect 32815 18748 32827 18751
rect 33134 18748 33140 18760
rect 32815 18720 33140 18748
rect 32815 18717 32827 18720
rect 32769 18711 32827 18717
rect 25961 18683 26019 18689
rect 24688 18652 25912 18680
rect 24489 18643 24547 18649
rect 16356 18584 17448 18612
rect 17497 18615 17555 18621
rect 16356 18572 16362 18584
rect 17497 18581 17509 18615
rect 17543 18612 17555 18615
rect 17586 18612 17592 18624
rect 17543 18584 17592 18612
rect 17543 18581 17555 18584
rect 17497 18575 17555 18581
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 18046 18572 18052 18624
rect 18104 18612 18110 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 18104 18584 18337 18612
rect 18104 18572 18110 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 18325 18575 18383 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 23290 18572 23296 18624
rect 23348 18612 23354 18624
rect 23753 18615 23811 18621
rect 23753 18612 23765 18615
rect 23348 18584 23765 18612
rect 23348 18572 23354 18584
rect 23753 18581 23765 18584
rect 23799 18581 23811 18615
rect 23753 18575 23811 18581
rect 24578 18572 24584 18624
rect 24636 18612 24642 18624
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 24636 18584 24685 18612
rect 24636 18572 24642 18584
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 25884 18612 25912 18652
rect 25961 18649 25973 18683
rect 26007 18680 26019 18683
rect 26697 18683 26755 18689
rect 26697 18680 26709 18683
rect 26007 18652 26709 18680
rect 26007 18649 26019 18652
rect 25961 18643 26019 18649
rect 26697 18649 26709 18652
rect 26743 18649 26755 18683
rect 28350 18680 28356 18692
rect 28311 18652 28356 18680
rect 26697 18643 26755 18649
rect 28350 18640 28356 18652
rect 28408 18640 28414 18692
rect 30745 18683 30803 18689
rect 30745 18649 30757 18683
rect 30791 18680 30803 18683
rect 31018 18680 31024 18692
rect 30791 18652 31024 18680
rect 30791 18649 30803 18652
rect 30745 18643 30803 18649
rect 31018 18640 31024 18652
rect 31076 18640 31082 18692
rect 26234 18612 26240 18624
rect 25884 18584 26240 18612
rect 24673 18575 24731 18581
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 26878 18572 26884 18624
rect 26936 18612 26942 18624
rect 32784 18612 32812 18711
rect 33134 18708 33140 18720
rect 33192 18708 33198 18760
rect 33336 18757 33364 18788
rect 43622 18776 43628 18828
rect 43680 18816 43686 18828
rect 46293 18819 46351 18825
rect 46293 18816 46305 18819
rect 43680 18788 46305 18816
rect 43680 18776 43686 18788
rect 46293 18785 46305 18788
rect 46339 18785 46351 18819
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 46293 18779 46351 18785
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 33321 18751 33379 18757
rect 33321 18717 33333 18751
rect 33367 18717 33379 18751
rect 33321 18711 33379 18717
rect 33597 18751 33655 18757
rect 33597 18717 33609 18751
rect 33643 18748 33655 18751
rect 33962 18748 33968 18760
rect 33643 18720 33968 18748
rect 33643 18717 33655 18720
rect 33597 18711 33655 18717
rect 33962 18708 33968 18720
rect 34020 18708 34026 18760
rect 37090 18748 37096 18760
rect 37051 18720 37096 18748
rect 37090 18708 37096 18720
rect 37148 18708 37154 18760
rect 43806 18708 43812 18760
rect 43864 18748 43870 18760
rect 43993 18751 44051 18757
rect 43993 18748 44005 18751
rect 43864 18720 44005 18748
rect 43864 18708 43870 18720
rect 43993 18717 44005 18720
rect 44039 18717 44051 18751
rect 44174 18748 44180 18760
rect 44135 18720 44180 18748
rect 43993 18711 44051 18717
rect 44174 18708 44180 18720
rect 44232 18708 44238 18760
rect 45186 18748 45192 18760
rect 45147 18720 45192 18748
rect 45186 18708 45192 18720
rect 45244 18708 45250 18760
rect 45370 18748 45376 18760
rect 45331 18720 45376 18748
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 33781 18683 33839 18689
rect 33781 18649 33793 18683
rect 33827 18680 33839 18683
rect 34606 18680 34612 18692
rect 33827 18652 34612 18680
rect 33827 18649 33839 18652
rect 33781 18643 33839 18649
rect 34606 18640 34612 18652
rect 34664 18640 34670 18692
rect 44082 18680 44088 18692
rect 44043 18652 44088 18680
rect 44082 18640 44088 18652
rect 44140 18640 44146 18692
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 26936 18584 32812 18612
rect 26936 18572 26942 18584
rect 37090 18572 37096 18624
rect 37148 18612 37154 18624
rect 45002 18612 45008 18624
rect 37148 18584 45008 18612
rect 37148 18572 37154 18584
rect 45002 18572 45008 18584
rect 45060 18572 45066 18624
rect 45278 18612 45284 18624
rect 45239 18584 45284 18612
rect 45278 18572 45284 18584
rect 45336 18572 45342 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1578 18368 1584 18420
rect 1636 18408 1642 18420
rect 14090 18408 14096 18420
rect 1636 18380 2774 18408
rect 14051 18380 14096 18408
rect 1636 18368 1642 18380
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 2746 18204 2774 18380
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 15838 18408 15844 18420
rect 15799 18380 15844 18408
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 18414 18408 18420 18420
rect 15948 18380 18420 18408
rect 3326 18300 3332 18352
rect 3384 18340 3390 18352
rect 15948 18340 15976 18380
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 18708 18380 20116 18408
rect 18708 18340 18736 18380
rect 19978 18340 19984 18352
rect 3384 18312 15976 18340
rect 16546 18312 18736 18340
rect 19550 18312 19984 18340
rect 3384 18300 3390 18312
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13872 18244 14013 18272
rect 13872 18232 13878 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 16298 18272 16304 18284
rect 15795 18244 16304 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 16546 18204 16574 18312
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 20088 18340 20116 18380
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 22005 18411 22063 18417
rect 22005 18408 22017 18411
rect 21876 18380 22017 18408
rect 21876 18368 21882 18380
rect 22005 18377 22017 18380
rect 22051 18377 22063 18411
rect 26878 18408 26884 18420
rect 22005 18371 22063 18377
rect 23124 18380 26884 18408
rect 23124 18340 23152 18380
rect 26878 18368 26884 18380
rect 26936 18368 26942 18420
rect 28810 18368 28816 18420
rect 28868 18408 28874 18420
rect 30009 18411 30067 18417
rect 30009 18408 30021 18411
rect 28868 18380 30021 18408
rect 28868 18368 28874 18380
rect 30009 18377 30021 18380
rect 30055 18377 30067 18411
rect 31018 18408 31024 18420
rect 30979 18380 31024 18408
rect 30009 18371 30067 18377
rect 31018 18368 31024 18380
rect 31076 18368 31082 18420
rect 43993 18411 44051 18417
rect 43993 18377 44005 18411
rect 44039 18408 44051 18411
rect 44450 18408 44456 18420
rect 44039 18380 44456 18408
rect 44039 18377 44051 18380
rect 43993 18371 44051 18377
rect 44450 18368 44456 18380
rect 44508 18408 44514 18420
rect 47670 18408 47676 18420
rect 44508 18380 46428 18408
rect 47631 18380 47676 18408
rect 44508 18368 44514 18380
rect 23290 18340 23296 18352
rect 20088 18312 23152 18340
rect 23251 18312 23296 18340
rect 23290 18300 23296 18312
rect 23348 18300 23354 18352
rect 28534 18300 28540 18352
rect 28592 18340 28598 18352
rect 29641 18343 29699 18349
rect 29641 18340 29653 18343
rect 28592 18312 29653 18340
rect 28592 18300 28598 18312
rect 29641 18309 29653 18312
rect 29687 18309 29699 18343
rect 29641 18303 29699 18309
rect 30558 18300 30564 18352
rect 30616 18340 30622 18352
rect 32306 18340 32312 18352
rect 30616 18312 31754 18340
rect 32267 18312 32312 18340
rect 30616 18300 30622 18312
rect 17586 18272 17592 18284
rect 17547 18244 17592 18272
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 18046 18272 18052 18284
rect 18007 18244 18052 18272
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 20956 18244 21833 18272
rect 20956 18232 20962 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 25409 18275 25467 18281
rect 25409 18272 25421 18275
rect 24912 18244 25421 18272
rect 24912 18232 24918 18244
rect 25409 18241 25421 18244
rect 25455 18272 25467 18275
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 25455 18244 26157 18272
rect 25455 18241 25467 18244
rect 25409 18235 25467 18241
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 28074 18272 28080 18284
rect 28035 18244 28080 18272
rect 26145 18235 26203 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 28721 18275 28779 18281
rect 28721 18241 28733 18275
rect 28767 18272 28779 18275
rect 28810 18272 28816 18284
rect 28767 18244 28816 18272
rect 28767 18241 28779 18244
rect 28721 18235 28779 18241
rect 28810 18232 28816 18244
rect 28868 18272 28874 18284
rect 29825 18275 29883 18281
rect 29825 18272 29837 18275
rect 28868 18244 29837 18272
rect 28868 18232 28874 18244
rect 29825 18241 29837 18244
rect 29871 18241 29883 18275
rect 30926 18272 30932 18284
rect 30887 18244 30932 18272
rect 29825 18235 29883 18241
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 31726 18272 31754 18312
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 34606 18340 34612 18352
rect 34567 18312 34612 18340
rect 34606 18300 34612 18312
rect 34664 18300 34670 18352
rect 45922 18340 45928 18352
rect 44192 18312 45928 18340
rect 32125 18275 32183 18281
rect 32125 18272 32137 18275
rect 31726 18244 32137 18272
rect 32125 18241 32137 18244
rect 32171 18241 32183 18275
rect 32125 18235 32183 18241
rect 33594 18232 33600 18284
rect 33652 18272 33658 18284
rect 44192 18281 44220 18312
rect 45922 18300 45928 18312
rect 45980 18300 45986 18352
rect 46400 18349 46428 18380
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 46385 18343 46443 18349
rect 46385 18309 46397 18343
rect 46431 18309 46443 18343
rect 46385 18303 46443 18309
rect 34425 18275 34483 18281
rect 34425 18272 34437 18275
rect 33652 18244 34437 18272
rect 33652 18232 33658 18244
rect 34425 18241 34437 18244
rect 34471 18241 34483 18275
rect 34425 18235 34483 18241
rect 44177 18275 44235 18281
rect 44177 18241 44189 18275
rect 44223 18241 44235 18275
rect 44726 18272 44732 18284
rect 44687 18244 44732 18272
rect 44177 18235 44235 18241
rect 44726 18232 44732 18244
rect 44784 18232 44790 18284
rect 45278 18232 45284 18284
rect 45336 18232 45342 18284
rect 46201 18275 46259 18281
rect 46201 18241 46213 18275
rect 46247 18241 46259 18275
rect 46201 18235 46259 18241
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 2746 18176 16574 18204
rect 17420 18176 18337 18204
rect 17420 18145 17448 18176
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 23109 18207 23167 18213
rect 18472 18176 22094 18204
rect 18472 18164 18478 18176
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 17405 18139 17463 18145
rect 1627 18108 2774 18136
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 2746 18068 2774 18108
rect 17405 18105 17417 18139
rect 17451 18105 17463 18139
rect 22066 18136 22094 18176
rect 23109 18173 23121 18207
rect 23155 18204 23167 18207
rect 23382 18204 23388 18216
rect 23155 18176 23388 18204
rect 23155 18173 23167 18176
rect 23109 18167 23167 18173
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 23569 18207 23627 18213
rect 23569 18173 23581 18207
rect 23615 18173 23627 18207
rect 23569 18167 23627 18173
rect 23584 18136 23612 18167
rect 28902 18164 28908 18216
rect 28960 18204 28966 18216
rect 28997 18207 29055 18213
rect 28997 18204 29009 18207
rect 28960 18176 29009 18204
rect 28960 18164 28966 18176
rect 28997 18173 29009 18176
rect 29043 18173 29055 18207
rect 28997 18167 29055 18173
rect 29089 18207 29147 18213
rect 29089 18173 29101 18207
rect 29135 18204 29147 18207
rect 29546 18204 29552 18216
rect 29135 18176 29552 18204
rect 29135 18173 29147 18176
rect 29089 18167 29147 18173
rect 29546 18164 29552 18176
rect 29604 18164 29610 18216
rect 30944 18204 30972 18232
rect 33686 18204 33692 18216
rect 30944 18176 33692 18204
rect 33686 18164 33692 18176
rect 33744 18164 33750 18216
rect 33965 18207 34023 18213
rect 33965 18173 33977 18207
rect 34011 18204 34023 18207
rect 34146 18204 34152 18216
rect 34011 18176 34152 18204
rect 34011 18173 34023 18176
rect 33965 18167 34023 18173
rect 34146 18164 34152 18176
rect 34204 18204 34210 18216
rect 36265 18207 36323 18213
rect 36265 18204 36277 18207
rect 34204 18176 36277 18204
rect 34204 18164 34210 18176
rect 36265 18173 36277 18176
rect 36311 18204 36323 18207
rect 41874 18204 41880 18216
rect 36311 18176 41880 18204
rect 36311 18173 36323 18176
rect 36265 18167 36323 18173
rect 41874 18164 41880 18176
rect 41932 18164 41938 18216
rect 45646 18204 45652 18216
rect 45607 18176 45652 18204
rect 45646 18164 45652 18176
rect 45704 18164 45710 18216
rect 45922 18164 45928 18216
rect 45980 18204 45986 18216
rect 46216 18204 46244 18235
rect 47486 18232 47492 18284
rect 47544 18272 47550 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47544 18244 47593 18272
rect 47544 18232 47550 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 45980 18176 46244 18204
rect 45980 18164 45986 18176
rect 27982 18136 27988 18148
rect 17405 18099 17463 18105
rect 19720 18108 20024 18136
rect 22066 18108 23612 18136
rect 25056 18108 27988 18136
rect 19720 18068 19748 18108
rect 2746 18040 19748 18068
rect 19797 18071 19855 18077
rect 19797 18037 19809 18071
rect 19843 18068 19855 18071
rect 19886 18068 19892 18080
rect 19843 18040 19892 18068
rect 19843 18037 19855 18040
rect 19797 18031 19855 18037
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 19996 18068 20024 18108
rect 25056 18068 25084 18108
rect 27982 18096 27988 18108
rect 28040 18096 28046 18148
rect 28169 18139 28227 18145
rect 28169 18105 28181 18139
rect 28215 18136 28227 18139
rect 29638 18136 29644 18148
rect 28215 18108 29644 18136
rect 28215 18105 28227 18108
rect 28169 18099 28227 18105
rect 29638 18096 29644 18108
rect 29696 18096 29702 18148
rect 30190 18096 30196 18148
rect 30248 18136 30254 18148
rect 37090 18136 37096 18148
rect 30248 18108 37096 18136
rect 30248 18096 30254 18108
rect 37090 18096 37096 18108
rect 37148 18096 37154 18148
rect 45186 18096 45192 18148
rect 45244 18136 45250 18148
rect 46569 18139 46627 18145
rect 46569 18136 46581 18139
rect 45244 18108 46581 18136
rect 45244 18096 45250 18108
rect 46569 18105 46581 18108
rect 46615 18105 46627 18139
rect 46569 18099 46627 18105
rect 25406 18068 25412 18080
rect 19996 18040 25084 18068
rect 25367 18040 25412 18068
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 26237 18071 26295 18077
rect 26237 18037 26249 18071
rect 26283 18068 26295 18071
rect 26326 18068 26332 18080
rect 26283 18040 26332 18068
rect 26283 18037 26295 18040
rect 26237 18031 26295 18037
rect 26326 18028 26332 18040
rect 26384 18028 26390 18080
rect 28534 18028 28540 18080
rect 28592 18068 28598 18080
rect 28813 18071 28871 18077
rect 28813 18068 28825 18071
rect 28592 18040 28825 18068
rect 28592 18028 28598 18040
rect 28813 18037 28825 18040
rect 28859 18037 28871 18071
rect 29086 18068 29092 18080
rect 29047 18040 29092 18068
rect 28813 18031 28871 18037
rect 29086 18028 29092 18040
rect 29144 18028 29150 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 22152 17836 22937 17864
rect 22152 17824 22158 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24949 17867 25007 17873
rect 24949 17864 24961 17867
rect 24084 17836 24961 17864
rect 24084 17824 24090 17836
rect 24949 17833 24961 17836
rect 24995 17833 25007 17867
rect 24949 17827 25007 17833
rect 44542 17824 44548 17876
rect 44600 17864 44606 17876
rect 45649 17867 45707 17873
rect 45649 17864 45661 17867
rect 44600 17836 45661 17864
rect 44600 17824 44606 17836
rect 45649 17833 45661 17836
rect 45695 17833 45707 17867
rect 45649 17827 45707 17833
rect 23750 17796 23756 17808
rect 23124 17768 23756 17796
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17728 20039 17731
rect 20254 17728 20260 17740
rect 20027 17700 20260 17728
rect 20027 17697 20039 17700
rect 19981 17691 20039 17697
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 23124 17669 23152 17768
rect 23750 17756 23756 17768
rect 23808 17756 23814 17808
rect 27706 17796 27712 17808
rect 25608 17768 27712 17796
rect 23382 17728 23388 17740
rect 23343 17700 23388 17728
rect 23382 17688 23388 17700
rect 23440 17728 23446 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 23440 17700 24409 17728
rect 23440 17688 23446 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17660 23351 17663
rect 24762 17660 24768 17672
rect 23339 17632 24768 17660
rect 23339 17629 23351 17632
rect 23293 17623 23351 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25608 17669 25636 17768
rect 27706 17756 27712 17768
rect 27764 17756 27770 17808
rect 28445 17799 28503 17805
rect 28445 17765 28457 17799
rect 28491 17796 28503 17799
rect 44726 17796 44732 17808
rect 28491 17768 44732 17796
rect 28491 17765 28503 17768
rect 28445 17759 28503 17765
rect 44726 17756 44732 17768
rect 44784 17796 44790 17808
rect 44784 17768 45508 17796
rect 44784 17756 44790 17768
rect 25685 17731 25743 17737
rect 25685 17697 25697 17731
rect 25731 17728 25743 17731
rect 25774 17728 25780 17740
rect 25731 17700 25780 17728
rect 25731 17697 25743 17700
rect 25685 17691 25743 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 25961 17731 26019 17737
rect 25961 17697 25973 17731
rect 26007 17728 26019 17731
rect 26234 17728 26240 17740
rect 26007 17700 26240 17728
rect 26007 17697 26019 17700
rect 25961 17691 26019 17697
rect 26234 17688 26240 17700
rect 26292 17688 26298 17740
rect 27890 17728 27896 17740
rect 26344 17700 27896 17728
rect 25593 17663 25651 17669
rect 25593 17629 25605 17663
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 11054 17592 11060 17604
rect 3568 17564 11060 17592
rect 3568 17552 3574 17564
rect 11054 17552 11060 17564
rect 11112 17552 11118 17604
rect 20162 17592 20168 17604
rect 20123 17564 20168 17592
rect 20162 17552 20168 17564
rect 20220 17552 20226 17604
rect 21821 17595 21879 17601
rect 21821 17561 21833 17595
rect 21867 17592 21879 17595
rect 21910 17592 21916 17604
rect 21867 17564 21916 17592
rect 21867 17561 21879 17564
rect 21821 17555 21879 17561
rect 21910 17552 21916 17564
rect 21968 17552 21974 17604
rect 24670 17592 24676 17604
rect 24583 17564 24676 17592
rect 24670 17552 24676 17564
rect 24728 17592 24734 17604
rect 25608 17592 25636 17623
rect 24728 17564 25636 17592
rect 24728 17552 24734 17564
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 24394 17524 24400 17536
rect 22244 17496 24400 17524
rect 22244 17484 22250 17496
rect 24394 17484 24400 17496
rect 24452 17524 24458 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 24452 17496 24593 17524
rect 24452 17484 24458 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24765 17527 24823 17533
rect 24765 17493 24777 17527
rect 24811 17524 24823 17527
rect 26344 17524 26372 17700
rect 27890 17688 27896 17700
rect 27948 17688 27954 17740
rect 44361 17731 44419 17737
rect 44361 17697 44373 17731
rect 44407 17728 44419 17731
rect 45370 17728 45376 17740
rect 44407 17700 45376 17728
rect 44407 17697 44419 17700
rect 44361 17691 44419 17697
rect 45370 17688 45376 17700
rect 45428 17688 45434 17740
rect 45480 17737 45508 17768
rect 45465 17731 45523 17737
rect 45465 17697 45477 17731
rect 45511 17697 45523 17731
rect 45465 17691 45523 17697
rect 26421 17663 26479 17669
rect 26421 17629 26433 17663
rect 26467 17660 26479 17663
rect 26970 17660 26976 17672
rect 26467 17632 26976 17660
rect 26467 17629 26479 17632
rect 26421 17623 26479 17629
rect 26970 17620 26976 17632
rect 27028 17660 27034 17672
rect 27065 17663 27123 17669
rect 27065 17660 27077 17663
rect 27028 17632 27077 17660
rect 27028 17620 27034 17632
rect 27065 17629 27077 17632
rect 27111 17629 27123 17663
rect 27798 17660 27804 17672
rect 27759 17632 27804 17660
rect 27065 17623 27123 17629
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 27982 17660 27988 17672
rect 27943 17632 27988 17660
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 29086 17660 29092 17672
rect 28675 17632 29092 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 29086 17620 29092 17632
rect 29144 17620 29150 17672
rect 29546 17620 29552 17672
rect 29604 17660 29610 17672
rect 29641 17663 29699 17669
rect 29641 17660 29653 17663
rect 29604 17632 29653 17660
rect 29604 17620 29610 17632
rect 29641 17629 29653 17632
rect 29687 17629 29699 17663
rect 29822 17660 29828 17672
rect 29783 17632 29828 17660
rect 29641 17623 29699 17629
rect 29822 17620 29828 17632
rect 29880 17620 29886 17672
rect 44269 17663 44327 17669
rect 44269 17629 44281 17663
rect 44315 17629 44327 17663
rect 44450 17660 44456 17672
rect 44411 17632 44456 17660
rect 44269 17623 44327 17629
rect 27893 17595 27951 17601
rect 27893 17561 27905 17595
rect 27939 17592 27951 17595
rect 28074 17592 28080 17604
rect 27939 17564 28080 17592
rect 27939 17561 27951 17564
rect 27893 17555 27951 17561
rect 28074 17552 28080 17564
rect 28132 17592 28138 17604
rect 28997 17595 29055 17601
rect 28132 17564 28856 17592
rect 28132 17552 28138 17564
rect 26510 17524 26516 17536
rect 24811 17496 26372 17524
rect 26471 17496 26516 17524
rect 24811 17493 24823 17496
rect 24765 17487 24823 17493
rect 26510 17484 26516 17496
rect 26568 17484 26574 17536
rect 27157 17527 27215 17533
rect 27157 17493 27169 17527
rect 27203 17524 27215 17527
rect 27246 17524 27252 17536
rect 27203 17496 27252 17524
rect 27203 17493 27215 17496
rect 27157 17487 27215 17493
rect 27246 17484 27252 17496
rect 27304 17484 27310 17536
rect 28626 17484 28632 17536
rect 28684 17524 28690 17536
rect 28828 17533 28856 17564
rect 28997 17561 29009 17595
rect 29043 17592 29055 17595
rect 29178 17592 29184 17604
rect 29043 17564 29184 17592
rect 29043 17561 29055 17564
rect 28997 17555 29055 17561
rect 29178 17552 29184 17564
rect 29236 17552 29242 17604
rect 44284 17592 44312 17623
rect 44450 17620 44456 17632
rect 44508 17620 44514 17672
rect 45005 17663 45063 17669
rect 45005 17629 45017 17663
rect 45051 17660 45063 17663
rect 45186 17660 45192 17672
rect 45051 17632 45192 17660
rect 45051 17629 45063 17632
rect 45005 17623 45063 17629
rect 45186 17620 45192 17632
rect 45244 17620 45250 17672
rect 46290 17660 46296 17672
rect 46251 17632 46296 17660
rect 46290 17620 46296 17632
rect 46348 17620 46354 17672
rect 45922 17592 45928 17604
rect 44284 17564 45928 17592
rect 45922 17552 45928 17564
rect 45980 17552 45986 17604
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 28721 17527 28779 17533
rect 28721 17524 28733 17527
rect 28684 17496 28733 17524
rect 28684 17484 28690 17496
rect 28721 17493 28733 17496
rect 28767 17493 28779 17527
rect 28721 17487 28779 17493
rect 28813 17527 28871 17533
rect 28813 17493 28825 17527
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 30653 17527 30711 17533
rect 30653 17493 30665 17527
rect 30699 17524 30711 17527
rect 33594 17524 33600 17536
rect 30699 17496 33600 17524
rect 30699 17493 30711 17496
rect 30653 17487 30711 17493
rect 33594 17484 33600 17496
rect 33652 17484 33658 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 27798 17320 27804 17332
rect 20272 17292 27804 17320
rect 5442 17212 5448 17264
rect 5500 17252 5506 17264
rect 20272 17252 20300 17292
rect 27798 17280 27804 17292
rect 27856 17320 27862 17332
rect 27856 17292 27936 17320
rect 27856 17280 27862 17292
rect 5500 17224 20300 17252
rect 21177 17255 21235 17261
rect 5500 17212 5506 17224
rect 21177 17221 21189 17255
rect 21223 17252 21235 17255
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21223 17224 22017 17252
rect 21223 17221 21235 17224
rect 21177 17215 21235 17221
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 24302 17212 24308 17264
rect 24360 17252 24366 17264
rect 24397 17255 24455 17261
rect 24397 17252 24409 17255
rect 24360 17224 24409 17252
rect 24360 17212 24366 17224
rect 24397 17221 24409 17224
rect 24443 17221 24455 17255
rect 26510 17252 26516 17264
rect 25622 17224 26516 17252
rect 24397 17215 24455 17221
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20990 17184 20996 17196
rect 20119 17156 20996 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20990 17144 20996 17156
rect 21048 17184 21054 17196
rect 27908 17193 27936 17292
rect 28626 17280 28632 17332
rect 28684 17320 28690 17332
rect 28813 17323 28871 17329
rect 28813 17320 28825 17323
rect 28684 17292 28825 17320
rect 28684 17280 28690 17292
rect 28813 17289 28825 17292
rect 28859 17320 28871 17323
rect 28994 17320 29000 17332
rect 28859 17292 29000 17320
rect 28859 17289 28871 17292
rect 28813 17283 28871 17289
rect 28994 17280 29000 17292
rect 29052 17280 29058 17332
rect 29641 17323 29699 17329
rect 29641 17289 29653 17323
rect 29687 17320 29699 17323
rect 29822 17320 29828 17332
rect 29687 17292 29828 17320
rect 29687 17289 29699 17292
rect 29641 17283 29699 17289
rect 29822 17280 29828 17292
rect 29880 17280 29886 17332
rect 30098 17320 30104 17332
rect 30024 17292 30104 17320
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 21048 17156 21097 17184
rect 21048 17144 21054 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 27893 17187 27951 17193
rect 27893 17153 27905 17187
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 27982 17144 27988 17196
rect 28040 17184 28046 17196
rect 28077 17187 28135 17193
rect 28077 17184 28089 17187
rect 28040 17156 28089 17184
rect 28040 17144 28046 17156
rect 28077 17153 28089 17156
rect 28123 17153 28135 17187
rect 28077 17147 28135 17153
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28629 17187 28687 17193
rect 28629 17184 28641 17187
rect 28592 17156 28641 17184
rect 28592 17144 28598 17156
rect 28629 17153 28641 17156
rect 28675 17153 28687 17187
rect 28810 17184 28816 17196
rect 28771 17156 28816 17184
rect 28629 17147 28687 17153
rect 28810 17144 28816 17156
rect 28868 17144 28874 17196
rect 29086 17144 29092 17196
rect 29144 17184 29150 17196
rect 29457 17187 29515 17193
rect 29457 17184 29469 17187
rect 29144 17156 29469 17184
rect 29144 17144 29150 17156
rect 29457 17153 29469 17156
rect 29503 17153 29515 17187
rect 29457 17147 29515 17153
rect 30024 17128 30052 17292
rect 30098 17280 30104 17292
rect 30156 17280 30162 17332
rect 47670 17320 47676 17332
rect 47631 17292 47676 17320
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 35802 17212 35808 17264
rect 35860 17252 35866 17264
rect 35860 17224 47624 17252
rect 35860 17212 35866 17224
rect 33594 17184 33600 17196
rect 33555 17156 33600 17184
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 47596 17193 47624 17224
rect 47581 17187 47639 17193
rect 47581 17153 47593 17187
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 21821 17119 21879 17125
rect 21821 17085 21833 17119
rect 21867 17116 21879 17119
rect 22186 17116 22192 17128
rect 21867 17088 22192 17116
rect 21867 17085 21879 17088
rect 21821 17079 21879 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 22281 17119 22339 17125
rect 22281 17085 22293 17119
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17116 24179 17119
rect 25406 17116 25412 17128
rect 24167 17088 25412 17116
rect 24167 17085 24179 17088
rect 24121 17079 24179 17085
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 22296 17048 22324 17079
rect 25406 17076 25412 17088
rect 25464 17076 25470 17128
rect 28994 17076 29000 17128
rect 29052 17116 29058 17128
rect 29273 17119 29331 17125
rect 29273 17116 29285 17119
rect 29052 17088 29285 17116
rect 29052 17076 29058 17088
rect 29273 17085 29285 17088
rect 29319 17085 29331 17119
rect 29273 17079 29331 17085
rect 30006 17076 30012 17128
rect 30064 17076 30070 17128
rect 33778 17116 33784 17128
rect 33739 17088 33784 17116
rect 33778 17076 33784 17088
rect 33836 17076 33842 17128
rect 35434 17116 35440 17128
rect 35395 17088 35440 17116
rect 35434 17076 35440 17088
rect 35492 17076 35498 17128
rect 45189 17119 45247 17125
rect 45189 17085 45201 17119
rect 45235 17085 45247 17119
rect 45189 17079 45247 17085
rect 45373 17119 45431 17125
rect 45373 17085 45385 17119
rect 45419 17116 45431 17119
rect 46658 17116 46664 17128
rect 45419 17088 46664 17116
rect 45419 17085 45431 17088
rect 45373 17079 45431 17085
rect 13872 17020 22324 17048
rect 27893 17051 27951 17057
rect 13872 17008 13878 17020
rect 27893 17017 27905 17051
rect 27939 17048 27951 17051
rect 29178 17048 29184 17060
rect 27939 17020 29184 17048
rect 27939 17017 27951 17020
rect 27893 17011 27951 17017
rect 29178 17008 29184 17020
rect 29236 17008 29242 17060
rect 45204 17048 45232 17079
rect 46658 17076 46664 17088
rect 46716 17076 46722 17128
rect 46842 17116 46848 17128
rect 46803 17088 46848 17116
rect 46842 17076 46848 17088
rect 46900 17076 46906 17128
rect 46750 17048 46756 17060
rect 45204 17020 46756 17048
rect 46750 17008 46756 17020
rect 46808 17008 46814 17060
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 25869 16983 25927 16989
rect 25869 16980 25881 16983
rect 24452 16952 25881 16980
rect 24452 16940 24458 16952
rect 25869 16949 25881 16952
rect 25915 16949 25927 16983
rect 25869 16943 25927 16949
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 24578 16776 24584 16788
rect 24539 16748 24584 16776
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 26326 16776 26332 16788
rect 25976 16748 26332 16776
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 20036 16612 20177 16640
rect 20036 16600 20042 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20990 16600 20996 16652
rect 21048 16640 21054 16652
rect 25976 16649 26004 16748
rect 26326 16736 26332 16748
rect 26384 16736 26390 16788
rect 29546 16776 29552 16788
rect 29507 16748 29552 16776
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 33778 16776 33784 16788
rect 33739 16748 33784 16776
rect 33778 16736 33784 16748
rect 33836 16736 33842 16788
rect 46290 16736 46296 16788
rect 46348 16776 46354 16788
rect 48133 16779 48191 16785
rect 48133 16776 48145 16779
rect 46348 16748 48145 16776
rect 46348 16736 46354 16748
rect 48133 16745 48145 16748
rect 48179 16745 48191 16779
rect 48133 16739 48191 16745
rect 45646 16708 45652 16720
rect 45020 16680 45652 16708
rect 25961 16643 26019 16649
rect 21048 16612 22508 16640
rect 21048 16600 21054 16612
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 22480 16581 22508 16612
rect 25961 16609 25973 16643
rect 26007 16609 26019 16643
rect 26234 16640 26240 16652
rect 26195 16612 26240 16640
rect 25961 16603 26019 16609
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 29178 16600 29184 16652
rect 29236 16640 29242 16652
rect 29236 16612 29592 16640
rect 29236 16600 29242 16612
rect 29564 16581 29592 16612
rect 29638 16600 29644 16652
rect 29696 16640 29702 16652
rect 45020 16649 45048 16680
rect 45646 16668 45652 16680
rect 45704 16668 45710 16720
rect 45005 16643 45063 16649
rect 29696 16612 29776 16640
rect 29696 16600 29702 16612
rect 29748 16581 29776 16612
rect 45005 16609 45017 16643
rect 45051 16609 45063 16643
rect 45462 16640 45468 16652
rect 45423 16612 45468 16640
rect 45005 16603 45063 16609
rect 45462 16600 45468 16612
rect 45520 16600 45526 16652
rect 46934 16600 46940 16652
rect 46992 16640 46998 16652
rect 46992 16612 47348 16640
rect 46992 16600 46998 16612
rect 47320 16584 47348 16612
rect 19521 16575 19579 16581
rect 19521 16572 19533 16575
rect 19484 16544 19533 16572
rect 19484 16532 19490 16544
rect 19521 16541 19533 16544
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 29549 16575 29607 16581
rect 29549 16541 29561 16575
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 33686 16572 33692 16584
rect 33647 16544 33692 16572
rect 29733 16535 29791 16541
rect 33686 16532 33692 16544
rect 33744 16532 33750 16584
rect 47302 16572 47308 16584
rect 47215 16544 47308 16572
rect 47302 16532 47308 16544
rect 47360 16532 47366 16584
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 20349 16507 20407 16513
rect 20349 16504 20361 16507
rect 19659 16476 20361 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 20349 16473 20361 16476
rect 20395 16473 20407 16507
rect 22002 16504 22008 16516
rect 21963 16476 22008 16504
rect 20349 16467 20407 16473
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 24394 16504 24400 16516
rect 24355 16476 24400 16504
rect 24394 16464 24400 16476
rect 24452 16464 24458 16516
rect 24613 16507 24671 16513
rect 24613 16473 24625 16507
rect 24659 16504 24671 16507
rect 25774 16504 25780 16516
rect 24659 16476 25780 16504
rect 24659 16473 24671 16476
rect 24613 16467 24671 16473
rect 25774 16464 25780 16476
rect 25832 16464 25838 16516
rect 27246 16464 27252 16516
rect 27304 16464 27310 16516
rect 45186 16504 45192 16516
rect 45147 16476 45192 16504
rect 45186 16464 45192 16476
rect 45244 16464 45250 16516
rect 46658 16464 46664 16516
rect 46716 16504 46722 16516
rect 47397 16507 47455 16513
rect 47397 16504 47409 16507
rect 46716 16476 47409 16504
rect 46716 16464 46722 16476
rect 47397 16473 47409 16476
rect 47443 16473 47455 16507
rect 47397 16467 47455 16473
rect 22557 16439 22615 16445
rect 22557 16405 22569 16439
rect 22603 16436 22615 16439
rect 22922 16436 22928 16448
rect 22603 16408 22928 16436
rect 22603 16405 22615 16408
rect 22557 16399 22615 16405
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 27706 16436 27712 16448
rect 27667 16408 27712 16436
rect 27706 16396 27712 16408
rect 27764 16396 27770 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 17402 16192 17408 16244
rect 17460 16232 17466 16244
rect 45186 16232 45192 16244
rect 17460 16204 22094 16232
rect 45147 16204 45192 16232
rect 17460 16192 17466 16204
rect 22066 16164 22094 16204
rect 45186 16192 45192 16204
rect 45244 16192 45250 16244
rect 45462 16164 45468 16176
rect 22066 16136 45468 16164
rect 45462 16124 45468 16136
rect 45520 16124 45526 16176
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2087 16068 2774 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2746 15892 2774 16068
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 13504 16068 18521 16096
rect 13504 16056 13510 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 22738 16096 22744 16108
rect 22699 16068 22744 16096
rect 18509 16059 18567 16065
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 29733 16099 29791 16105
rect 29733 16096 29745 16099
rect 27764 16068 29745 16096
rect 27764 16056 27770 16068
rect 29733 16065 29745 16068
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 45097 16099 45155 16105
rect 45097 16065 45109 16099
rect 45143 16096 45155 16099
rect 45738 16096 45744 16108
rect 45143 16068 45744 16096
rect 45143 16065 45155 16068
rect 45097 16059 45155 16065
rect 45738 16056 45744 16068
rect 45796 16096 45802 16108
rect 46658 16096 46664 16108
rect 45796 16068 46664 16096
rect 45796 16056 45802 16068
rect 46658 16056 46664 16068
rect 46716 16056 46722 16108
rect 46750 16056 46756 16108
rect 46808 16096 46814 16108
rect 47765 16099 47823 16105
rect 47765 16096 47777 16099
rect 46808 16068 47777 16096
rect 46808 16056 46814 16068
rect 47765 16065 47777 16068
rect 47811 16065 47823 16099
rect 47765 16059 47823 16065
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 16028 18751 16031
rect 19334 16028 19340 16040
rect 18739 16000 19340 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 22922 16028 22928 16040
rect 22883 16000 22928 16028
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 24581 16031 24639 16037
rect 24581 15997 24593 16031
rect 24627 15997 24639 16031
rect 29914 16028 29920 16040
rect 29875 16000 29920 16028
rect 24581 15991 24639 15997
rect 24596 15960 24624 15991
rect 29914 15988 29920 16000
rect 29972 15988 29978 16040
rect 31386 16028 31392 16040
rect 31347 16000 31392 16028
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 45554 16028 45560 16040
rect 31726 16000 45560 16028
rect 31726 15960 31754 16000
rect 45554 15988 45560 16000
rect 45612 15988 45618 16040
rect 24596 15932 31754 15960
rect 2866 15892 2872 15904
rect 2746 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15892 2930 15904
rect 17770 15892 17776 15904
rect 2924 15864 17776 15892
rect 2924 15852 2930 15864
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 19334 15688 19340 15700
rect 19295 15660 19340 15688
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 29914 15688 29920 15700
rect 29875 15660 29920 15688
rect 29914 15648 29920 15660
rect 29972 15648 29978 15700
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15484 19303 15487
rect 19334 15484 19340 15496
rect 19291 15456 19340 15484
rect 19291 15453 19303 15456
rect 19245 15447 19303 15453
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 29822 15484 29828 15496
rect 29783 15456 29828 15484
rect 29822 15444 29828 15456
rect 29880 15484 29886 15496
rect 30190 15484 30196 15496
rect 29880 15456 30196 15484
rect 29880 15444 29886 15456
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 19392 14980 21005 15008
rect 19392 14968 19398 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2314 14940 2320 14952
rect 1995 14912 2320 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 21085 14807 21143 14813
rect 21085 14773 21097 14807
rect 21131 14804 21143 14807
rect 21726 14804 21732 14816
rect 21131 14776 21732 14804
rect 21131 14773 21143 14776
rect 21085 14767 21143 14773
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 21726 14464 21732 14476
rect 21687 14436 21732 14464
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 22646 14464 22652 14476
rect 22607 14436 22652 14464
rect 22646 14424 22652 14436
rect 22704 14424 22710 14476
rect 26697 14467 26755 14473
rect 26697 14433 26709 14467
rect 26743 14464 26755 14467
rect 27430 14464 27436 14476
rect 26743 14436 27436 14464
rect 26743 14433 26755 14436
rect 26697 14427 26755 14433
rect 27430 14424 27436 14436
rect 27488 14424 27494 14476
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 2188 14368 2237 14396
rect 2188 14356 2194 14368
rect 2225 14365 2237 14368
rect 2271 14396 2283 14399
rect 21085 14399 21143 14405
rect 2271 14368 2774 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2746 14260 2774 14368
rect 21085 14365 21097 14399
rect 21131 14396 21143 14399
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 21131 14368 21557 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 21545 14365 21557 14368
rect 21591 14365 21603 14399
rect 21545 14359 21603 14365
rect 26881 14331 26939 14337
rect 26881 14297 26893 14331
rect 26927 14328 26939 14331
rect 27062 14328 27068 14340
rect 26927 14300 27068 14328
rect 26927 14297 26939 14300
rect 26881 14291 26939 14297
rect 27062 14288 27068 14300
rect 27120 14288 27126 14340
rect 28442 14288 28448 14340
rect 28500 14328 28506 14340
rect 28537 14331 28595 14337
rect 28537 14328 28549 14331
rect 28500 14300 28549 14328
rect 28500 14288 28506 14300
rect 28537 14297 28549 14300
rect 28583 14297 28595 14331
rect 28537 14291 28595 14297
rect 34698 14260 34704 14272
rect 2746 14232 34704 14260
rect 34698 14220 34704 14232
rect 34756 14220 34762 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 27062 14056 27068 14068
rect 27023 14028 27068 14056
rect 27062 14016 27068 14028
rect 27120 14016 27126 14068
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 8803 13892 26985 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 26973 13889 26985 13892
rect 27019 13920 27031 13923
rect 29822 13920 29828 13932
rect 27019 13892 29828 13920
rect 27019 13889 27031 13892
rect 26973 13883 27031 13889
rect 29822 13880 29828 13892
rect 29880 13880 29886 13932
rect 46658 13920 46664 13932
rect 46619 13892 46664 13920
rect 46658 13880 46664 13892
rect 46716 13880 46722 13932
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8168 13824 8861 13852
rect 8168 13812 8174 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 10870 13716 10876 13728
rect 4028 13688 10876 13716
rect 4028 13676 4034 13688
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 46474 13676 46480 13728
rect 46532 13716 46538 13728
rect 46753 13719 46811 13725
rect 46753 13716 46765 13719
rect 46532 13688 46765 13716
rect 46532 13676 46538 13688
rect 46753 13685 46765 13688
rect 46799 13685 46811 13719
rect 46753 13679 46811 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 46474 13376 46480 13388
rect 46435 13348 46480 13376
rect 46474 13336 46480 13348
rect 46532 13336 46538 13388
rect 46290 13308 46296 13320
rect 46251 13280 46296 13308
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 46290 12792 46296 12844
rect 46348 12832 46354 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 46348 12804 47777 12832
rect 46348 12792 46354 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 32950 12628 32956 12640
rect 2179 12600 32956 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 32950 12588 32956 12600
rect 33008 12588 33014 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 47670 11064 47676 11076
rect 46523 11036 47676 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 47670 11024 47676 11036
rect 47728 11024 47734 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 15562 10996 15568 11008
rect 3200 10968 15568 10996
rect 3200 10956 3206 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 47670 10792 47676 10804
rect 47631 10764 47676 10792
rect 47670 10752 47676 10764
rect 47728 10752 47734 10804
rect 34698 10616 34704 10668
rect 34756 10656 34762 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 34756 10628 47593 10656
rect 34756 10616 34762 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47029 10455 47087 10461
rect 47029 10452 47041 10455
rect 46348 10424 47041 10452
rect 46348 10412 46354 10424
rect 47029 10421 47041 10424
rect 47075 10421 47087 10455
rect 47029 10415 47087 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 46477 9979 46535 9985
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 46934 9976 46940 9988
rect 46523 9948 46940 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 46934 9936 46940 9948
rect 46992 9936 46998 9988
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 46934 9636 46940 9648
rect 46895 9608 46940 9636
rect 46934 9596 46940 9608
rect 46992 9596 46998 9648
rect 45646 9528 45652 9580
rect 45704 9568 45710 9580
rect 46845 9571 46903 9577
rect 46845 9568 46857 9571
rect 45704 9540 46857 9568
rect 45704 9528 45710 9540
rect 46845 9537 46857 9540
rect 46891 9568 46903 9571
rect 47302 9568 47308 9580
rect 46891 9540 47308 9568
rect 46891 9537 46903 9540
rect 46845 9531 46903 9537
rect 47302 9528 47308 9540
rect 47360 9528 47366 9580
rect 47854 9568 47860 9580
rect 47815 9540 47860 9568
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 45830 9392 45836 9444
rect 45888 9432 45894 9444
rect 48041 9435 48099 9441
rect 48041 9432 48053 9435
rect 45888 9404 48053 9432
rect 45888 9392 45894 9404
rect 48041 9401 48053 9404
rect 48087 9401 48099 9435
rect 48041 9395 48099 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47854 8956 47860 8968
rect 47815 8928 47860 8956
rect 47854 8916 47860 8928
rect 47912 8916 47918 8968
rect 32214 8780 32220 8832
rect 32272 8820 32278 8832
rect 48041 8823 48099 8829
rect 48041 8820 48053 8823
rect 32272 8792 48053 8820
rect 32272 8780 32278 8792
rect 48041 8789 48053 8792
rect 48087 8789 48099 8823
rect 48041 8783 48099 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 46106 8480 46112 8492
rect 46067 8452 46112 8480
rect 46106 8440 46112 8452
rect 46164 8440 46170 8492
rect 2038 8304 2044 8356
rect 2096 8344 2102 8356
rect 2096 8316 45876 8344
rect 2096 8304 2102 8316
rect 39114 8236 39120 8288
rect 39172 8276 39178 8288
rect 45738 8276 45744 8288
rect 39172 8248 45744 8276
rect 39172 8236 39178 8248
rect 45738 8236 45744 8248
rect 45796 8236 45802 8288
rect 45848 8285 45876 8316
rect 45833 8279 45891 8285
rect 45833 8245 45845 8279
rect 45879 8276 45891 8279
rect 46201 8279 46259 8285
rect 46201 8276 46213 8279
rect 45879 8248 46213 8276
rect 45879 8245 45891 8248
rect 45833 8239 45891 8245
rect 46201 8245 46213 8248
rect 46247 8245 46259 8279
rect 46201 8239 46259 8245
rect 46382 8236 46388 8288
rect 46440 8276 46446 8288
rect 46569 8279 46627 8285
rect 46569 8276 46581 8279
rect 46440 8248 46581 8276
rect 46440 8236 46446 8248
rect 46569 8245 46581 8248
rect 46615 8245 46627 8279
rect 46569 8239 46627 8245
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 45922 7896 45928 7948
rect 45980 7936 45986 7948
rect 47213 7939 47271 7945
rect 47213 7936 47225 7939
rect 45980 7908 47225 7936
rect 45980 7896 45986 7908
rect 47213 7905 47225 7908
rect 47259 7905 47271 7939
rect 47213 7899 47271 7905
rect 46382 7868 46388 7880
rect 46343 7840 46388 7868
rect 46382 7828 46388 7840
rect 46440 7828 46446 7880
rect 46934 7800 46940 7812
rect 46895 7772 46940 7800
rect 46934 7760 46940 7772
rect 46992 7760 46998 7812
rect 47029 7803 47087 7809
rect 47029 7769 47041 7803
rect 47075 7769 47087 7803
rect 47029 7763 47087 7769
rect 46201 7735 46259 7741
rect 46201 7701 46213 7735
rect 46247 7732 46259 7735
rect 47044 7732 47072 7763
rect 46247 7704 47072 7732
rect 46247 7701 46259 7704
rect 46201 7695 46259 7701
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 46934 7488 46940 7540
rect 46992 7528 46998 7540
rect 47949 7531 48007 7537
rect 47949 7528 47961 7531
rect 46992 7500 47961 7528
rect 46992 7488 46998 7500
rect 47949 7497 47961 7500
rect 47995 7497 48007 7531
rect 47949 7491 48007 7497
rect 46106 7460 46112 7472
rect 46067 7432 46112 7460
rect 46106 7420 46112 7432
rect 46164 7420 46170 7472
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 46014 7324 46020 7336
rect 45975 7296 46020 7324
rect 46014 7284 46020 7296
rect 46072 7284 46078 7336
rect 46293 7327 46351 7333
rect 46293 7293 46305 7327
rect 46339 7293 46351 7327
rect 46293 7287 46351 7293
rect 45922 7216 45928 7268
rect 45980 7256 45986 7268
rect 46308 7256 46336 7287
rect 45980 7228 46336 7256
rect 45980 7216 45986 7228
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 28350 6848 28356 6860
rect 3476 6820 28356 6848
rect 3476 6808 3482 6820
rect 28350 6808 28356 6820
rect 28408 6808 28414 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47210 6740 47216 6792
rect 47268 6780 47274 6792
rect 47581 6783 47639 6789
rect 47581 6780 47593 6783
rect 47268 6752 47593 6780
rect 47268 6740 47274 6752
rect 47581 6749 47593 6752
rect 47627 6749 47639 6783
rect 47581 6743 47639 6749
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 48038 6440 48044 6452
rect 47999 6412 48044 6440
rect 48038 6400 48044 6412
rect 48096 6400 48102 6452
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 40126 5652 40132 5704
rect 40184 5692 40190 5704
rect 40221 5695 40279 5701
rect 40221 5692 40233 5695
rect 40184 5664 40233 5692
rect 40184 5652 40190 5664
rect 40221 5661 40233 5664
rect 40267 5661 40279 5695
rect 40221 5655 40279 5661
rect 40034 5516 40040 5568
rect 40092 5556 40098 5568
rect 40313 5559 40371 5565
rect 40313 5556 40325 5559
rect 40092 5528 40325 5556
rect 40092 5516 40098 5528
rect 40313 5525 40325 5528
rect 40359 5525 40371 5559
rect 40313 5519 40371 5525
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 37274 5352 37280 5364
rect 22066 5324 37280 5352
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 22066 5284 22094 5324
rect 37274 5312 37280 5324
rect 37332 5312 37338 5364
rect 37366 5312 37372 5364
rect 37424 5352 37430 5364
rect 38657 5355 38715 5361
rect 38657 5352 38669 5355
rect 37424 5324 38669 5352
rect 37424 5312 37430 5324
rect 38657 5321 38669 5324
rect 38703 5321 38715 5355
rect 48041 5355 48099 5361
rect 48041 5352 48053 5355
rect 38657 5315 38715 5321
rect 38764 5324 48053 5352
rect 4028 5256 22094 5284
rect 37461 5287 37519 5293
rect 4028 5244 4034 5256
rect 37461 5253 37473 5287
rect 37507 5284 37519 5287
rect 37550 5284 37556 5296
rect 37507 5256 37556 5284
rect 37507 5253 37519 5256
rect 37461 5247 37519 5253
rect 37550 5244 37556 5256
rect 37608 5244 37614 5296
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 20254 5216 20260 5228
rect 19659 5188 20260 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 23014 5216 23020 5228
rect 22603 5188 23020 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 23014 5176 23020 5188
rect 23072 5176 23078 5228
rect 23474 5216 23480 5228
rect 23435 5188 23480 5216
rect 23474 5176 23480 5188
rect 23532 5176 23538 5228
rect 37366 5148 37372 5160
rect 37327 5120 37372 5148
rect 37366 5108 37372 5120
rect 37424 5108 37430 5160
rect 38286 5148 38292 5160
rect 38247 5120 38292 5148
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 22649 5083 22707 5089
rect 22649 5049 22661 5083
rect 22695 5080 22707 5083
rect 23750 5080 23756 5092
rect 22695 5052 23756 5080
rect 22695 5049 22707 5052
rect 22649 5043 22707 5049
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 30098 5040 30104 5092
rect 30156 5080 30162 5092
rect 38764 5080 38792 5324
rect 48041 5321 48053 5324
rect 48087 5321 48099 5355
rect 48041 5315 48099 5321
rect 42334 5244 42340 5296
rect 42392 5284 42398 5296
rect 42613 5287 42671 5293
rect 42613 5284 42625 5287
rect 42392 5256 42625 5284
rect 42392 5244 42398 5256
rect 42613 5253 42625 5256
rect 42659 5253 42671 5287
rect 42613 5247 42671 5253
rect 40034 5216 40040 5228
rect 39995 5188 40040 5216
rect 40034 5176 40040 5188
rect 40092 5176 40098 5228
rect 43809 5219 43867 5225
rect 43809 5216 43821 5219
rect 43364 5188 43821 5216
rect 40218 5148 40224 5160
rect 40179 5120 40224 5148
rect 40218 5108 40224 5120
rect 40276 5108 40282 5160
rect 41874 5148 41880 5160
rect 41835 5120 41880 5148
rect 41874 5108 41880 5120
rect 41932 5108 41938 5160
rect 42521 5151 42579 5157
rect 42521 5148 42533 5151
rect 41984 5120 42533 5148
rect 30156 5052 38792 5080
rect 30156 5040 30162 5052
rect 19705 5015 19763 5021
rect 19705 4981 19717 5015
rect 19751 5012 19763 5015
rect 20070 5012 20076 5024
rect 19751 4984 20076 5012
rect 19751 4981 19763 4984
rect 19705 4975 19763 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 23293 5015 23351 5021
rect 23293 4981 23305 5015
rect 23339 5012 23351 5015
rect 24762 5012 24768 5024
rect 23339 4984 24768 5012
rect 23339 4981 23351 4984
rect 23293 4975 23351 4981
rect 24762 4972 24768 4984
rect 24820 4972 24826 5024
rect 37366 4972 37372 5024
rect 37424 5012 37430 5024
rect 41984 5012 42012 5120
rect 42521 5117 42533 5120
rect 42567 5148 42579 5151
rect 43364 5148 43392 5188
rect 43809 5185 43821 5188
rect 43855 5185 43867 5219
rect 43809 5179 43867 5185
rect 46750 5176 46756 5228
rect 46808 5216 46814 5228
rect 47857 5219 47915 5225
rect 47857 5216 47869 5219
rect 46808 5188 47869 5216
rect 46808 5176 46814 5188
rect 47857 5185 47869 5188
rect 47903 5185 47915 5219
rect 47857 5179 47915 5185
rect 42567 5120 43392 5148
rect 43533 5151 43591 5157
rect 42567 5117 42579 5120
rect 42521 5111 42579 5117
rect 43533 5117 43545 5151
rect 43579 5148 43591 5151
rect 43714 5148 43720 5160
rect 43579 5120 43720 5148
rect 43579 5117 43591 5120
rect 43533 5111 43591 5117
rect 43714 5108 43720 5120
rect 43772 5108 43778 5160
rect 37424 4984 42012 5012
rect 37424 4972 37430 4984
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 40218 4808 40224 4820
rect 40179 4780 40224 4808
rect 40218 4768 40224 4780
rect 40276 4768 40282 4820
rect 42334 4808 42340 4820
rect 42295 4780 42340 4808
rect 42334 4768 42340 4780
rect 42392 4768 42398 4820
rect 39209 4743 39267 4749
rect 39209 4709 39221 4743
rect 39255 4740 39267 4743
rect 40126 4740 40132 4752
rect 39255 4712 40132 4740
rect 39255 4709 39267 4712
rect 39209 4703 39267 4709
rect 40126 4700 40132 4712
rect 40184 4700 40190 4752
rect 46106 4700 46112 4752
rect 46164 4740 46170 4752
rect 46164 4712 47624 4740
rect 46164 4700 46170 4712
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 47486 4672 47492 4684
rect 21324 4644 23612 4672
rect 21324 4632 21330 4644
rect 19334 4604 19340 4616
rect 19295 4576 19340 4604
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 21634 4604 21640 4616
rect 21595 4576 21640 4604
rect 21634 4564 21640 4576
rect 21692 4564 21698 4616
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 22554 4604 22560 4616
rect 22327 4576 22560 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 23198 4604 23204 4616
rect 22971 4576 23204 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 23584 4613 23612 4644
rect 46676 4644 47492 4672
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 39117 4607 39175 4613
rect 39117 4573 39129 4607
rect 39163 4573 39175 4607
rect 40402 4604 40408 4616
rect 40363 4576 40408 4604
rect 39117 4567 39175 4573
rect 22186 4496 22192 4548
rect 22244 4536 22250 4548
rect 23017 4539 23075 4545
rect 23017 4536 23029 4539
rect 22244 4508 23029 4536
rect 22244 4496 22250 4508
rect 23017 4505 23029 4508
rect 23063 4505 23075 4539
rect 39132 4536 39160 4567
rect 40402 4564 40408 4576
rect 40460 4564 40466 4616
rect 40770 4564 40776 4616
rect 40828 4604 40834 4616
rect 40865 4607 40923 4613
rect 40865 4604 40877 4607
rect 40828 4576 40877 4604
rect 40828 4564 40834 4576
rect 40865 4573 40877 4576
rect 40911 4573 40923 4607
rect 40865 4567 40923 4573
rect 40957 4607 41015 4613
rect 40957 4573 40969 4607
rect 41003 4604 41015 4607
rect 41509 4607 41567 4613
rect 41509 4604 41521 4607
rect 41003 4576 41521 4604
rect 41003 4573 41015 4576
rect 40957 4567 41015 4573
rect 41509 4573 41521 4576
rect 41555 4573 41567 4607
rect 41509 4567 41567 4573
rect 42521 4607 42579 4613
rect 42521 4573 42533 4607
rect 42567 4604 42579 4607
rect 42886 4604 42892 4616
rect 42567 4576 42892 4604
rect 42567 4573 42579 4576
rect 42521 4567 42579 4573
rect 42886 4564 42892 4576
rect 42944 4564 42950 4616
rect 46676 4613 46704 4644
rect 47486 4632 47492 4644
rect 47544 4632 47550 4684
rect 47596 4681 47624 4712
rect 47581 4675 47639 4681
rect 47581 4641 47593 4675
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 46661 4607 46719 4613
rect 46661 4573 46673 4607
rect 46707 4573 46719 4607
rect 46661 4567 46719 4573
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47305 4607 47363 4613
rect 47305 4604 47317 4607
rect 46900 4576 47317 4604
rect 46900 4564 46906 4576
rect 47305 4573 47317 4576
rect 47351 4573 47363 4607
rect 47305 4567 47363 4573
rect 41601 4539 41659 4545
rect 41601 4536 41613 4539
rect 39132 4508 41613 4536
rect 23017 4499 23075 4505
rect 41601 4505 41613 4508
rect 41647 4505 41659 4539
rect 41601 4499 41659 4505
rect 19426 4468 19432 4480
rect 19387 4440 19432 4468
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 20441 4471 20499 4477
rect 20441 4437 20453 4471
rect 20487 4468 20499 4471
rect 20622 4468 20628 4480
rect 20487 4440 20628 4468
rect 20487 4437 20499 4440
rect 20441 4431 20499 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21082 4468 21088 4480
rect 21043 4440 21088 4468
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22278 4468 22284 4480
rect 21775 4440 22284 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 22373 4471 22431 4477
rect 22373 4437 22385 4471
rect 22419 4468 22431 4471
rect 22462 4468 22468 4480
rect 22419 4440 22468 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 23290 4428 23296 4480
rect 23348 4468 23354 4480
rect 23661 4471 23719 4477
rect 23661 4468 23673 4471
rect 23348 4440 23673 4468
rect 23348 4428 23354 4440
rect 23661 4437 23673 4440
rect 23707 4437 23719 4471
rect 23661 4431 23719 4437
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46753 4471 46811 4477
rect 46753 4468 46765 4471
rect 46532 4440 46765 4468
rect 46532 4428 46538 4440
rect 46753 4437 46765 4440
rect 46799 4437 46811 4471
rect 46753 4431 46811 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 20717 4267 20775 4273
rect 19720 4236 20208 4264
rect 7392 4168 7604 4196
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2774 4128 2780 4140
rect 2735 4100 2780 4128
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 7392 4060 7420 4168
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 3476 4032 7420 4060
rect 3476 4020 3482 4032
rect 7484 3992 7512 4091
rect 7576 4060 7604 4168
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 17862 4128 17868 4140
rect 10091 4100 17868 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 18380 4100 18613 4128
rect 18380 4088 18386 4100
rect 18601 4097 18613 4100
rect 18647 4097 18659 4131
rect 19242 4128 19248 4140
rect 19203 4100 19248 4128
rect 18601 4091 18659 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19720 4060 19748 4236
rect 19794 4156 19800 4208
rect 19852 4196 19858 4208
rect 20073 4199 20131 4205
rect 20073 4196 20085 4199
rect 19852 4168 20085 4196
rect 19852 4156 19858 4168
rect 20073 4165 20085 4168
rect 20119 4165 20131 4199
rect 20180 4196 20208 4236
rect 20717 4233 20729 4267
rect 20763 4264 20775 4267
rect 20990 4264 20996 4276
rect 20763 4236 20996 4264
rect 20763 4233 20775 4236
rect 20717 4227 20775 4233
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21692 4236 21925 4264
rect 21692 4224 21698 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 22554 4264 22560 4276
rect 22515 4236 22560 4264
rect 21913 4227 21971 4233
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 37277 4267 37335 4273
rect 37277 4233 37289 4267
rect 37323 4264 37335 4267
rect 37550 4264 37556 4276
rect 37323 4236 37556 4264
rect 37323 4233 37335 4236
rect 37277 4227 37335 4233
rect 37550 4224 37556 4236
rect 37608 4224 37614 4276
rect 40402 4224 40408 4276
rect 40460 4264 40466 4276
rect 40865 4267 40923 4273
rect 40865 4264 40877 4267
rect 40460 4236 40877 4264
rect 40460 4224 40466 4236
rect 40865 4233 40877 4236
rect 40911 4233 40923 4267
rect 40865 4227 40923 4233
rect 22370 4196 22376 4208
rect 20180 4168 22376 4196
rect 20073 4159 20131 4165
rect 22370 4156 22376 4168
rect 22428 4156 22434 4208
rect 25409 4199 25467 4205
rect 25409 4196 25421 4199
rect 25240 4168 25421 4196
rect 25240 4140 25268 4168
rect 25409 4165 25421 4168
rect 25455 4165 25467 4199
rect 25409 4159 25467 4165
rect 25501 4199 25559 4205
rect 25501 4165 25513 4199
rect 25547 4196 25559 4199
rect 25590 4196 25596 4208
rect 25547 4168 25596 4196
rect 25547 4165 25559 4168
rect 25501 4159 25559 4165
rect 25590 4156 25596 4168
rect 25648 4156 25654 4208
rect 40037 4199 40095 4205
rect 40037 4165 40049 4199
rect 40083 4196 40095 4199
rect 40770 4196 40776 4208
rect 40083 4168 40776 4196
rect 40083 4165 40095 4168
rect 40037 4159 40095 4165
rect 40770 4156 40776 4168
rect 40828 4156 40834 4208
rect 42797 4199 42855 4205
rect 42797 4165 42809 4199
rect 42843 4196 42855 4199
rect 43254 4196 43260 4208
rect 42843 4168 43260 4196
rect 42843 4165 42855 4168
rect 42797 4159 42855 4165
rect 43254 4156 43260 4168
rect 43312 4156 43318 4208
rect 43714 4196 43720 4208
rect 43675 4168 43720 4196
rect 43714 4156 43720 4168
rect 43772 4156 43778 4208
rect 46658 4196 46664 4208
rect 46619 4168 46664 4196
rect 46658 4156 46664 4168
rect 46716 4156 46722 4208
rect 47765 4199 47823 4205
rect 47765 4165 47777 4199
rect 47811 4196 47823 4199
rect 47854 4196 47860 4208
rect 47811 4168 47860 4196
rect 47811 4165 47823 4168
rect 47765 4159 47823 4165
rect 47854 4156 47860 4168
rect 47912 4156 47918 4208
rect 19978 4128 19984 4140
rect 19939 4100 19984 4128
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20622 4128 20628 4140
rect 20583 4100 20628 4128
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21082 4088 21088 4140
rect 21140 4128 21146 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21140 4100 21833 4128
rect 21140 4088 21146 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 22336 4100 22477 4128
rect 22336 4088 22342 4100
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 23109 4131 23167 4137
rect 23109 4128 23121 4131
rect 22612 4100 23121 4128
rect 22612 4088 22618 4100
rect 23109 4097 23121 4100
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 23382 4088 23388 4140
rect 23440 4128 23446 4140
rect 23753 4131 23811 4137
rect 23753 4128 23765 4131
rect 23440 4100 23765 4128
rect 23440 4088 23446 4100
rect 23753 4097 23765 4100
rect 23799 4097 23811 4131
rect 23753 4091 23811 4097
rect 24320 4100 24900 4128
rect 7576 4032 19748 4060
rect 19904 4032 20852 4060
rect 19904 3992 19932 4032
rect 7484 3964 19932 3992
rect 20824 3992 20852 4032
rect 20898 4020 20904 4072
rect 20956 4060 20962 4072
rect 24320 4060 24348 4100
rect 20956 4032 24348 4060
rect 20956 4020 20962 4032
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 24872 4060 24900 4100
rect 25222 4088 25228 4140
rect 25280 4088 25286 4140
rect 28810 4128 28816 4140
rect 26252 4100 28816 4128
rect 26252 4060 26280 4100
rect 28810 4088 28816 4100
rect 28868 4088 28874 4140
rect 30101 4131 30159 4137
rect 30101 4097 30113 4131
rect 30147 4128 30159 4131
rect 30926 4128 30932 4140
rect 30147 4100 30932 4128
rect 30147 4097 30159 4100
rect 30101 4091 30159 4097
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 37461 4131 37519 4137
rect 37461 4097 37473 4131
rect 37507 4128 37519 4131
rect 37734 4128 37740 4140
rect 37507 4100 37740 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 37734 4088 37740 4100
rect 37792 4088 37798 4140
rect 40494 4128 40500 4140
rect 39592 4100 40356 4128
rect 40455 4100 40500 4128
rect 39592 4072 39620 4100
rect 24452 4032 24808 4060
rect 24872 4032 26280 4060
rect 26421 4063 26479 4069
rect 24452 4020 24458 4032
rect 24670 3992 24676 4004
rect 20824 3964 24676 3992
rect 24670 3952 24676 3964
rect 24728 3952 24734 4004
rect 24780 3992 24808 4032
rect 26421 4029 26433 4063
rect 26467 4060 26479 4063
rect 26602 4060 26608 4072
rect 26467 4032 26608 4060
rect 26467 4029 26479 4032
rect 26421 4023 26479 4029
rect 26602 4020 26608 4032
rect 26660 4060 26666 4072
rect 28534 4060 28540 4072
rect 26660 4032 28540 4060
rect 26660 4020 26666 4032
rect 28534 4020 28540 4032
rect 28592 4020 28598 4072
rect 39390 4060 39396 4072
rect 39351 4032 39396 4060
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 39574 4060 39580 4072
rect 39535 4032 39580 4060
rect 39574 4020 39580 4032
rect 39632 4020 39638 4072
rect 40218 4060 40224 4072
rect 39960 4032 40224 4060
rect 30193 3995 30251 4001
rect 30193 3992 30205 3995
rect 24780 3964 30205 3992
rect 30193 3961 30205 3964
rect 30239 3961 30251 3995
rect 39960 3992 39988 4032
rect 40218 4020 40224 4032
rect 40276 4020 40282 4072
rect 40328 4060 40356 4100
rect 40494 4088 40500 4100
rect 40552 4088 40558 4140
rect 40681 4131 40739 4137
rect 40681 4097 40693 4131
rect 40727 4097 40739 4131
rect 46014 4128 46020 4140
rect 40681 4091 40739 4097
rect 43640 4100 46020 4128
rect 40696 4060 40724 4091
rect 40328 4032 40724 4060
rect 40770 4020 40776 4072
rect 40828 4060 40834 4072
rect 42705 4063 42763 4069
rect 42705 4060 42717 4063
rect 40828 4032 42717 4060
rect 40828 4020 40834 4032
rect 42705 4029 42717 4032
rect 42751 4060 42763 4063
rect 43640 4060 43668 4100
rect 46014 4088 46020 4100
rect 46072 4088 46078 4140
rect 42751 4032 43668 4060
rect 42751 4029 42763 4032
rect 42705 4023 42763 4029
rect 43714 4020 43720 4072
rect 43772 4060 43778 4072
rect 48041 4063 48099 4069
rect 48041 4060 48053 4063
rect 43772 4032 48053 4060
rect 43772 4020 43778 4032
rect 48041 4029 48053 4032
rect 48087 4029 48099 4063
rect 48041 4023 48099 4029
rect 46845 3995 46903 4001
rect 46845 3992 46857 3995
rect 30193 3955 30251 3961
rect 30300 3964 39988 3992
rect 40236 3964 43668 3992
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2004 3896 2237 3924
rect 2004 3884 2010 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6604 3896 6837 3924
rect 6604 3884 6610 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 7558 3924 7564 3936
rect 7519 3896 7564 3924
rect 6825 3887 6883 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7984 3896 8309 3924
rect 7984 3884 7990 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9364 3896 9505 3924
rect 9364 3884 9370 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 10134 3924 10140 3936
rect 10095 3896 10140 3924
rect 9493 3887 9551 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11572 3896 11713 3924
rect 11572 3884 11578 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 17644 3896 18705 3924
rect 17644 3884 17650 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19337 3927 19395 3933
rect 19337 3924 19349 3927
rect 18932 3896 19349 3924
rect 18932 3884 18938 3896
rect 19337 3893 19349 3896
rect 19383 3893 19395 3927
rect 19337 3887 19395 3893
rect 23106 3884 23112 3936
rect 23164 3924 23170 3936
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 23164 3896 23213 3924
rect 23164 3884 23170 3896
rect 23201 3893 23213 3896
rect 23247 3893 23259 3927
rect 23842 3924 23848 3936
rect 23803 3896 23848 3924
rect 23201 3887 23259 3893
rect 23842 3884 23848 3896
rect 23900 3884 23906 3936
rect 24578 3884 24584 3936
rect 24636 3924 24642 3936
rect 24857 3927 24915 3933
rect 24857 3924 24869 3927
rect 24636 3896 24869 3924
rect 24636 3884 24642 3896
rect 24857 3893 24869 3896
rect 24903 3893 24915 3927
rect 24857 3887 24915 3893
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 30300 3924 30328 3964
rect 25372 3896 30328 3924
rect 25372 3884 25378 3896
rect 30374 3884 30380 3936
rect 30432 3924 30438 3936
rect 40236 3924 40264 3964
rect 30432 3896 40264 3924
rect 30432 3884 30438 3896
rect 40310 3884 40316 3936
rect 40368 3924 40374 3936
rect 43530 3924 43536 3936
rect 40368 3896 43536 3924
rect 40368 3884 40374 3896
rect 43530 3884 43536 3896
rect 43588 3884 43594 3936
rect 43640 3924 43668 3964
rect 45526 3964 46857 3992
rect 45526 3924 45554 3964
rect 46845 3961 46857 3964
rect 46891 3961 46903 3995
rect 46845 3955 46903 3961
rect 43640 3896 45554 3924
rect 46109 3927 46167 3933
rect 46109 3893 46121 3927
rect 46155 3924 46167 3927
rect 46290 3924 46296 3936
rect 46155 3896 46296 3924
rect 46155 3893 46167 3896
rect 46109 3887 46167 3893
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 17681 3723 17739 3729
rect 17681 3689 17693 3723
rect 17727 3720 17739 3723
rect 19242 3720 19248 3732
rect 17727 3692 19248 3720
rect 17727 3689 17739 3692
rect 17681 3683 17739 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19613 3723 19671 3729
rect 19613 3689 19625 3723
rect 19659 3720 19671 3723
rect 20346 3720 20352 3732
rect 19659 3692 20352 3720
rect 19659 3689 19671 3692
rect 19613 3683 19671 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 35526 3720 35532 3732
rect 22066 3692 35532 3720
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 22066 3652 22094 3692
rect 35526 3680 35532 3692
rect 35584 3680 35590 3732
rect 40313 3723 40371 3729
rect 35866 3692 40172 3720
rect 22554 3652 22560 3664
rect 3936 3624 22094 3652
rect 22515 3624 22560 3652
rect 3936 3612 3942 3624
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 23198 3652 23204 3664
rect 23159 3624 23204 3652
rect 23198 3612 23204 3624
rect 23256 3612 23262 3664
rect 30374 3652 30380 3664
rect 24688 3624 30380 3652
rect 7098 3584 7104 3596
rect 7059 3556 7104 3584
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 10134 3584 10140 3596
rect 9539 3556 10140 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3553 10747 3587
rect 10689 3547 10747 3553
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 1820 3488 2881 3516
rect 1820 3476 1826 3488
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 2869 3479 2927 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6135 3488 6561 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1360 3420 1869 3448
rect 1360 3408 1366 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 6730 3448 6736 3460
rect 6691 3420 6736 3448
rect 1857 3411 1915 3417
rect 6730 3408 6736 3420
rect 6788 3408 6794 3460
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 10704 3448 10732 3547
rect 20438 3544 20444 3596
rect 20496 3584 20502 3596
rect 20625 3587 20683 3593
rect 20625 3584 20637 3587
rect 20496 3556 20637 3584
rect 20496 3544 20502 3556
rect 20625 3553 20637 3556
rect 20671 3553 20683 3587
rect 20625 3547 20683 3553
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 24688 3584 24716 3624
rect 30374 3612 30380 3624
rect 30432 3612 30438 3664
rect 35866 3652 35894 3692
rect 39390 3652 39396 3664
rect 31726 3624 35894 3652
rect 37660 3624 39396 3652
rect 20864 3556 24716 3584
rect 20864 3544 20870 3556
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 25593 3587 25651 3593
rect 25593 3584 25605 3587
rect 24820 3556 25605 3584
rect 24820 3544 24826 3556
rect 25593 3553 25605 3556
rect 25639 3553 25651 3587
rect 26602 3584 26608 3596
rect 26563 3556 26608 3584
rect 25593 3547 25651 3553
rect 26602 3544 26608 3556
rect 26660 3544 26666 3596
rect 12066 3516 12072 3528
rect 12027 3488 12072 3516
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 17586 3516 17592 3528
rect 17547 3488 17592 3516
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17828 3488 18245 3516
rect 17828 3476 17834 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3516 19579 3519
rect 19794 3516 19800 3528
rect 19567 3488 19800 3516
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 22462 3516 22468 3528
rect 22423 3488 22468 3516
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 23106 3516 23112 3528
rect 23067 3488 23112 3516
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27249 3519 27307 3525
rect 27249 3516 27261 3519
rect 26752 3488 27261 3516
rect 26752 3476 26758 3488
rect 27249 3485 27261 3488
rect 27295 3485 27307 3519
rect 27249 3479 27307 3485
rect 27338 3476 27344 3528
rect 27396 3516 27402 3528
rect 31726 3516 31754 3624
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 37274 3584 37280 3596
rect 35492 3556 37280 3584
rect 35492 3544 35498 3556
rect 37274 3544 37280 3556
rect 37332 3544 37338 3596
rect 37660 3593 37688 3624
rect 39390 3612 39396 3624
rect 39448 3612 39454 3664
rect 40144 3652 40172 3692
rect 40313 3689 40325 3723
rect 40359 3720 40371 3723
rect 40494 3720 40500 3732
rect 40359 3692 40500 3720
rect 40359 3689 40371 3692
rect 40313 3683 40371 3689
rect 40494 3680 40500 3692
rect 40552 3680 40558 3732
rect 44266 3652 44272 3664
rect 40144 3624 44272 3652
rect 44266 3612 44272 3624
rect 44324 3612 44330 3664
rect 37645 3587 37703 3593
rect 37645 3584 37657 3587
rect 37476 3556 37657 3584
rect 32950 3516 32956 3528
rect 27396 3488 31754 3516
rect 32911 3488 32956 3516
rect 27396 3476 27402 3488
rect 32950 3476 32956 3488
rect 33008 3476 33014 3528
rect 33778 3516 33784 3528
rect 33739 3488 33784 3516
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 20346 3448 20352 3460
rect 9088 3420 10732 3448
rect 11624 3420 18460 3448
rect 20307 3420 20352 3448
rect 9088 3408 9094 3420
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 11624 3380 11652 3420
rect 2179 3352 11652 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12161 3383 12219 3389
rect 12161 3380 12173 3383
rect 11756 3352 12173 3380
rect 11756 3340 11762 3352
rect 12161 3349 12173 3352
rect 12207 3349 12219 3383
rect 12161 3343 12219 3349
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 14056 3352 14197 3380
rect 14056 3340 14062 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 18325 3383 18383 3389
rect 18325 3380 18337 3383
rect 18288 3352 18337 3380
rect 18288 3340 18294 3352
rect 18325 3349 18337 3352
rect 18371 3349 18383 3383
rect 18432 3380 18460 3420
rect 20346 3408 20352 3420
rect 20404 3408 20410 3460
rect 25694 3451 25752 3457
rect 25694 3417 25706 3451
rect 25740 3448 25752 3451
rect 25740 3420 25820 3448
rect 25740 3417 25752 3420
rect 25694 3411 25752 3417
rect 20898 3380 20904 3392
rect 18432 3352 20904 3380
rect 18325 3343 18383 3349
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 24486 3380 24492 3392
rect 21968 3352 24492 3380
rect 21968 3340 21974 3352
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25792 3380 25820 3420
rect 30006 3408 30012 3460
rect 30064 3448 30070 3460
rect 37476 3448 37504 3556
rect 37645 3553 37657 3556
rect 37691 3553 37703 3587
rect 38286 3584 38292 3596
rect 38247 3556 38292 3584
rect 37645 3547 37703 3553
rect 38286 3544 38292 3556
rect 38344 3544 38350 3596
rect 40221 3587 40279 3593
rect 40221 3553 40233 3587
rect 40267 3584 40279 3587
rect 41690 3584 41696 3596
rect 40267 3556 41696 3584
rect 40267 3553 40279 3556
rect 40221 3547 40279 3553
rect 41690 3544 41696 3556
rect 41748 3544 41754 3596
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 42794 3544 42800 3596
rect 42852 3584 42858 3596
rect 44085 3587 44143 3593
rect 44085 3584 44097 3587
rect 42852 3556 44097 3584
rect 42852 3544 42858 3556
rect 44085 3553 44097 3556
rect 44131 3553 44143 3587
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 44085 3547 44143 3553
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 39114 3476 39120 3528
rect 39172 3516 39178 3528
rect 39574 3516 39580 3528
rect 39172 3488 39580 3516
rect 39172 3476 39178 3488
rect 39574 3476 39580 3488
rect 39632 3516 39638 3528
rect 39945 3519 40003 3525
rect 39945 3516 39957 3519
rect 39632 3488 39957 3516
rect 39632 3476 39638 3488
rect 39945 3485 39957 3488
rect 39991 3485 40003 3519
rect 40954 3516 40960 3528
rect 40915 3488 40960 3516
rect 39945 3479 40003 3485
rect 40954 3476 40960 3488
rect 41012 3476 41018 3528
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 42760 3488 43269 3516
rect 42760 3476 42766 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 43257 3479 43315 3485
rect 30064 3420 37504 3448
rect 37737 3451 37795 3457
rect 30064 3408 30070 3420
rect 37737 3417 37749 3451
rect 37783 3448 37795 3451
rect 38654 3448 38660 3460
rect 37783 3420 38660 3448
rect 37783 3417 37795 3420
rect 37737 3411 37795 3417
rect 38654 3408 38660 3420
rect 38712 3408 38718 3460
rect 39758 3408 39764 3460
rect 39816 3448 39822 3460
rect 41141 3451 41199 3457
rect 41141 3448 41153 3451
rect 39816 3420 41153 3448
rect 39816 3408 39822 3420
rect 41141 3417 41153 3420
rect 41187 3417 41199 3451
rect 43272 3448 43300 3479
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45646 3516 45652 3528
rect 45607 3488 45652 3516
rect 45646 3476 45652 3488
rect 45704 3476 45710 3528
rect 46198 3448 46204 3460
rect 43272 3420 46204 3448
rect 41141 3411 41199 3417
rect 46198 3408 46204 3420
rect 46256 3408 46262 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 27065 3383 27123 3389
rect 27065 3380 27077 3383
rect 25792 3352 27077 3380
rect 27065 3349 27077 3352
rect 27111 3349 27123 3383
rect 27065 3343 27123 3349
rect 33045 3383 33103 3389
rect 33045 3349 33057 3383
rect 33091 3380 33103 3383
rect 33134 3380 33140 3392
rect 33091 3352 33140 3380
rect 33091 3349 33103 3352
rect 33045 3343 33103 3349
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 39942 3340 39948 3392
rect 40000 3380 40006 3392
rect 40497 3383 40555 3389
rect 40497 3380 40509 3383
rect 40000 3352 40509 3380
rect 40000 3340 40006 3352
rect 40497 3349 40509 3352
rect 40543 3349 40555 3383
rect 40497 3343 40555 3349
rect 42978 3340 42984 3392
rect 43036 3380 43042 3392
rect 43349 3383 43407 3389
rect 43349 3380 43361 3383
rect 43036 3352 43361 3380
rect 43036 3340 43042 3352
rect 43349 3349 43361 3352
rect 43395 3349 43407 3383
rect 43349 3343 43407 3349
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 6730 3176 6736 3188
rect 6691 3148 6736 3176
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 14090 3176 14096 3188
rect 6886 3148 14096 3176
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 6638 3040 6644 3052
rect 6551 3012 6644 3040
rect 6638 3000 6644 3012
rect 6696 3040 6702 3052
rect 6886 3040 6914 3148
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 18322 3176 18328 3188
rect 18283 3148 18328 3176
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 18969 3179 19027 3185
rect 18969 3145 18981 3179
rect 19015 3176 19027 3179
rect 19334 3176 19340 3188
rect 19015 3148 19340 3176
rect 19015 3145 19027 3148
rect 18969 3139 19027 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 24394 3176 24400 3188
rect 20404 3148 24400 3176
rect 20404 3136 20410 3148
rect 24394 3136 24400 3148
rect 24452 3136 24458 3188
rect 24486 3136 24492 3188
rect 24544 3176 24550 3188
rect 33778 3176 33784 3188
rect 24544 3148 31754 3176
rect 24544 3136 24550 3148
rect 8110 3108 8116 3120
rect 8071 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13998 3108 14004 3120
rect 13959 3080 14004 3108
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 18690 3108 18696 3120
rect 17420 3080 18696 3108
rect 7926 3040 7932 3052
rect 6696 3012 6914 3040
rect 7887 3012 7932 3040
rect 6696 3000 6702 3012
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 17420 3049 17448 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 21177 3111 21235 3117
rect 21177 3077 21189 3111
rect 21223 3108 21235 3111
rect 23382 3108 23388 3120
rect 21223 3080 23388 3108
rect 21223 3077 21235 3080
rect 21177 3071 21235 3077
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 24762 3108 24768 3120
rect 24723 3080 24768 3108
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 25222 3108 25228 3120
rect 24912 3080 25228 3108
rect 24912 3068 24918 3080
rect 25222 3068 25228 3080
rect 25280 3108 25286 3120
rect 30006 3108 30012 3120
rect 25280 3080 30012 3108
rect 25280 3068 25286 3080
rect 30006 3068 30012 3080
rect 30064 3068 30070 3120
rect 31726 3108 31754 3148
rect 32968 3148 33784 3176
rect 32214 3108 32220 3120
rect 31726 3080 32220 3108
rect 32214 3068 32220 3080
rect 32272 3068 32278 3120
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 18230 3040 18236 3052
rect 18191 3012 18236 3040
rect 17405 3003 17463 3009
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 18874 3040 18880 3052
rect 18835 3012 18880 3040
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7800 2944 8401 2972
rect 7800 2932 7806 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11020 2944 11989 2972
rect 11020 2932 11026 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15252 2944 17325 2972
rect 15252 2932 15258 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17770 2972 17776 2984
rect 17731 2944 17776 2972
rect 17313 2935 17371 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 19536 2972 19564 3003
rect 20162 3000 20168 3052
rect 20220 3040 20226 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20220 3012 20361 3040
rect 20220 3000 20226 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3040 21143 3043
rect 22186 3040 22192 3052
rect 21131 3012 22192 3040
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22370 3040 22376 3052
rect 22331 3012 22376 3040
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3040 23167 3043
rect 23290 3040 23296 3052
rect 23155 3012 23296 3040
rect 23155 3009 23167 3012
rect 23109 3003 23167 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23750 3040 23756 3052
rect 23711 3012 23756 3040
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 32968 3049 32996 3148
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 37734 3176 37740 3188
rect 37695 3148 37740 3176
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 39758 3176 39764 3188
rect 39719 3148 39764 3176
rect 39758 3136 39764 3148
rect 39816 3136 39822 3188
rect 40954 3136 40960 3188
rect 41012 3176 41018 3188
rect 41049 3179 41107 3185
rect 41049 3176 41061 3179
rect 41012 3148 41061 3176
rect 41012 3136 41018 3148
rect 41049 3145 41061 3148
rect 41095 3145 41107 3179
rect 41049 3139 41107 3145
rect 47762 3136 47768 3188
rect 47820 3176 47826 3188
rect 47857 3179 47915 3185
rect 47857 3176 47869 3179
rect 47820 3148 47869 3176
rect 47820 3136 47826 3148
rect 47857 3145 47869 3148
rect 47903 3145 47915 3179
rect 47857 3139 47915 3145
rect 33134 3108 33140 3120
rect 33095 3080 33140 3108
rect 33134 3068 33140 3080
rect 33192 3068 33198 3120
rect 42702 3108 42708 3120
rect 35866 3080 42708 3108
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 27120 3012 27169 3040
rect 27120 3000 27126 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 32953 3043 33011 3049
rect 32953 3009 32965 3043
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 22002 2972 22008 2984
rect 19536 2944 22008 2972
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 23017 2975 23075 2981
rect 23017 2941 23029 2975
rect 23063 2972 23075 2975
rect 24854 2972 24860 2984
rect 23063 2944 24860 2972
rect 23063 2941 23075 2944
rect 23017 2935 23075 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 12124 2876 31754 2904
rect 12124 2864 12130 2876
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 18690 2836 18696 2848
rect 13412 2808 18696 2836
rect 13412 2796 13418 2808
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19613 2839 19671 2845
rect 19613 2805 19625 2839
rect 19659 2836 19671 2839
rect 21266 2836 21272 2848
rect 19659 2808 21272 2836
rect 19659 2805 19671 2808
rect 19613 2799 19671 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 23566 2796 23572 2848
rect 23624 2836 23630 2848
rect 23845 2839 23903 2845
rect 23845 2836 23857 2839
rect 23624 2808 23857 2836
rect 23624 2796 23630 2808
rect 23845 2805 23857 2808
rect 23891 2805 23903 2839
rect 23845 2799 23903 2805
rect 27341 2839 27399 2845
rect 27341 2805 27353 2839
rect 27387 2836 27399 2839
rect 31294 2836 31300 2848
rect 27387 2808 31300 2836
rect 27387 2805 27399 2808
rect 27341 2799 27399 2805
rect 31294 2796 31300 2808
rect 31352 2796 31358 2848
rect 31726 2836 31754 2876
rect 32950 2836 32956 2848
rect 31726 2808 32956 2836
rect 32950 2796 32956 2808
rect 33008 2836 33014 2848
rect 35866 2836 35894 3080
rect 42702 3068 42708 3080
rect 42760 3068 42766 3120
rect 42978 3108 42984 3120
rect 42939 3080 42984 3108
rect 42978 3068 42984 3080
rect 43036 3068 43042 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 38654 3040 38660 3052
rect 37323 3012 38660 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 38654 3000 38660 3012
rect 38712 3000 38718 3052
rect 39942 3040 39948 3052
rect 39903 3012 39948 3040
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 40405 3043 40463 3049
rect 40405 3009 40417 3043
rect 40451 3040 40463 3043
rect 40770 3040 40776 3052
rect 40451 3012 40776 3040
rect 40451 3009 40463 3012
rect 40405 3003 40463 3009
rect 39390 2932 39396 2984
rect 39448 2972 39454 2984
rect 40420 2972 40448 3003
rect 40770 3000 40776 3012
rect 40828 3000 40834 3052
rect 42794 3040 42800 3052
rect 42755 3012 42800 3040
rect 42794 3000 42800 3012
rect 42852 3000 42858 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3040 47823 3043
rect 48314 3040 48320 3052
rect 47811 3012 48320 3040
rect 47811 3009 47823 3012
rect 47765 3003 47823 3009
rect 48314 3000 48320 3012
rect 48372 3000 48378 3052
rect 39448 2944 40448 2972
rect 40589 2975 40647 2981
rect 39448 2932 39454 2944
rect 40589 2941 40601 2975
rect 40635 2972 40647 2975
rect 41690 2972 41696 2984
rect 40635 2944 41696 2972
rect 40635 2941 40647 2944
rect 40589 2935 40647 2941
rect 41690 2932 41696 2944
rect 41748 2932 41754 2984
rect 43162 2932 43168 2984
rect 43220 2972 43226 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 43220 2944 43269 2972
rect 43220 2932 43226 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 37274 2864 37280 2916
rect 37332 2904 37338 2916
rect 45094 2904 45100 2916
rect 37332 2876 45100 2904
rect 37332 2864 37338 2876
rect 45094 2864 45100 2876
rect 45152 2864 45158 2916
rect 37366 2836 37372 2848
rect 33008 2808 35894 2836
rect 37327 2808 37372 2836
rect 33008 2796 33014 2808
rect 37366 2796 37372 2808
rect 37424 2796 37430 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 19978 2632 19984 2644
rect 19939 2604 19984 2632
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20530 2592 20536 2644
rect 20588 2632 20594 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20588 2604 20913 2632
rect 20588 2592 20594 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 22370 2632 22376 2644
rect 22331 2604 22376 2632
rect 20901 2595 20959 2601
rect 22370 2592 22376 2604
rect 22428 2592 22434 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 25961 2635 26019 2641
rect 25961 2601 25973 2635
rect 26007 2632 26019 2635
rect 28074 2632 28080 2644
rect 26007 2604 28080 2632
rect 26007 2601 26019 2604
rect 25961 2595 26019 2601
rect 28074 2592 28080 2604
rect 28132 2592 28138 2644
rect 28166 2592 28172 2644
rect 28224 2632 28230 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 28224 2604 28641 2632
rect 28224 2592 28230 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 28629 2595 28687 2601
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 30340 2604 35572 2632
rect 30340 2592 30346 2604
rect 3970 2564 3976 2576
rect 1412 2536 3976 2564
rect 1412 2505 1440 2536
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 15194 2564 15200 2576
rect 6886 2536 15200 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 1397 2459 1455 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 6886 2496 6914 2536
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 19337 2567 19395 2573
rect 19337 2533 19349 2567
rect 19383 2564 19395 2567
rect 20254 2564 20260 2576
rect 19383 2536 20260 2564
rect 19383 2533 19395 2536
rect 19337 2527 19395 2533
rect 20254 2524 20260 2536
rect 20312 2524 20318 2576
rect 26145 2567 26203 2573
rect 22066 2536 23980 2564
rect 5307 2468 6914 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 15841 2499 15899 2505
rect 7064 2468 7109 2496
rect 7064 2456 7070 2468
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 22066 2496 22094 2536
rect 23842 2496 23848 2508
rect 15887 2468 22094 2496
rect 22940 2468 23848 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19426 2428 19432 2440
rect 19291 2400 19432 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19889 2431 19947 2437
rect 19889 2397 19901 2431
rect 19935 2428 19947 2431
rect 20070 2428 20076 2440
rect 19935 2400 20076 2428
rect 19935 2397 19947 2400
rect 19889 2391 19947 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20680 2400 20729 2428
rect 20680 2388 20686 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 22940 2437 22968 2468
rect 23842 2456 23848 2468
rect 23900 2456 23906 2508
rect 23952 2496 23980 2536
rect 26145 2533 26157 2567
rect 26191 2564 26203 2567
rect 26694 2564 26700 2576
rect 26191 2536 26700 2564
rect 26191 2533 26203 2536
rect 26145 2527 26203 2533
rect 26694 2524 26700 2536
rect 26752 2524 26758 2576
rect 35544 2564 35572 2604
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 36357 2635 36415 2641
rect 36357 2632 36369 2635
rect 35676 2604 36369 2632
rect 35676 2592 35682 2604
rect 36357 2601 36369 2604
rect 36403 2601 36415 2635
rect 39114 2632 39120 2644
rect 39075 2604 39120 2632
rect 36357 2595 36415 2601
rect 39114 2592 39120 2604
rect 39172 2592 39178 2644
rect 41690 2632 41696 2644
rect 41651 2604 41696 2632
rect 41690 2592 41696 2604
rect 41748 2592 41754 2644
rect 42518 2632 42524 2644
rect 42479 2604 42524 2632
rect 42518 2592 42524 2604
rect 42576 2592 42582 2644
rect 42886 2632 42892 2644
rect 42847 2604 42892 2632
rect 42886 2592 42892 2604
rect 42944 2592 42950 2644
rect 38289 2567 38347 2573
rect 38289 2564 38301 2567
rect 35544 2536 38301 2564
rect 38289 2533 38301 2536
rect 38335 2533 38347 2567
rect 38289 2527 38347 2533
rect 41233 2567 41291 2573
rect 41233 2533 41245 2567
rect 41279 2564 41291 2567
rect 43070 2564 43076 2576
rect 41279 2536 43076 2564
rect 41279 2533 41291 2536
rect 41233 2527 41291 2533
rect 43070 2524 43076 2536
rect 43128 2524 43134 2576
rect 27249 2499 27307 2505
rect 23952 2468 27200 2496
rect 22925 2431 22983 2437
rect 21232 2400 22416 2428
rect 21232 2388 21238 2400
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 2774 2360 2780 2372
rect 1627 2332 2780 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7558 2360 7564 2372
rect 6779 2332 7564 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 4172 2292 4200 2323
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8444 2332 9413 2360
rect 8444 2320 8450 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21968 2332 22293 2360
rect 21968 2320 21974 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22388 2360 22416 2400
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 23566 2428 23572 2440
rect 23527 2400 23572 2428
rect 22925 2391 22983 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25556 2400 25697 2428
rect 25556 2388 25562 2400
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26476 2400 26985 2428
rect 26476 2388 26482 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 27172 2428 27200 2468
rect 27249 2465 27261 2499
rect 27295 2496 27307 2499
rect 27982 2496 27988 2508
rect 27295 2468 27988 2496
rect 27295 2465 27307 2468
rect 27249 2459 27307 2465
rect 27982 2456 27988 2468
rect 28040 2456 28046 2508
rect 28092 2468 31064 2496
rect 28092 2428 28120 2468
rect 27172 2400 28120 2428
rect 26973 2391 27031 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 28408 2400 28457 2428
rect 28408 2388 28414 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29696 2400 29929 2428
rect 29696 2388 29702 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 22388 2332 23796 2360
rect 22281 2323 22339 2329
rect 4430 2292 4436 2304
rect 2648 2264 4200 2292
rect 4391 2264 4436 2292
rect 2648 2252 2654 2264
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 7006 2292 7012 2304
rect 6512 2264 7012 2292
rect 6512 2252 6518 2264
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 16850 2292 16856 2304
rect 16811 2264 16856 2292
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 23661 2295 23719 2301
rect 23661 2292 23673 2295
rect 22060 2264 23673 2292
rect 22060 2252 22066 2264
rect 23661 2261 23673 2264
rect 23707 2261 23719 2295
rect 23768 2292 23796 2332
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 28074 2320 28080 2372
rect 28132 2360 28138 2372
rect 31036 2360 31064 2468
rect 31202 2456 31208 2508
rect 31260 2496 31266 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 31260 2468 40509 2496
rect 31260 2456 31266 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 43254 2496 43260 2508
rect 40497 2459 40555 2465
rect 42444 2468 43260 2496
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35492 2400 35725 2428
rect 35492 2388 35498 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 37366 2428 37372 2440
rect 35713 2391 35771 2397
rect 35866 2400 37372 2428
rect 35866 2360 35894 2400
rect 37366 2388 37372 2400
rect 37424 2388 37430 2440
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 38068 2400 38117 2428
rect 38068 2388 38074 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39301 2431 39359 2437
rect 39301 2397 39313 2431
rect 39347 2428 39359 2431
rect 39942 2428 39948 2440
rect 39347 2400 39948 2428
rect 39347 2397 39359 2400
rect 39301 2391 39359 2397
rect 39942 2388 39948 2400
rect 40000 2388 40006 2440
rect 41230 2388 41236 2440
rect 41288 2428 41294 2440
rect 42444 2437 42472 2468
rect 43254 2456 43260 2468
rect 43312 2496 43318 2508
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 43312 2468 46489 2496
rect 43312 2456 43318 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 47394 2456 47400 2508
rect 47452 2496 47458 2508
rect 47857 2499 47915 2505
rect 47857 2496 47869 2499
rect 47452 2468 47869 2496
rect 47452 2456 47458 2468
rect 47857 2465 47869 2468
rect 47903 2465 47915 2499
rect 47857 2459 47915 2465
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 41288 2400 41889 2428
rect 41288 2388 41294 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 42429 2431 42487 2437
rect 42429 2397 42441 2431
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 46201 2431 46259 2437
rect 46201 2397 46213 2431
rect 46247 2428 46259 2431
rect 47026 2428 47032 2440
rect 46247 2400 47032 2428
rect 46247 2397 46259 2400
rect 46201 2391 46259 2397
rect 28132 2332 30788 2360
rect 31036 2332 35894 2360
rect 28132 2320 28138 2332
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 23768 2264 24961 2292
rect 23661 2255 23719 2261
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 29730 2292 29736 2304
rect 29691 2264 29736 2292
rect 24949 2255 25007 2261
rect 29730 2252 29736 2264
rect 29788 2252 29794 2304
rect 30760 2292 30788 2332
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 36136 2332 36277 2360
rect 36136 2320 36142 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 39390 2320 39396 2372
rect 39448 2360 39454 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39448 2332 40325 2360
rect 39448 2320 39454 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 35529 2295 35587 2301
rect 35529 2292 35541 2295
rect 30760 2264 35541 2292
rect 35529 2261 35541 2264
rect 35575 2261 35587 2295
rect 35529 2255 35587 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 43916 2292 43944 2391
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 47673 2431 47731 2437
rect 47673 2397 47685 2431
rect 47719 2428 47731 2431
rect 48038 2428 48044 2440
rect 47719 2400 48044 2428
rect 47719 2397 47731 2400
rect 47673 2391 47731 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 45373 2363 45431 2369
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 45462 2292 45468 2304
rect 38712 2264 43944 2292
rect 45423 2264 45468 2292
rect 38712 2252 38718 2264
rect 45462 2252 45468 2264
rect 45520 2252 45526 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 23934 2088 23940 2100
rect 9732 2060 23940 2088
rect 9732 2048 9738 2060
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 4430 1980 4436 2032
rect 4488 2020 4494 2032
rect 29546 2020 29552 2032
rect 4488 1992 29552 2020
rect 4488 1980 4494 1992
rect 29546 1980 29552 1992
rect 29604 1980 29610 2032
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 3568 1924 6914 1952
rect 3568 1912 3574 1924
rect 6886 1884 6914 1924
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 26786 1952 26792 1964
rect 16908 1924 26792 1952
rect 16908 1912 16914 1924
rect 26786 1912 26792 1924
rect 26844 1912 26850 1964
rect 28718 1912 28724 1964
rect 28776 1952 28782 1964
rect 45462 1952 45468 1964
rect 28776 1924 45468 1952
rect 28776 1912 28782 1924
rect 45462 1912 45468 1924
rect 45520 1912 45526 1964
rect 28442 1884 28448 1896
rect 6886 1856 28448 1884
rect 28442 1844 28448 1856
rect 28500 1844 28506 1896
rect 29730 1844 29736 1896
rect 29788 1884 29794 1896
rect 42518 1884 42524 1896
rect 29788 1856 42524 1884
rect 29788 1844 29794 1856
rect 42518 1844 42524 1856
rect 42576 1844 42582 1896
<< via1 >>
rect 45560 47880 45612 47932
rect 46112 47880 46164 47932
rect 40040 47404 40092 47456
rect 41236 47404 41288 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 21916 47200 21968 47252
rect 36912 47200 36964 47252
rect 46848 47200 46900 47252
rect 20536 47132 20588 47184
rect 28908 47132 28960 47184
rect 35348 47132 35400 47184
rect 44456 47132 44508 47184
rect 47768 47132 47820 47184
rect 30748 47107 30800 47116
rect 1952 46996 2004 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5816 46996 5868 47048
rect 7380 47039 7432 47048
rect 7380 47005 7389 47039
rect 7389 47005 7423 47039
rect 7423 47005 7432 47039
rect 7380 46996 7432 47005
rect 9036 46996 9088 47048
rect 11612 47039 11664 47048
rect 11612 47005 11621 47039
rect 11621 47005 11655 47039
rect 11655 47005 11664 47039
rect 11612 46996 11664 47005
rect 12256 46996 12308 47048
rect 12900 46996 12952 47048
rect 13820 46996 13872 47048
rect 14372 47039 14424 47048
rect 14372 47005 14381 47039
rect 14381 47005 14415 47039
rect 14415 47005 14424 47039
rect 14372 46996 14424 47005
rect 16488 46996 16540 47048
rect 17776 46996 17828 47048
rect 20996 47039 21048 47048
rect 20996 47005 21005 47039
rect 21005 47005 21039 47039
rect 21039 47005 21048 47039
rect 20996 46996 21048 47005
rect 2504 46928 2556 46980
rect 4068 46971 4120 46980
rect 2596 46860 2648 46912
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 7472 46928 7524 46980
rect 9496 46928 9548 46980
rect 11704 46928 11756 46980
rect 12440 46928 12492 46980
rect 2872 46903 2924 46912
rect 2872 46869 2881 46903
rect 2881 46869 2915 46903
rect 2915 46869 2924 46903
rect 4896 46903 4948 46912
rect 2872 46860 2924 46869
rect 4896 46869 4905 46903
rect 4905 46869 4939 46903
rect 4939 46869 4948 46903
rect 4896 46860 4948 46869
rect 18696 46860 18748 46912
rect 20628 46928 20680 46980
rect 19984 46860 20036 46912
rect 24584 46996 24636 47048
rect 25412 47039 25464 47048
rect 25412 47005 25421 47039
rect 25421 47005 25455 47039
rect 25455 47005 25464 47039
rect 25412 46996 25464 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 29368 46928 29420 46980
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 39304 47064 39356 47116
rect 48320 47064 48372 47116
rect 34704 46996 34756 47048
rect 38108 46996 38160 47048
rect 41880 47039 41932 47048
rect 41880 47005 41889 47039
rect 41889 47005 41923 47039
rect 41923 47005 41932 47039
rect 41880 46996 41932 47005
rect 43812 46996 43864 47048
rect 44456 46996 44508 47048
rect 47676 46996 47728 47048
rect 37372 46928 37424 46980
rect 39304 46928 39356 46980
rect 43076 46928 43128 46980
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 3884 46588 3936 46640
rect 24584 46563 24636 46572
rect 24584 46529 24593 46563
rect 24593 46529 24627 46563
rect 24627 46529 24636 46563
rect 24584 46520 24636 46529
rect 12072 46452 12124 46504
rect 13544 46452 13596 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 19248 46495 19300 46504
rect 14280 46452 14332 46461
rect 19248 46461 19257 46495
rect 19257 46461 19291 46495
rect 19291 46461 19300 46495
rect 19248 46452 19300 46461
rect 20444 46495 20496 46504
rect 18604 46384 18656 46436
rect 20444 46461 20453 46495
rect 20453 46461 20487 46495
rect 20487 46461 20496 46495
rect 20444 46452 20496 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 32220 46384 32272 46436
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47952 46563 48004 46572
rect 47952 46529 47961 46563
rect 47961 46529 47995 46563
rect 47995 46529 48004 46563
rect 47952 46520 48004 46529
rect 34428 46495 34480 46504
rect 34428 46461 34437 46495
rect 34437 46461 34471 46495
rect 34471 46461 34480 46495
rect 34428 46452 34480 46461
rect 34796 46452 34848 46504
rect 38292 46495 38344 46504
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 45192 46495 45244 46504
rect 42524 46384 42576 46436
rect 45192 46461 45201 46495
rect 45201 46461 45235 46495
rect 45235 46461 45244 46495
rect 45192 46452 45244 46461
rect 46756 46495 46808 46504
rect 46756 46461 46765 46495
rect 46765 46461 46799 46495
rect 46799 46461 46808 46495
rect 46756 46452 46808 46461
rect 46664 46384 46716 46436
rect 2320 46316 2372 46368
rect 2412 46316 2464 46368
rect 10968 46316 11020 46368
rect 38660 46316 38712 46368
rect 39948 46316 40000 46368
rect 41236 46359 41288 46368
rect 41236 46325 41245 46359
rect 41245 46325 41279 46359
rect 41279 46325 41288 46359
rect 41236 46316 41288 46325
rect 47308 46316 47360 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 12072 46155 12124 46164
rect 12072 46121 12081 46155
rect 12081 46121 12115 46155
rect 12115 46121 12124 46155
rect 12072 46112 12124 46121
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 18604 46155 18656 46164
rect 18604 46121 18613 46155
rect 18613 46121 18647 46155
rect 18647 46121 18656 46155
rect 18604 46112 18656 46121
rect 19248 46112 19300 46164
rect 24768 46112 24820 46164
rect 32312 46112 32364 46164
rect 34428 46112 34480 46164
rect 34796 46155 34848 46164
rect 34796 46121 34805 46155
rect 34805 46121 34839 46155
rect 34839 46121 34848 46155
rect 34796 46112 34848 46121
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 45192 46112 45244 46164
rect 2412 45976 2464 46028
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 20996 45976 21048 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25412 45976 25464 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 11980 45951 12032 45960
rect 11980 45917 11989 45951
rect 11989 45917 12023 45951
rect 12023 45917 12032 45951
rect 11980 45908 12032 45917
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 14096 45908 14148 45917
rect 18696 45908 18748 45960
rect 24584 45951 24636 45960
rect 24584 45917 24593 45951
rect 24593 45917 24627 45951
rect 24627 45917 24636 45951
rect 24584 45908 24636 45917
rect 32588 45908 32640 45960
rect 35440 45908 35492 45960
rect 41236 46019 41288 46028
rect 41236 45985 41245 46019
rect 41245 45985 41279 46019
rect 41279 45985 41288 46019
rect 41236 45976 41288 45985
rect 41972 46019 42024 46028
rect 41972 45985 41981 46019
rect 41981 45985 42015 46019
rect 42015 45985 42024 46019
rect 41972 45976 42024 45985
rect 45100 46044 45152 46096
rect 45652 46044 45704 46096
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 2228 45840 2280 45892
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 41420 45883 41472 45892
rect 41420 45849 41429 45883
rect 41429 45849 41463 45883
rect 41463 45849 41472 45883
rect 41420 45840 41472 45849
rect 45744 45908 45796 45960
rect 46296 45840 46348 45892
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 26884 45772 26936 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 2228 45611 2280 45620
rect 2228 45577 2237 45611
rect 2237 45577 2271 45611
rect 2271 45577 2280 45611
rect 2228 45568 2280 45577
rect 11980 45568 12032 45620
rect 20904 45611 20956 45620
rect 1952 45432 2004 45484
rect 20904 45577 20913 45611
rect 20913 45577 20947 45611
rect 20947 45577 20956 45611
rect 20904 45568 20956 45577
rect 24584 45568 24636 45620
rect 36176 45568 36228 45620
rect 42616 45568 42668 45620
rect 45560 45568 45612 45620
rect 25412 45543 25464 45552
rect 25412 45509 25421 45543
rect 25421 45509 25455 45543
rect 25455 45509 25464 45543
rect 25412 45500 25464 45509
rect 41420 45500 41472 45552
rect 25780 45432 25832 45484
rect 41052 45475 41104 45484
rect 41052 45441 41061 45475
rect 41061 45441 41095 45475
rect 41095 45441 41104 45475
rect 41052 45432 41104 45441
rect 32588 45364 32640 45416
rect 24584 45296 24636 45348
rect 41880 45432 41932 45484
rect 42892 45407 42944 45416
rect 42892 45373 42901 45407
rect 42901 45373 42935 45407
rect 42935 45373 42944 45407
rect 42892 45364 42944 45373
rect 44088 45407 44140 45416
rect 44088 45373 44097 45407
rect 44097 45373 44131 45407
rect 44131 45373 44140 45407
rect 44088 45364 44140 45373
rect 44916 45364 44968 45416
rect 45192 45407 45244 45416
rect 45192 45373 45201 45407
rect 45201 45373 45235 45407
rect 45235 45373 45244 45407
rect 45192 45364 45244 45373
rect 45744 45407 45796 45416
rect 45744 45373 45753 45407
rect 45753 45373 45787 45407
rect 45787 45373 45796 45407
rect 45744 45364 45796 45373
rect 46848 45296 46900 45348
rect 48044 45271 48096 45280
rect 48044 45237 48053 45271
rect 48053 45237 48087 45271
rect 48087 45237 48096 45271
rect 48044 45228 48096 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 42892 45067 42944 45076
rect 42892 45033 42901 45067
rect 42901 45033 42935 45067
rect 42935 45033 42944 45067
rect 42892 45024 42944 45033
rect 44456 45067 44508 45076
rect 44456 45033 44465 45067
rect 44465 45033 44499 45067
rect 44499 45033 44508 45067
rect 44456 45024 44508 45033
rect 45192 45024 45244 45076
rect 45376 45024 45428 45076
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 45560 44820 45612 44872
rect 45744 44820 45796 44872
rect 47676 44752 47728 44804
rect 47860 44684 47912 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 46480 44480 46532 44532
rect 46664 44480 46716 44532
rect 44916 44387 44968 44396
rect 44916 44353 44925 44387
rect 44925 44353 44959 44387
rect 44959 44353 44968 44387
rect 44916 44344 44968 44353
rect 46296 44387 46348 44396
rect 46296 44353 46305 44387
rect 46305 44353 46339 44387
rect 46339 44353 46348 44387
rect 46296 44344 46348 44353
rect 47492 44344 47544 44396
rect 47400 44276 47452 44328
rect 41052 44208 41104 44260
rect 47584 44208 47636 44260
rect 46480 44140 46532 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 46480 43843 46532 43852
rect 46480 43809 46489 43843
rect 46489 43809 46523 43843
rect 46523 43809 46532 43843
rect 46480 43800 46532 43809
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 47676 43435 47728 43444
rect 47676 43401 47685 43435
rect 47685 43401 47719 43435
rect 47719 43401 47728 43435
rect 47676 43392 47728 43401
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 47400 43256 47452 43308
rect 1492 43188 1544 43240
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 46296 42168 46348 42220
rect 47860 42168 47912 42220
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46480 41216 46532 41268
rect 14096 41080 14148 41132
rect 46848 41080 46900 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 39212 40876 39264 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 26976 40536 27028 40588
rect 26608 40468 26660 40520
rect 47032 40511 47084 40520
rect 47032 40477 47041 40511
rect 47041 40477 47075 40511
rect 47075 40477 47084 40511
rect 47032 40468 47084 40477
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 2044 40443 2096 40452
rect 2044 40409 2053 40443
rect 2053 40409 2087 40443
rect 2087 40409 2096 40443
rect 2044 40400 2096 40409
rect 26240 40375 26292 40384
rect 26240 40341 26249 40375
rect 26249 40341 26283 40375
rect 26283 40341 26292 40375
rect 26240 40332 26292 40341
rect 26884 40332 26936 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 26424 40128 26476 40180
rect 23480 40060 23532 40112
rect 19248 39992 19300 40044
rect 47584 40035 47636 40044
rect 47584 40001 47593 40035
rect 47593 40001 47627 40035
rect 47627 40001 47636 40035
rect 47584 39992 47636 40001
rect 23848 39924 23900 39976
rect 25136 39924 25188 39976
rect 19984 39831 20036 39840
rect 19984 39797 19993 39831
rect 19993 39797 20027 39831
rect 20027 39797 20036 39831
rect 19984 39788 20036 39797
rect 46480 39788 46532 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 23480 39584 23532 39636
rect 25136 39627 25188 39636
rect 25136 39593 25145 39627
rect 25145 39593 25179 39627
rect 25179 39593 25188 39627
rect 25136 39584 25188 39593
rect 26056 39584 26108 39636
rect 26608 39627 26660 39636
rect 26240 39516 26292 39568
rect 26608 39593 26617 39627
rect 26617 39593 26651 39627
rect 26651 39593 26660 39627
rect 26608 39584 26660 39593
rect 47032 39516 47084 39568
rect 18144 39380 18196 39432
rect 22100 39380 22152 39432
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 26424 39380 26476 39432
rect 18972 39312 19024 39364
rect 19984 39312 20036 39364
rect 20996 39287 21048 39296
rect 20996 39253 21005 39287
rect 21005 39253 21039 39287
rect 21039 39253 21048 39287
rect 20996 39244 21048 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 18972 39083 19024 39092
rect 18972 39049 18981 39083
rect 18981 39049 19015 39083
rect 19015 39049 19024 39083
rect 18972 39040 19024 39049
rect 20996 39040 21048 39092
rect 25136 38972 25188 39024
rect 21824 38904 21876 38956
rect 23480 38904 23532 38956
rect 29920 38947 29972 38956
rect 20076 38879 20128 38888
rect 20076 38845 20085 38879
rect 20085 38845 20119 38879
rect 20119 38845 20128 38879
rect 20076 38836 20128 38845
rect 20168 38879 20220 38888
rect 20168 38845 20177 38879
rect 20177 38845 20211 38879
rect 20211 38845 20220 38879
rect 20168 38836 20220 38845
rect 22008 38836 22060 38888
rect 23848 38879 23900 38888
rect 23848 38845 23857 38879
rect 23857 38845 23891 38879
rect 23891 38845 23900 38879
rect 23848 38836 23900 38845
rect 24124 38879 24176 38888
rect 24124 38845 24133 38879
rect 24133 38845 24167 38879
rect 24167 38845 24176 38879
rect 24124 38836 24176 38845
rect 24768 38836 24820 38888
rect 29920 38913 29929 38947
rect 29929 38913 29963 38947
rect 29963 38913 29972 38947
rect 29920 38904 29972 38913
rect 45560 38904 45612 38956
rect 47860 38947 47912 38956
rect 47860 38913 47869 38947
rect 47869 38913 47903 38947
rect 47903 38913 47912 38947
rect 47860 38904 47912 38913
rect 27252 38879 27304 38888
rect 19248 38700 19300 38752
rect 22100 38743 22152 38752
rect 22100 38709 22109 38743
rect 22109 38709 22143 38743
rect 22143 38709 22152 38743
rect 23296 38743 23348 38752
rect 22100 38700 22152 38709
rect 23296 38709 23305 38743
rect 23305 38709 23339 38743
rect 23339 38709 23348 38743
rect 23296 38700 23348 38709
rect 25320 38700 25372 38752
rect 27252 38845 27261 38879
rect 27261 38845 27295 38879
rect 27295 38845 27304 38879
rect 27252 38836 27304 38845
rect 27344 38836 27396 38888
rect 30012 38879 30064 38888
rect 30012 38845 30021 38879
rect 30021 38845 30055 38879
rect 30055 38845 30064 38879
rect 30012 38836 30064 38845
rect 30104 38879 30156 38888
rect 30104 38845 30113 38879
rect 30113 38845 30147 38879
rect 30147 38845 30156 38879
rect 30104 38836 30156 38845
rect 29828 38768 29880 38820
rect 29000 38700 29052 38752
rect 46388 38700 46440 38752
rect 46572 38700 46624 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 20076 38496 20128 38548
rect 24124 38496 24176 38548
rect 25136 38539 25188 38548
rect 25136 38505 25145 38539
rect 25145 38505 25179 38539
rect 25179 38505 25188 38539
rect 25136 38496 25188 38505
rect 25320 38496 25372 38548
rect 29920 38496 29972 38548
rect 20444 38360 20496 38412
rect 23480 38360 23532 38412
rect 24768 38360 24820 38412
rect 18512 38292 18564 38344
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 20536 38335 20588 38344
rect 20536 38301 20545 38335
rect 20545 38301 20579 38335
rect 20579 38301 20588 38335
rect 20536 38292 20588 38301
rect 21180 38292 21232 38344
rect 22008 38335 22060 38344
rect 22008 38301 22017 38335
rect 22017 38301 22051 38335
rect 22051 38301 22060 38335
rect 22008 38292 22060 38301
rect 24952 38292 25004 38344
rect 26516 38360 26568 38412
rect 27528 38403 27580 38412
rect 26424 38292 26476 38344
rect 27528 38369 27537 38403
rect 27537 38369 27571 38403
rect 27571 38369 27580 38403
rect 27528 38360 27580 38369
rect 29828 38360 29880 38412
rect 46388 38403 46440 38412
rect 46388 38369 46397 38403
rect 46397 38369 46431 38403
rect 46431 38369 46440 38403
rect 46388 38360 46440 38369
rect 48044 38403 48096 38412
rect 48044 38369 48053 38403
rect 48053 38369 48087 38403
rect 48087 38369 48096 38403
rect 48044 38360 48096 38369
rect 27344 38292 27396 38344
rect 29000 38335 29052 38344
rect 29000 38301 29009 38335
rect 29009 38301 29043 38335
rect 29043 38301 29052 38335
rect 29000 38292 29052 38301
rect 46112 38292 46164 38344
rect 22376 38224 22428 38276
rect 23296 38224 23348 38276
rect 25964 38267 26016 38276
rect 25964 38233 25973 38267
rect 25973 38233 26007 38267
rect 26007 38233 26016 38267
rect 25964 38224 26016 38233
rect 19340 38199 19392 38208
rect 19340 38165 19349 38199
rect 19349 38165 19383 38199
rect 19383 38165 19392 38199
rect 19340 38156 19392 38165
rect 20536 38156 20588 38208
rect 23756 38199 23808 38208
rect 23756 38165 23765 38199
rect 23765 38165 23799 38199
rect 23799 38165 23808 38199
rect 23756 38156 23808 38165
rect 26424 38199 26476 38208
rect 26424 38165 26433 38199
rect 26433 38165 26467 38199
rect 26467 38165 26476 38199
rect 26424 38156 26476 38165
rect 27160 38156 27212 38208
rect 27344 38199 27396 38208
rect 27344 38165 27353 38199
rect 27353 38165 27387 38199
rect 27387 38165 27396 38199
rect 27344 38156 27396 38165
rect 31116 38224 31168 38276
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 11704 37952 11756 38004
rect 22192 37952 22244 38004
rect 22376 37995 22428 38004
rect 22376 37961 22385 37995
rect 22385 37961 22419 37995
rect 22419 37961 22428 37995
rect 22376 37952 22428 37961
rect 24952 37995 25004 38004
rect 24952 37961 24961 37995
rect 24961 37961 24995 37995
rect 24995 37961 25004 37995
rect 24952 37952 25004 37961
rect 27252 37952 27304 38004
rect 30012 37952 30064 38004
rect 31116 37995 31168 38004
rect 31116 37961 31125 37995
rect 31125 37961 31159 37995
rect 31159 37961 31168 37995
rect 31116 37952 31168 37961
rect 17500 37748 17552 37800
rect 18144 37884 18196 37936
rect 19340 37884 19392 37936
rect 21824 37884 21876 37936
rect 20996 37816 21048 37868
rect 22560 37859 22612 37868
rect 22560 37825 22569 37859
rect 22569 37825 22603 37859
rect 22603 37825 22612 37859
rect 22560 37816 22612 37825
rect 18236 37748 18288 37800
rect 19432 37748 19484 37800
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 25412 37791 25464 37800
rect 25412 37757 25421 37791
rect 25421 37757 25455 37791
rect 25455 37757 25464 37791
rect 25412 37748 25464 37757
rect 25780 37884 25832 37936
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 27528 37748 27580 37800
rect 20168 37680 20220 37732
rect 20536 37723 20588 37732
rect 20536 37689 20545 37723
rect 20545 37689 20579 37723
rect 20579 37689 20588 37723
rect 20536 37680 20588 37689
rect 22192 37680 22244 37732
rect 30932 37816 30984 37868
rect 33232 37816 33284 37868
rect 46296 37816 46348 37868
rect 30012 37748 30064 37800
rect 34704 37748 34756 37800
rect 19340 37655 19392 37664
rect 19340 37621 19349 37655
rect 19349 37621 19383 37655
rect 19383 37621 19392 37655
rect 19340 37612 19392 37621
rect 23480 37612 23532 37664
rect 23664 37612 23716 37664
rect 27896 37612 27948 37664
rect 30104 37612 30156 37664
rect 32680 37612 32732 37664
rect 46480 37612 46532 37664
rect 47768 37655 47820 37664
rect 47768 37621 47777 37655
rect 47777 37621 47811 37655
rect 47811 37621 47820 37655
rect 47768 37612 47820 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 18236 37451 18288 37460
rect 18236 37417 18245 37451
rect 18245 37417 18279 37451
rect 18279 37417 18288 37451
rect 18236 37408 18288 37417
rect 22560 37408 22612 37460
rect 27344 37451 27396 37460
rect 27344 37417 27353 37451
rect 27353 37417 27387 37451
rect 27387 37417 27396 37451
rect 27344 37408 27396 37417
rect 30012 37451 30064 37460
rect 30012 37417 30021 37451
rect 30021 37417 30055 37451
rect 30055 37417 30064 37451
rect 30012 37408 30064 37417
rect 20076 37272 20128 37324
rect 23664 37315 23716 37324
rect 23664 37281 23673 37315
rect 23673 37281 23707 37315
rect 23707 37281 23716 37315
rect 23664 37272 23716 37281
rect 1768 37204 1820 37256
rect 19340 37204 19392 37256
rect 23756 37204 23808 37256
rect 24676 37247 24728 37256
rect 24676 37213 24685 37247
rect 24685 37213 24719 37247
rect 24719 37213 24728 37247
rect 24676 37204 24728 37213
rect 25136 37204 25188 37256
rect 27344 37272 27396 37324
rect 26516 37247 26568 37256
rect 26516 37213 26525 37247
rect 26525 37213 26559 37247
rect 26559 37213 26568 37247
rect 26516 37204 26568 37213
rect 29644 37315 29696 37324
rect 25596 37136 25648 37188
rect 29644 37281 29653 37315
rect 29653 37281 29687 37315
rect 29687 37281 29696 37315
rect 29644 37272 29696 37281
rect 29920 37272 29972 37324
rect 32680 37315 32732 37324
rect 32680 37281 32689 37315
rect 32689 37281 32723 37315
rect 32723 37281 32732 37315
rect 32680 37272 32732 37281
rect 34704 37272 34756 37324
rect 35256 37315 35308 37324
rect 35256 37281 35265 37315
rect 35265 37281 35299 37315
rect 35299 37281 35308 37315
rect 35256 37272 35308 37281
rect 46480 37315 46532 37324
rect 46480 37281 46489 37315
rect 46489 37281 46523 37315
rect 46523 37281 46532 37315
rect 46480 37272 46532 37281
rect 48136 37315 48188 37324
rect 48136 37281 48145 37315
rect 48145 37281 48179 37315
rect 48179 37281 48188 37315
rect 48136 37272 48188 37281
rect 29828 37204 29880 37256
rect 35348 37204 35400 37256
rect 33692 37136 33744 37188
rect 47768 37136 47820 37188
rect 19984 37068 20036 37120
rect 23572 37111 23624 37120
rect 23572 37077 23581 37111
rect 23581 37077 23615 37111
rect 23615 37077 23624 37111
rect 24768 37111 24820 37120
rect 23572 37068 23624 37077
rect 24768 37077 24777 37111
rect 24777 37077 24811 37111
rect 24811 37077 24820 37111
rect 24768 37068 24820 37077
rect 28172 37068 28224 37120
rect 33968 37068 34020 37120
rect 34704 37111 34756 37120
rect 34704 37077 34713 37111
rect 34713 37077 34747 37111
rect 34747 37077 34756 37111
rect 34704 37068 34756 37077
rect 35164 37111 35216 37120
rect 35164 37077 35173 37111
rect 35173 37077 35207 37111
rect 35207 37077 35216 37111
rect 35164 37068 35216 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 19984 36864 20036 36916
rect 23572 36864 23624 36916
rect 24768 36864 24820 36916
rect 23756 36796 23808 36848
rect 24860 36796 24912 36848
rect 25136 36839 25188 36848
rect 25136 36805 25145 36839
rect 25145 36805 25179 36839
rect 25179 36805 25188 36839
rect 25136 36796 25188 36805
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 19248 36771 19300 36780
rect 19248 36737 19257 36771
rect 19257 36737 19291 36771
rect 19291 36737 19300 36771
rect 19248 36728 19300 36737
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 20260 36771 20312 36780
rect 20260 36737 20269 36771
rect 20269 36737 20303 36771
rect 20303 36737 20312 36771
rect 20260 36728 20312 36737
rect 22100 36771 22152 36780
rect 22100 36737 22109 36771
rect 22109 36737 22143 36771
rect 22143 36737 22152 36771
rect 22100 36728 22152 36737
rect 23940 36728 23992 36780
rect 25044 36728 25096 36780
rect 25320 36728 25372 36780
rect 26516 36864 26568 36916
rect 30104 36864 30156 36916
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 20444 36660 20496 36712
rect 25596 36660 25648 36712
rect 25964 36728 26016 36780
rect 26240 36771 26292 36780
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 26240 36728 26292 36737
rect 27344 36771 27396 36780
rect 27344 36737 27353 36771
rect 27353 36737 27387 36771
rect 27387 36737 27396 36771
rect 27344 36728 27396 36737
rect 30380 36796 30432 36848
rect 31116 36796 31168 36848
rect 29644 36728 29696 36780
rect 26516 36660 26568 36712
rect 26608 36660 26660 36712
rect 29828 36703 29880 36712
rect 29828 36669 29837 36703
rect 29837 36669 29871 36703
rect 29871 36669 29880 36703
rect 29828 36660 29880 36669
rect 30104 36703 30156 36712
rect 30104 36669 30113 36703
rect 30113 36669 30147 36703
rect 30147 36669 30156 36703
rect 30104 36660 30156 36669
rect 30196 36660 30248 36712
rect 33232 36864 33284 36916
rect 34704 36864 34756 36916
rect 35164 36864 35216 36916
rect 33968 36728 34020 36780
rect 34612 36703 34664 36712
rect 34612 36669 34621 36703
rect 34621 36669 34655 36703
rect 34655 36669 34664 36703
rect 34612 36660 34664 36669
rect 12440 36592 12492 36644
rect 26792 36592 26844 36644
rect 22192 36567 22244 36576
rect 22192 36533 22201 36567
rect 22201 36533 22235 36567
rect 22235 36533 22244 36567
rect 22192 36524 22244 36533
rect 24860 36524 24912 36576
rect 25964 36524 26016 36576
rect 26148 36524 26200 36576
rect 30840 36524 30892 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 2044 36252 2096 36304
rect 19248 36252 19300 36304
rect 19616 36252 19668 36304
rect 19984 36252 20036 36304
rect 19524 36227 19576 36236
rect 19524 36193 19533 36227
rect 19533 36193 19567 36227
rect 19567 36193 19576 36227
rect 19524 36184 19576 36193
rect 20996 36184 21048 36236
rect 22468 36184 22520 36236
rect 24676 36320 24728 36372
rect 25412 36320 25464 36372
rect 25044 36252 25096 36304
rect 26240 36320 26292 36372
rect 29092 36320 29144 36372
rect 29644 36320 29696 36372
rect 30104 36320 30156 36372
rect 31116 36320 31168 36372
rect 33692 36320 33744 36372
rect 26148 36295 26200 36304
rect 26148 36261 26157 36295
rect 26157 36261 26191 36295
rect 26191 36261 26200 36295
rect 26148 36252 26200 36261
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 19340 36159 19392 36168
rect 19340 36125 19349 36159
rect 19349 36125 19383 36159
rect 19383 36125 19392 36159
rect 19340 36116 19392 36125
rect 21180 36159 21232 36168
rect 20352 36048 20404 36100
rect 21180 36125 21189 36159
rect 21189 36125 21223 36159
rect 21223 36125 21232 36159
rect 21180 36116 21232 36125
rect 24860 36159 24912 36168
rect 18512 35980 18564 36032
rect 21088 35980 21140 36032
rect 22192 36048 22244 36100
rect 24860 36125 24869 36159
rect 24869 36125 24903 36159
rect 24903 36125 24912 36159
rect 24860 36116 24912 36125
rect 25044 36048 25096 36100
rect 22376 35980 22428 36032
rect 26516 36048 26568 36100
rect 26792 36091 26844 36100
rect 26792 36057 26801 36091
rect 26801 36057 26835 36091
rect 26835 36057 26844 36091
rect 26792 36048 26844 36057
rect 28080 36048 28132 36100
rect 29000 36159 29052 36168
rect 29000 36125 29009 36159
rect 29009 36125 29043 36159
rect 29043 36125 29052 36159
rect 29000 36116 29052 36125
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 30196 36184 30248 36236
rect 30472 36116 30524 36168
rect 30932 36159 30984 36168
rect 30932 36125 30941 36159
rect 30941 36125 30975 36159
rect 30975 36125 30984 36159
rect 30932 36116 30984 36125
rect 32312 36116 32364 36168
rect 31300 36048 31352 36100
rect 27068 35980 27120 36032
rect 30196 35980 30248 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 17500 35776 17552 35828
rect 21180 35776 21232 35828
rect 21364 35776 21416 35828
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 17960 35683 18012 35692
rect 17960 35649 17969 35683
rect 17969 35649 18003 35683
rect 18003 35649 18012 35683
rect 17960 35640 18012 35649
rect 21088 35708 21140 35760
rect 19340 35683 19392 35692
rect 19340 35649 19349 35683
rect 19349 35649 19383 35683
rect 19383 35649 19392 35683
rect 19340 35640 19392 35649
rect 19432 35683 19484 35692
rect 19432 35649 19441 35683
rect 19441 35649 19475 35683
rect 19475 35649 19484 35683
rect 19432 35640 19484 35649
rect 20352 35683 20404 35692
rect 20352 35649 20361 35683
rect 20361 35649 20395 35683
rect 20395 35649 20404 35683
rect 20352 35640 20404 35649
rect 16672 35504 16724 35556
rect 1860 35436 1912 35488
rect 16948 35436 17000 35488
rect 20444 35572 20496 35624
rect 19984 35504 20036 35556
rect 19248 35436 19300 35488
rect 20996 35504 21048 35556
rect 22468 35776 22520 35828
rect 30380 35776 30432 35828
rect 31300 35819 31352 35828
rect 31300 35785 31309 35819
rect 31309 35785 31343 35819
rect 31343 35785 31352 35819
rect 31300 35776 31352 35785
rect 29000 35708 29052 35760
rect 29920 35708 29972 35760
rect 30196 35708 30248 35760
rect 22376 35683 22428 35692
rect 22376 35649 22385 35683
rect 22385 35649 22419 35683
rect 22419 35649 22428 35683
rect 22376 35640 22428 35649
rect 30288 35683 30340 35692
rect 30288 35649 30297 35683
rect 30297 35649 30331 35683
rect 30331 35649 30340 35683
rect 30288 35640 30340 35649
rect 48136 35683 48188 35692
rect 48136 35649 48145 35683
rect 48145 35649 48179 35683
rect 48179 35649 48188 35683
rect 48136 35640 48188 35649
rect 22192 35615 22244 35624
rect 22192 35581 22201 35615
rect 22201 35581 22235 35615
rect 22235 35581 22244 35615
rect 22192 35572 22244 35581
rect 28080 35572 28132 35624
rect 29184 35572 29236 35624
rect 30472 35572 30524 35624
rect 29000 35504 29052 35556
rect 29920 35504 29972 35556
rect 20536 35479 20588 35488
rect 20536 35445 20545 35479
rect 20545 35445 20579 35479
rect 20579 35445 20588 35479
rect 20536 35436 20588 35445
rect 30840 35436 30892 35488
rect 47124 35436 47176 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 20444 35232 20496 35284
rect 21180 35232 21232 35284
rect 22008 35232 22060 35284
rect 29000 35275 29052 35284
rect 29000 35241 29009 35275
rect 29009 35241 29043 35275
rect 29043 35241 29052 35275
rect 29000 35232 29052 35241
rect 34612 35232 34664 35284
rect 17960 35164 18012 35216
rect 16672 35071 16724 35080
rect 16672 35037 16681 35071
rect 16681 35037 16715 35071
rect 16715 35037 16724 35071
rect 16672 35028 16724 35037
rect 16948 35071 17000 35080
rect 16948 35037 16957 35071
rect 16957 35037 16991 35071
rect 16991 35037 17000 35071
rect 16948 35028 17000 35037
rect 19340 35139 19392 35148
rect 19340 35105 19349 35139
rect 19349 35105 19383 35139
rect 19383 35105 19392 35139
rect 19340 35096 19392 35105
rect 20352 35096 20404 35148
rect 22192 35096 22244 35148
rect 17592 35071 17644 35080
rect 17592 35037 17601 35071
rect 17601 35037 17635 35071
rect 17635 35037 17644 35071
rect 17592 35028 17644 35037
rect 17776 35071 17828 35080
rect 17776 35037 17785 35071
rect 17785 35037 17819 35071
rect 17819 35037 17828 35071
rect 17776 35028 17828 35037
rect 18236 35028 18288 35080
rect 19248 35028 19300 35080
rect 20536 35028 20588 35080
rect 23480 35028 23532 35080
rect 24124 35028 24176 35080
rect 19156 34960 19208 35012
rect 22928 34960 22980 35012
rect 27988 35003 28040 35012
rect 27988 34969 27997 35003
rect 27997 34969 28031 35003
rect 28031 34969 28040 35003
rect 27988 34960 28040 34969
rect 28632 35003 28684 35012
rect 28632 34969 28641 35003
rect 28641 34969 28675 35003
rect 28675 34969 28684 35003
rect 28632 34960 28684 34969
rect 29276 35096 29328 35148
rect 29828 35096 29880 35148
rect 33968 35139 34020 35148
rect 33968 35105 33977 35139
rect 33977 35105 34011 35139
rect 34011 35105 34020 35139
rect 33968 35096 34020 35105
rect 35348 35139 35400 35148
rect 35348 35105 35357 35139
rect 35357 35105 35391 35139
rect 35391 35105 35400 35139
rect 35348 35096 35400 35105
rect 35808 35096 35860 35148
rect 29184 35028 29236 35080
rect 30012 35071 30064 35080
rect 30012 35037 30021 35071
rect 30021 35037 30055 35071
rect 30055 35037 30064 35071
rect 30012 35028 30064 35037
rect 29736 34960 29788 35012
rect 30104 34960 30156 35012
rect 18052 34892 18104 34944
rect 21456 34892 21508 34944
rect 23572 34892 23624 34944
rect 30472 35028 30524 35080
rect 31208 35028 31260 35080
rect 32588 34960 32640 35012
rect 34796 35028 34848 35080
rect 47032 35028 47084 35080
rect 47860 35028 47912 35080
rect 48044 35028 48096 35080
rect 34060 34960 34112 35012
rect 33508 34935 33560 34944
rect 33508 34901 33517 34935
rect 33517 34901 33551 34935
rect 33551 34901 33560 34935
rect 33508 34892 33560 34901
rect 34520 34892 34572 34944
rect 35624 34892 35676 34944
rect 47860 34892 47912 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 17592 34688 17644 34740
rect 18052 34620 18104 34672
rect 18512 34620 18564 34672
rect 19340 34688 19392 34740
rect 25504 34688 25556 34740
rect 30012 34688 30064 34740
rect 32588 34731 32640 34740
rect 17500 34595 17552 34604
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 20168 34527 20220 34536
rect 20168 34493 20177 34527
rect 20177 34493 20211 34527
rect 20211 34493 20220 34527
rect 20168 34484 20220 34493
rect 22192 34620 22244 34672
rect 23572 34620 23624 34672
rect 24124 34620 24176 34672
rect 20444 34595 20496 34604
rect 20444 34561 20453 34595
rect 20453 34561 20487 34595
rect 20487 34561 20496 34595
rect 20444 34552 20496 34561
rect 22008 34552 22060 34604
rect 24768 34595 24820 34604
rect 24768 34561 24777 34595
rect 24777 34561 24811 34595
rect 24811 34561 24820 34595
rect 24768 34552 24820 34561
rect 25044 34595 25096 34604
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 26424 34620 26476 34672
rect 25044 34552 25096 34561
rect 22836 34527 22888 34536
rect 22836 34493 22845 34527
rect 22845 34493 22879 34527
rect 22879 34493 22888 34527
rect 22836 34484 22888 34493
rect 22560 34416 22612 34468
rect 19156 34348 19208 34400
rect 21272 34348 21324 34400
rect 25228 34484 25280 34536
rect 27252 34552 27304 34604
rect 29184 34620 29236 34672
rect 32588 34697 32597 34731
rect 32597 34697 32631 34731
rect 32631 34697 32640 34731
rect 32588 34688 32640 34697
rect 34612 34688 34664 34740
rect 35624 34731 35676 34740
rect 28356 34552 28408 34604
rect 29736 34595 29788 34604
rect 29736 34561 29745 34595
rect 29745 34561 29779 34595
rect 29779 34561 29788 34595
rect 29736 34552 29788 34561
rect 31116 34552 31168 34604
rect 31576 34595 31628 34604
rect 31576 34561 31585 34595
rect 31585 34561 31619 34595
rect 31619 34561 31628 34595
rect 35624 34697 35633 34731
rect 35633 34697 35667 34731
rect 35667 34697 35676 34731
rect 35624 34688 35676 34697
rect 32496 34595 32548 34604
rect 31576 34552 31628 34561
rect 32496 34561 32505 34595
rect 32505 34561 32539 34595
rect 32539 34561 32548 34595
rect 32496 34552 32548 34561
rect 34060 34595 34112 34604
rect 34060 34561 34069 34595
rect 34069 34561 34103 34595
rect 34103 34561 34112 34595
rect 34060 34552 34112 34561
rect 34612 34552 34664 34604
rect 34796 34552 34848 34604
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 35532 34552 35584 34561
rect 47768 34595 47820 34604
rect 47768 34561 47777 34595
rect 47777 34561 47811 34595
rect 47811 34561 47820 34595
rect 47768 34552 47820 34561
rect 24216 34416 24268 34468
rect 26424 34484 26476 34536
rect 29276 34527 29328 34536
rect 29276 34493 29285 34527
rect 29285 34493 29319 34527
rect 29319 34493 29328 34527
rect 29276 34484 29328 34493
rect 29920 34484 29972 34536
rect 27436 34416 27488 34468
rect 24308 34391 24360 34400
rect 24308 34357 24317 34391
rect 24317 34357 24351 34391
rect 24351 34357 24360 34391
rect 24308 34348 24360 34357
rect 24952 34391 25004 34400
rect 24952 34357 24961 34391
rect 24961 34357 24995 34391
rect 24995 34357 25004 34391
rect 27344 34391 27396 34400
rect 24952 34348 25004 34357
rect 27344 34357 27353 34391
rect 27353 34357 27387 34391
rect 27387 34357 27396 34391
rect 27344 34348 27396 34357
rect 33508 34416 33560 34468
rect 30748 34391 30800 34400
rect 30748 34357 30757 34391
rect 30757 34357 30791 34391
rect 30791 34357 30800 34391
rect 30748 34348 30800 34357
rect 33968 34391 34020 34400
rect 33968 34357 33977 34391
rect 33977 34357 34011 34391
rect 34011 34357 34020 34391
rect 33968 34348 34020 34357
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 20168 34144 20220 34196
rect 20812 34144 20864 34196
rect 21364 34187 21416 34196
rect 21364 34153 21373 34187
rect 21373 34153 21407 34187
rect 21407 34153 21416 34187
rect 21364 34144 21416 34153
rect 22836 34144 22888 34196
rect 24768 34144 24820 34196
rect 27160 34144 27212 34196
rect 27436 34144 27488 34196
rect 35532 34144 35584 34196
rect 9496 34076 9548 34128
rect 20444 34051 20496 34060
rect 20444 34017 20453 34051
rect 20453 34017 20487 34051
rect 20487 34017 20496 34051
rect 20444 34008 20496 34017
rect 29276 34076 29328 34128
rect 27712 34008 27764 34060
rect 28908 34008 28960 34060
rect 30748 34008 30800 34060
rect 32864 34008 32916 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 47584 34051 47636 34060
rect 47584 34017 47593 34051
rect 47593 34017 47627 34051
rect 47627 34017 47636 34051
rect 47584 34008 47636 34017
rect 1584 33983 1636 33992
rect 1584 33949 1593 33983
rect 1593 33949 1627 33983
rect 1627 33949 1636 33983
rect 1584 33940 1636 33949
rect 20352 33940 20404 33992
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 21456 33983 21508 33992
rect 21456 33949 21465 33983
rect 21465 33949 21499 33983
rect 21499 33949 21508 33983
rect 21456 33940 21508 33949
rect 22744 33983 22796 33992
rect 22744 33949 22753 33983
rect 22753 33949 22787 33983
rect 22787 33949 22796 33983
rect 22744 33940 22796 33949
rect 22836 33940 22888 33992
rect 23296 33983 23348 33992
rect 20904 33872 20956 33924
rect 23296 33949 23305 33983
rect 23305 33949 23339 33983
rect 23339 33949 23348 33983
rect 23296 33940 23348 33949
rect 23756 33872 23808 33924
rect 24308 33872 24360 33924
rect 1952 33804 2004 33856
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 25412 33915 25464 33924
rect 25412 33881 25421 33915
rect 25421 33881 25455 33915
rect 25455 33881 25464 33915
rect 25412 33872 25464 33881
rect 26424 33872 26476 33924
rect 27252 33872 27304 33924
rect 27436 33872 27488 33924
rect 29184 33940 29236 33992
rect 29736 33940 29788 33992
rect 30012 33940 30064 33992
rect 30104 33983 30156 33992
rect 30104 33949 30113 33983
rect 30113 33949 30147 33983
rect 30147 33949 30156 33983
rect 30104 33940 30156 33949
rect 30288 33983 30340 33992
rect 30288 33949 30297 33983
rect 30297 33949 30331 33983
rect 30331 33949 30340 33983
rect 30288 33940 30340 33949
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 31116 33872 31168 33924
rect 20720 33804 20772 33813
rect 26332 33804 26384 33856
rect 29552 33804 29604 33856
rect 31300 33804 31352 33856
rect 32772 33847 32824 33856
rect 32772 33813 32781 33847
rect 32781 33813 32815 33847
rect 32815 33813 32824 33847
rect 32772 33804 32824 33813
rect 34520 33940 34572 33992
rect 34612 33940 34664 33992
rect 34796 33940 34848 33992
rect 35164 33940 35216 33992
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 19064 33600 19116 33652
rect 20720 33600 20772 33652
rect 22744 33600 22796 33652
rect 23756 33600 23808 33652
rect 23848 33600 23900 33652
rect 24216 33600 24268 33652
rect 23572 33532 23624 33584
rect 14372 33464 14424 33516
rect 20996 33464 21048 33516
rect 23664 33507 23716 33516
rect 23664 33473 23673 33507
rect 23673 33473 23707 33507
rect 23707 33473 23716 33507
rect 23664 33464 23716 33473
rect 27344 33532 27396 33584
rect 29184 33600 29236 33652
rect 30012 33643 30064 33652
rect 30012 33609 30021 33643
rect 30021 33609 30055 33643
rect 30055 33609 30064 33643
rect 30012 33600 30064 33609
rect 35164 33643 35216 33652
rect 35164 33609 35173 33643
rect 35173 33609 35207 33643
rect 35207 33609 35216 33643
rect 35164 33600 35216 33609
rect 47768 33600 47820 33652
rect 28908 33532 28960 33584
rect 29092 33532 29144 33584
rect 29276 33532 29328 33584
rect 31024 33532 31076 33584
rect 23848 33464 23900 33516
rect 24124 33464 24176 33516
rect 24676 33507 24728 33516
rect 24676 33473 24685 33507
rect 24685 33473 24719 33507
rect 24719 33473 24728 33507
rect 24676 33464 24728 33473
rect 27436 33507 27488 33516
rect 27436 33473 27445 33507
rect 27445 33473 27479 33507
rect 27479 33473 27488 33507
rect 27436 33464 27488 33473
rect 29460 33507 29512 33516
rect 29460 33473 29469 33507
rect 29469 33473 29503 33507
rect 29503 33473 29512 33507
rect 29460 33464 29512 33473
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 1676 33439 1728 33448
rect 1676 33405 1685 33439
rect 1685 33405 1719 33439
rect 1719 33405 1728 33439
rect 1676 33396 1728 33405
rect 21088 33396 21140 33448
rect 26976 33396 27028 33448
rect 27712 33396 27764 33448
rect 28448 33396 28500 33448
rect 28724 33396 28776 33448
rect 29920 33396 29972 33448
rect 32772 33532 32824 33584
rect 32496 33464 32548 33516
rect 33048 33464 33100 33516
rect 34796 33464 34848 33516
rect 46756 33507 46808 33516
rect 46756 33473 46765 33507
rect 46765 33473 46799 33507
rect 46799 33473 46808 33507
rect 46756 33464 46808 33473
rect 47492 33464 47544 33516
rect 20812 33328 20864 33380
rect 19800 33260 19852 33312
rect 22928 33303 22980 33312
rect 22928 33269 22937 33303
rect 22937 33269 22971 33303
rect 22971 33269 22980 33303
rect 22928 33260 22980 33269
rect 23572 33260 23624 33312
rect 26240 33260 26292 33312
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 31576 33328 31628 33380
rect 29552 33303 29604 33312
rect 27160 33260 27212 33269
rect 29552 33269 29561 33303
rect 29561 33269 29595 33303
rect 29595 33269 29604 33303
rect 29552 33260 29604 33269
rect 29644 33260 29696 33312
rect 32404 33303 32456 33312
rect 32404 33269 32413 33303
rect 32413 33269 32447 33303
rect 32447 33269 32456 33303
rect 32404 33260 32456 33269
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1952 33099 2004 33108
rect 1952 33065 1961 33099
rect 1961 33065 1995 33099
rect 1995 33065 2004 33099
rect 1952 33056 2004 33065
rect 20996 33099 21048 33108
rect 20996 33065 21005 33099
rect 21005 33065 21039 33099
rect 21039 33065 21048 33099
rect 20996 33056 21048 33065
rect 23848 33056 23900 33108
rect 25412 33056 25464 33108
rect 20904 32988 20956 33040
rect 1676 32852 1728 32904
rect 1952 32852 2004 32904
rect 18236 32920 18288 32972
rect 19800 32963 19852 32972
rect 2228 32716 2280 32768
rect 18144 32716 18196 32768
rect 19800 32929 19809 32963
rect 19809 32929 19843 32963
rect 19843 32929 19852 32963
rect 19800 32920 19852 32929
rect 20076 32920 20128 32972
rect 21456 32920 21508 32972
rect 20536 32852 20588 32904
rect 23664 32895 23716 32904
rect 23664 32861 23673 32895
rect 23673 32861 23707 32895
rect 23707 32861 23716 32895
rect 23664 32852 23716 32861
rect 24308 32988 24360 33040
rect 27252 33056 27304 33108
rect 27528 33056 27580 33108
rect 29184 33056 29236 33108
rect 31116 33056 31168 33108
rect 34796 33099 34848 33108
rect 34796 33065 34805 33099
rect 34805 33065 34839 33099
rect 34839 33065 34848 33099
rect 34796 33056 34848 33065
rect 27344 32988 27396 33040
rect 29644 32988 29696 33040
rect 25320 32920 25372 32972
rect 25964 32920 26016 32972
rect 28264 32920 28316 32972
rect 24952 32852 25004 32904
rect 25412 32895 25464 32904
rect 20352 32784 20404 32836
rect 22836 32784 22888 32836
rect 23020 32784 23072 32836
rect 25412 32861 25421 32895
rect 25421 32861 25455 32895
rect 25455 32861 25464 32895
rect 25412 32852 25464 32861
rect 26332 32895 26384 32904
rect 26332 32861 26341 32895
rect 26341 32861 26375 32895
rect 26375 32861 26384 32895
rect 26332 32852 26384 32861
rect 27988 32852 28040 32904
rect 28448 32895 28500 32904
rect 28448 32861 28457 32895
rect 28457 32861 28491 32895
rect 28491 32861 28500 32895
rect 28448 32852 28500 32861
rect 28540 32852 28592 32904
rect 28908 32852 28960 32904
rect 29460 32852 29512 32904
rect 29736 32920 29788 32972
rect 31024 32963 31076 32972
rect 31024 32929 31033 32963
rect 31033 32929 31067 32963
rect 31067 32929 31076 32963
rect 31024 32920 31076 32929
rect 31300 32963 31352 32972
rect 31300 32929 31309 32963
rect 31309 32929 31343 32963
rect 31343 32929 31352 32963
rect 31300 32920 31352 32929
rect 30380 32852 30432 32904
rect 32404 32852 32456 32904
rect 33048 32852 33100 32904
rect 35716 32852 35768 32904
rect 26148 32784 26200 32836
rect 27528 32784 27580 32836
rect 31392 32784 31444 32836
rect 46940 32784 46992 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 23296 32716 23348 32768
rect 25412 32716 25464 32768
rect 25504 32716 25556 32768
rect 29552 32716 29604 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 3792 32512 3844 32564
rect 2228 32487 2280 32496
rect 2228 32453 2237 32487
rect 2237 32453 2271 32487
rect 2271 32453 2280 32487
rect 2228 32444 2280 32453
rect 18144 32487 18196 32496
rect 18144 32453 18153 32487
rect 18153 32453 18187 32487
rect 18187 32453 18196 32487
rect 18144 32444 18196 32453
rect 23664 32512 23716 32564
rect 1860 32376 1912 32428
rect 19248 32376 19300 32428
rect 4620 32308 4672 32360
rect 1400 32172 1452 32224
rect 7472 32172 7524 32224
rect 17684 32172 17736 32224
rect 19156 32308 19208 32360
rect 20352 32376 20404 32428
rect 20536 32419 20588 32428
rect 20536 32385 20545 32419
rect 20545 32385 20579 32419
rect 20579 32385 20588 32419
rect 20536 32376 20588 32385
rect 20904 32376 20956 32428
rect 21456 32376 21508 32428
rect 24032 32376 24084 32428
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 24584 32308 24636 32360
rect 25964 32444 26016 32496
rect 28356 32512 28408 32564
rect 28448 32512 28500 32564
rect 28908 32512 28960 32564
rect 29000 32512 29052 32564
rect 32864 32512 32916 32564
rect 46940 32555 46992 32564
rect 46940 32521 46949 32555
rect 46949 32521 46983 32555
rect 46983 32521 46992 32555
rect 46940 32512 46992 32521
rect 29460 32444 29512 32496
rect 26148 32376 26200 32428
rect 26240 32419 26292 32428
rect 26240 32385 26249 32419
rect 26249 32385 26283 32419
rect 26283 32385 26292 32419
rect 27436 32419 27488 32428
rect 26240 32376 26292 32385
rect 27436 32385 27445 32419
rect 27445 32385 27479 32419
rect 27479 32385 27488 32419
rect 27436 32376 27488 32385
rect 28264 32376 28316 32428
rect 29736 32419 29788 32428
rect 29736 32385 29745 32419
rect 29745 32385 29779 32419
rect 29779 32385 29788 32419
rect 29736 32376 29788 32385
rect 30932 32376 30984 32428
rect 31392 32376 31444 32428
rect 46480 32376 46532 32428
rect 47400 32376 47452 32428
rect 47952 32419 48004 32428
rect 47952 32385 47961 32419
rect 47961 32385 47995 32419
rect 47995 32385 48004 32419
rect 47952 32376 48004 32385
rect 29184 32308 29236 32360
rect 29828 32351 29880 32360
rect 29828 32317 29837 32351
rect 29837 32317 29871 32351
rect 29871 32317 29880 32351
rect 29828 32308 29880 32317
rect 29920 32351 29972 32360
rect 29920 32317 29929 32351
rect 29929 32317 29963 32351
rect 29963 32317 29972 32351
rect 29920 32308 29972 32317
rect 18880 32172 18932 32224
rect 20076 32215 20128 32224
rect 20076 32181 20085 32215
rect 20085 32181 20119 32215
rect 20119 32181 20128 32215
rect 20076 32172 20128 32181
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 24216 32172 24268 32224
rect 25780 32240 25832 32292
rect 25504 32215 25556 32224
rect 25504 32181 25513 32215
rect 25513 32181 25547 32215
rect 25547 32181 25556 32215
rect 25504 32172 25556 32181
rect 25596 32172 25648 32224
rect 28540 32215 28592 32224
rect 28540 32181 28549 32215
rect 28549 32181 28583 32215
rect 28583 32181 28592 32215
rect 28540 32172 28592 32181
rect 29184 32172 29236 32224
rect 30748 32172 30800 32224
rect 31484 32172 31536 32224
rect 32036 32172 32088 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3884 31968 3936 32020
rect 1952 31900 2004 31952
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 3792 31875 3844 31884
rect 3792 31841 3801 31875
rect 3801 31841 3835 31875
rect 3835 31841 3844 31875
rect 3792 31832 3844 31841
rect 8300 31900 8352 31952
rect 4620 31875 4672 31884
rect 4620 31841 4629 31875
rect 4629 31841 4663 31875
rect 4663 31841 4672 31875
rect 4620 31832 4672 31841
rect 5448 31832 5500 31884
rect 15200 31832 15252 31884
rect 19248 31968 19300 32020
rect 20076 31968 20128 32020
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 17684 31832 17736 31884
rect 17776 31807 17828 31816
rect 17776 31773 17785 31807
rect 17785 31773 17819 31807
rect 17819 31773 17828 31807
rect 17776 31764 17828 31773
rect 19156 31832 19208 31884
rect 18236 31764 18288 31816
rect 19432 31832 19484 31884
rect 24124 31968 24176 32020
rect 26976 31968 27028 32020
rect 29736 31968 29788 32020
rect 41696 31968 41748 32020
rect 47584 31968 47636 32020
rect 24584 31900 24636 31952
rect 24768 31900 24820 31952
rect 27896 31900 27948 31952
rect 29920 31900 29972 31952
rect 32496 31943 32548 31952
rect 32496 31909 32505 31943
rect 32505 31909 32539 31943
rect 32539 31909 32548 31943
rect 32496 31900 32548 31909
rect 20720 31764 20772 31816
rect 20996 31764 21048 31816
rect 22928 31832 22980 31884
rect 25412 31832 25464 31884
rect 25596 31832 25648 31884
rect 28264 31832 28316 31884
rect 22008 31807 22060 31816
rect 22008 31773 22017 31807
rect 22017 31773 22051 31807
rect 22051 31773 22060 31807
rect 22008 31764 22060 31773
rect 24032 31807 24084 31816
rect 24032 31773 24041 31807
rect 24041 31773 24075 31807
rect 24075 31773 24084 31807
rect 24032 31764 24084 31773
rect 24216 31807 24268 31816
rect 24216 31773 24225 31807
rect 24225 31773 24259 31807
rect 24259 31773 24268 31807
rect 24216 31764 24268 31773
rect 25780 31764 25832 31816
rect 26976 31764 27028 31816
rect 27436 31764 27488 31816
rect 27712 31764 27764 31816
rect 31392 31832 31444 31884
rect 29092 31764 29144 31816
rect 30104 31807 30156 31816
rect 30104 31773 30113 31807
rect 30113 31773 30147 31807
rect 30147 31773 30156 31807
rect 30104 31764 30156 31773
rect 31484 31764 31536 31816
rect 32864 31832 32916 31884
rect 45836 31764 45888 31816
rect 47492 31900 47544 31952
rect 46756 31875 46808 31884
rect 46756 31841 46765 31875
rect 46765 31841 46799 31875
rect 46799 31841 46808 31875
rect 46756 31832 46808 31841
rect 47584 31875 47636 31884
rect 47584 31841 47593 31875
rect 47593 31841 47627 31875
rect 47627 31841 47636 31875
rect 47584 31832 47636 31841
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 12900 31696 12952 31748
rect 15016 31739 15068 31748
rect 15016 31705 15025 31739
rect 15025 31705 15059 31739
rect 15059 31705 15068 31739
rect 15016 31696 15068 31705
rect 22284 31739 22336 31748
rect 22284 31705 22293 31739
rect 22293 31705 22327 31739
rect 22327 31705 22336 31739
rect 22284 31696 22336 31705
rect 23572 31696 23624 31748
rect 30380 31739 30432 31748
rect 30380 31705 30389 31739
rect 30389 31705 30423 31739
rect 30423 31705 30432 31739
rect 30380 31696 30432 31705
rect 34796 31696 34848 31748
rect 18328 31671 18380 31680
rect 18328 31637 18337 31671
rect 18337 31637 18371 31671
rect 18371 31637 18380 31671
rect 18328 31628 18380 31637
rect 25136 31671 25188 31680
rect 25136 31637 25145 31671
rect 25145 31637 25179 31671
rect 25179 31637 25188 31671
rect 25136 31628 25188 31637
rect 25596 31671 25648 31680
rect 25596 31637 25605 31671
rect 25605 31637 25639 31671
rect 25639 31637 25648 31671
rect 25596 31628 25648 31637
rect 28908 31628 28960 31680
rect 34704 31671 34756 31680
rect 34704 31637 34713 31671
rect 34713 31637 34747 31671
rect 34747 31637 34756 31671
rect 34704 31628 34756 31637
rect 35348 31628 35400 31680
rect 36820 31628 36872 31680
rect 43076 31628 43128 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 12900 31467 12952 31476
rect 12900 31433 12909 31467
rect 12909 31433 12943 31467
rect 12943 31433 12952 31467
rect 12900 31424 12952 31433
rect 15016 31424 15068 31476
rect 19156 31424 19208 31476
rect 22284 31424 22336 31476
rect 2044 31288 2096 31340
rect 14740 31331 14792 31340
rect 14740 31297 14749 31331
rect 14749 31297 14783 31331
rect 14783 31297 14792 31331
rect 14740 31288 14792 31297
rect 19432 31288 19484 31340
rect 25136 31424 25188 31476
rect 27988 31424 28040 31476
rect 24124 31356 24176 31408
rect 29828 31424 29880 31476
rect 30380 31424 30432 31476
rect 31392 31424 31444 31476
rect 24584 31288 24636 31340
rect 25412 31288 25464 31340
rect 26976 31288 27028 31340
rect 27620 31288 27672 31340
rect 28724 31288 28776 31340
rect 29736 31331 29788 31340
rect 29736 31297 29745 31331
rect 29745 31297 29779 31331
rect 29779 31297 29788 31331
rect 29736 31288 29788 31297
rect 30748 31331 30800 31340
rect 30748 31297 30757 31331
rect 30757 31297 30791 31331
rect 30791 31297 30800 31331
rect 30748 31288 30800 31297
rect 32220 31288 32272 31340
rect 36820 31424 36872 31476
rect 35716 31331 35768 31340
rect 35716 31297 35725 31331
rect 35725 31297 35759 31331
rect 35759 31297 35768 31331
rect 35716 31288 35768 31297
rect 18328 31220 18380 31272
rect 24768 31220 24820 31272
rect 25596 31220 25648 31272
rect 29644 31220 29696 31272
rect 32036 31220 32088 31272
rect 25504 31152 25556 31204
rect 18972 31084 19024 31136
rect 28080 31152 28132 31204
rect 31760 31152 31812 31204
rect 32404 31220 32456 31272
rect 33876 31220 33928 31272
rect 25964 31084 26016 31136
rect 30656 31084 30708 31136
rect 35348 31084 35400 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 23572 30880 23624 30932
rect 26976 30923 27028 30932
rect 26976 30889 26985 30923
rect 26985 30889 27019 30923
rect 27019 30889 27028 30923
rect 26976 30880 27028 30889
rect 29644 30923 29696 30932
rect 29644 30889 29653 30923
rect 29653 30889 29687 30923
rect 29687 30889 29696 30923
rect 29644 30880 29696 30889
rect 33048 30880 33100 30932
rect 33876 30923 33928 30932
rect 33876 30889 33885 30923
rect 33885 30889 33919 30923
rect 33919 30889 33928 30923
rect 33876 30880 33928 30889
rect 34796 30880 34848 30932
rect 17868 30787 17920 30796
rect 17868 30753 17877 30787
rect 17877 30753 17911 30787
rect 17911 30753 17920 30787
rect 17868 30744 17920 30753
rect 12532 30719 12584 30728
rect 12532 30685 12541 30719
rect 12541 30685 12575 30719
rect 12575 30685 12584 30719
rect 12532 30676 12584 30685
rect 13452 30676 13504 30728
rect 14188 30676 14240 30728
rect 16304 30719 16356 30728
rect 16304 30685 16313 30719
rect 16313 30685 16347 30719
rect 16347 30685 16356 30719
rect 16304 30676 16356 30685
rect 20168 30676 20220 30728
rect 15016 30651 15068 30660
rect 15016 30617 15025 30651
rect 15025 30617 15059 30651
rect 15059 30617 15068 30651
rect 15016 30608 15068 30617
rect 16580 30608 16632 30660
rect 19432 30608 19484 30660
rect 24308 30676 24360 30728
rect 26792 30744 26844 30796
rect 27068 30744 27120 30796
rect 25964 30719 26016 30728
rect 25964 30685 25971 30719
rect 25971 30685 26016 30719
rect 25964 30676 26016 30685
rect 26148 30719 26200 30728
rect 26148 30685 26157 30719
rect 26157 30685 26191 30719
rect 26191 30685 26200 30719
rect 26148 30676 26200 30685
rect 28080 30744 28132 30796
rect 29184 30744 29236 30796
rect 25228 30608 25280 30660
rect 25688 30608 25740 30660
rect 27528 30676 27580 30728
rect 28356 30719 28408 30728
rect 28356 30685 28365 30719
rect 28365 30685 28399 30719
rect 28399 30685 28408 30719
rect 28356 30676 28408 30685
rect 29552 30719 29604 30728
rect 29552 30685 29561 30719
rect 29561 30685 29595 30719
rect 29595 30685 29604 30719
rect 29552 30676 29604 30685
rect 32036 30744 32088 30796
rect 35808 30744 35860 30796
rect 31484 30719 31536 30728
rect 31484 30685 31493 30719
rect 31493 30685 31527 30719
rect 31527 30685 31536 30719
rect 31484 30676 31536 30685
rect 34704 30676 34756 30728
rect 39304 30676 39356 30728
rect 27896 30608 27948 30660
rect 28448 30608 28500 30660
rect 29000 30608 29052 30660
rect 30104 30608 30156 30660
rect 32220 30608 32272 30660
rect 12440 30540 12492 30592
rect 13084 30583 13136 30592
rect 13084 30549 13093 30583
rect 13093 30549 13127 30583
rect 13127 30549 13136 30583
rect 13084 30540 13136 30549
rect 19340 30540 19392 30592
rect 20352 30583 20404 30592
rect 20352 30549 20361 30583
rect 20361 30549 20395 30583
rect 20395 30549 20404 30583
rect 20352 30540 20404 30549
rect 24860 30540 24912 30592
rect 27344 30583 27396 30592
rect 27344 30549 27353 30583
rect 27353 30549 27387 30583
rect 27387 30549 27396 30583
rect 27344 30540 27396 30549
rect 31760 30540 31812 30592
rect 35164 30583 35216 30592
rect 35164 30549 35173 30583
rect 35173 30549 35207 30583
rect 35207 30549 35216 30583
rect 35164 30540 35216 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 14372 30336 14424 30388
rect 16304 30336 16356 30388
rect 12440 30311 12492 30320
rect 12440 30277 12449 30311
rect 12449 30277 12483 30311
rect 12483 30277 12492 30311
rect 12440 30268 12492 30277
rect 13084 30268 13136 30320
rect 14096 30268 14148 30320
rect 14740 30268 14792 30320
rect 9772 30243 9824 30252
rect 9772 30209 9781 30243
rect 9781 30209 9815 30243
rect 9815 30209 9824 30243
rect 9772 30200 9824 30209
rect 9220 30132 9272 30184
rect 14280 30200 14332 30252
rect 19340 30268 19392 30320
rect 20352 30200 20404 30252
rect 24400 30268 24452 30320
rect 26148 30336 26200 30388
rect 26976 30336 27028 30388
rect 27528 30336 27580 30388
rect 27344 30268 27396 30320
rect 27804 30268 27856 30320
rect 28080 30243 28132 30252
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 35164 30336 35216 30388
rect 28448 30268 28500 30320
rect 34520 30243 34572 30252
rect 16672 30175 16724 30184
rect 9680 29996 9732 30048
rect 10324 30039 10376 30048
rect 10324 30005 10333 30039
rect 10333 30005 10367 30039
rect 10367 30005 10376 30039
rect 10324 29996 10376 30005
rect 16672 30141 16681 30175
rect 16681 30141 16715 30175
rect 16715 30141 16724 30175
rect 16672 30132 16724 30141
rect 17500 30132 17552 30184
rect 18972 30175 19024 30184
rect 15476 30064 15528 30116
rect 12624 29996 12676 30048
rect 15384 29996 15436 30048
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 15844 29996 15896 30048
rect 18972 30141 18981 30175
rect 18981 30141 19015 30175
rect 19015 30141 19024 30175
rect 18972 30132 19024 30141
rect 22100 30132 22152 30184
rect 22652 30132 22704 30184
rect 24860 30132 24912 30184
rect 34520 30209 34529 30243
rect 34529 30209 34563 30243
rect 34563 30209 34572 30243
rect 34520 30200 34572 30209
rect 34612 30200 34664 30252
rect 34796 30200 34848 30252
rect 30012 30132 30064 30184
rect 28356 30064 28408 30116
rect 32496 30064 32548 30116
rect 20904 29996 20956 30048
rect 22284 29996 22336 30048
rect 25688 29996 25740 30048
rect 28540 29996 28592 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12072 29792 12124 29844
rect 16672 29792 16724 29844
rect 17500 29835 17552 29844
rect 17500 29801 17509 29835
rect 17509 29801 17543 29835
rect 17543 29801 17552 29835
rect 17500 29792 17552 29801
rect 20168 29792 20220 29844
rect 20812 29792 20864 29844
rect 21824 29792 21876 29844
rect 11888 29724 11940 29776
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9680 29656 9732 29665
rect 11704 29656 11756 29708
rect 9312 29588 9364 29640
rect 12164 29631 12216 29640
rect 12164 29597 12173 29631
rect 12173 29597 12207 29631
rect 12207 29597 12216 29631
rect 12164 29588 12216 29597
rect 15016 29656 15068 29708
rect 15384 29699 15436 29708
rect 15384 29665 15393 29699
rect 15393 29665 15427 29699
rect 15427 29665 15436 29699
rect 15384 29656 15436 29665
rect 20812 29656 20864 29708
rect 21088 29699 21140 29708
rect 21088 29665 21097 29699
rect 21097 29665 21131 29699
rect 21131 29665 21140 29699
rect 21088 29656 21140 29665
rect 21732 29656 21784 29708
rect 14280 29631 14332 29640
rect 10324 29520 10376 29572
rect 11244 29452 11296 29504
rect 12992 29520 13044 29572
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 18420 29588 18472 29640
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 20720 29588 20772 29640
rect 13084 29452 13136 29504
rect 15476 29520 15528 29572
rect 16764 29520 16816 29572
rect 21088 29520 21140 29572
rect 22100 29631 22152 29640
rect 22100 29597 22109 29631
rect 22109 29597 22143 29631
rect 22143 29597 22152 29631
rect 22100 29588 22152 29597
rect 22284 29588 22336 29640
rect 24400 29792 24452 29844
rect 26056 29792 26108 29844
rect 27068 29835 27120 29844
rect 27068 29801 27077 29835
rect 27077 29801 27111 29835
rect 27111 29801 27120 29835
rect 27068 29792 27120 29801
rect 27988 29792 28040 29844
rect 28356 29792 28408 29844
rect 28540 29835 28592 29844
rect 28540 29801 28549 29835
rect 28549 29801 28583 29835
rect 28583 29801 28592 29835
rect 28540 29792 28592 29801
rect 29920 29792 29972 29844
rect 30932 29835 30984 29844
rect 30932 29801 30941 29835
rect 30941 29801 30975 29835
rect 30975 29801 30984 29835
rect 30932 29792 30984 29801
rect 26516 29724 26568 29776
rect 26884 29724 26936 29776
rect 46848 29792 46900 29844
rect 24308 29588 24360 29640
rect 26148 29588 26200 29640
rect 26329 29631 26381 29640
rect 26329 29597 26338 29631
rect 26338 29597 26372 29631
rect 26372 29597 26381 29631
rect 26329 29588 26381 29597
rect 27804 29656 27856 29708
rect 28724 29588 28776 29640
rect 30656 29656 30708 29708
rect 32864 29656 32916 29708
rect 29736 29631 29788 29640
rect 29736 29597 29743 29631
rect 29743 29597 29788 29631
rect 29736 29588 29788 29597
rect 30012 29631 30064 29640
rect 30012 29597 30026 29631
rect 30026 29597 30060 29631
rect 30060 29597 30064 29631
rect 30012 29588 30064 29597
rect 19340 29452 19392 29504
rect 20720 29452 20772 29504
rect 22008 29452 22060 29504
rect 28264 29520 28316 29572
rect 28448 29563 28500 29572
rect 28448 29529 28457 29563
rect 28457 29529 28491 29563
rect 28491 29529 28500 29563
rect 28448 29520 28500 29529
rect 28540 29520 28592 29572
rect 30196 29588 30248 29640
rect 24400 29452 24452 29504
rect 26240 29452 26292 29504
rect 27528 29452 27580 29504
rect 31484 29588 31536 29640
rect 48136 29631 48188 29640
rect 48136 29597 48145 29631
rect 48145 29597 48179 29631
rect 48179 29597 48188 29631
rect 48136 29588 48188 29597
rect 32864 29520 32916 29572
rect 32772 29452 32824 29504
rect 34060 29452 34112 29504
rect 47400 29452 47452 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 9772 29248 9824 29300
rect 12440 29248 12492 29300
rect 13084 29291 13136 29300
rect 13084 29257 13093 29291
rect 13093 29257 13127 29291
rect 13127 29257 13136 29291
rect 13084 29248 13136 29257
rect 14280 29248 14332 29300
rect 14372 29248 14424 29300
rect 16580 29248 16632 29300
rect 11704 29180 11756 29232
rect 12992 29223 13044 29232
rect 12992 29189 13001 29223
rect 13001 29189 13035 29223
rect 13035 29189 13044 29223
rect 12992 29180 13044 29189
rect 15752 29180 15804 29232
rect 20904 29223 20956 29232
rect 20904 29189 20913 29223
rect 20913 29189 20947 29223
rect 20947 29189 20956 29223
rect 20904 29180 20956 29189
rect 21088 29223 21140 29232
rect 21088 29189 21097 29223
rect 21097 29189 21131 29223
rect 21131 29189 21140 29223
rect 21088 29180 21140 29189
rect 22100 29248 22152 29300
rect 26884 29180 26936 29232
rect 29000 29248 29052 29300
rect 8484 29112 8536 29164
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 12072 29155 12124 29164
rect 12072 29121 12081 29155
rect 12081 29121 12115 29155
rect 12115 29121 12124 29155
rect 12072 29112 12124 29121
rect 9956 29044 10008 29096
rect 12164 29044 12216 29096
rect 16028 29112 16080 29164
rect 19064 29155 19116 29164
rect 19064 29121 19073 29155
rect 19073 29121 19107 29155
rect 19107 29121 19116 29155
rect 19064 29112 19116 29121
rect 22008 29155 22060 29164
rect 22008 29121 22017 29155
rect 22017 29121 22051 29155
rect 22051 29121 22060 29155
rect 22008 29112 22060 29121
rect 22744 29155 22796 29164
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 13360 29044 13412 29096
rect 22284 29087 22336 29096
rect 22284 29053 22293 29087
rect 22293 29053 22327 29087
rect 22327 29053 22336 29087
rect 22284 29044 22336 29053
rect 22376 29044 22428 29096
rect 26976 29112 27028 29164
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27804 29155 27856 29164
rect 27804 29121 27813 29155
rect 27813 29121 27847 29155
rect 27847 29121 27856 29155
rect 27804 29112 27856 29121
rect 27988 29112 28040 29164
rect 28724 29112 28776 29164
rect 29184 29112 29236 29164
rect 32404 29248 32456 29300
rect 32864 29248 32916 29300
rect 34520 29248 34572 29300
rect 29920 29180 29972 29232
rect 31024 29180 31076 29232
rect 32956 29112 33008 29164
rect 34060 29155 34112 29164
rect 34060 29121 34069 29155
rect 34069 29121 34103 29155
rect 34103 29121 34112 29155
rect 34060 29112 34112 29121
rect 28540 29044 28592 29096
rect 30012 29044 30064 29096
rect 32496 29044 32548 29096
rect 33968 29044 34020 29096
rect 35348 29044 35400 29096
rect 11244 28976 11296 29028
rect 17960 28976 18012 29028
rect 18696 28976 18748 29028
rect 26148 28976 26200 29028
rect 26424 28976 26476 29028
rect 28724 28976 28776 29028
rect 21272 28951 21324 28960
rect 21272 28917 21281 28951
rect 21281 28917 21315 28951
rect 21315 28917 21324 28951
rect 21272 28908 21324 28917
rect 22836 28908 22888 28960
rect 26240 28908 26292 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 12624 28704 12676 28756
rect 15476 28704 15528 28756
rect 18328 28704 18380 28756
rect 22744 28704 22796 28756
rect 26332 28704 26384 28756
rect 29736 28704 29788 28756
rect 31024 28704 31076 28756
rect 34060 28704 34112 28756
rect 34796 28704 34848 28756
rect 3792 28636 3844 28688
rect 3976 28568 4028 28620
rect 16396 28568 16448 28620
rect 22284 28636 22336 28688
rect 23112 28636 23164 28688
rect 18696 28611 18748 28620
rect 18696 28577 18705 28611
rect 18705 28577 18739 28611
rect 18739 28577 18748 28611
rect 18696 28568 18748 28577
rect 21088 28568 21140 28620
rect 14188 28500 14240 28552
rect 18512 28500 18564 28552
rect 19340 28500 19392 28552
rect 20904 28500 20956 28552
rect 21548 28543 21600 28552
rect 21548 28509 21557 28543
rect 21557 28509 21591 28543
rect 21591 28509 21600 28543
rect 21548 28500 21600 28509
rect 26424 28568 26476 28620
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 22928 28500 22980 28552
rect 23296 28500 23348 28552
rect 23572 28500 23624 28552
rect 24308 28500 24360 28552
rect 26332 28500 26384 28552
rect 27252 28500 27304 28552
rect 28080 28568 28132 28620
rect 10048 28432 10100 28484
rect 16120 28475 16172 28484
rect 10416 28364 10468 28416
rect 14648 28407 14700 28416
rect 14648 28373 14657 28407
rect 14657 28373 14691 28407
rect 14691 28373 14700 28407
rect 14648 28364 14700 28373
rect 16120 28441 16129 28475
rect 16129 28441 16163 28475
rect 16163 28441 16172 28475
rect 16120 28432 16172 28441
rect 18236 28432 18288 28484
rect 21272 28432 21324 28484
rect 27620 28432 27672 28484
rect 27804 28432 27856 28484
rect 19248 28364 19300 28416
rect 20536 28364 20588 28416
rect 21180 28407 21232 28416
rect 21180 28373 21189 28407
rect 21189 28373 21223 28407
rect 21223 28373 21232 28407
rect 21180 28364 21232 28373
rect 22928 28364 22980 28416
rect 24492 28407 24544 28416
rect 24492 28373 24501 28407
rect 24501 28373 24535 28407
rect 24535 28373 24544 28407
rect 24492 28364 24544 28373
rect 25320 28364 25372 28416
rect 26516 28364 26568 28416
rect 27068 28364 27120 28416
rect 29184 28636 29236 28688
rect 28908 28611 28960 28620
rect 28908 28577 28917 28611
rect 28917 28577 28951 28611
rect 28951 28577 28960 28611
rect 28908 28568 28960 28577
rect 32404 28611 32456 28620
rect 32404 28577 32413 28611
rect 32413 28577 32447 28611
rect 32447 28577 32456 28611
rect 32404 28568 32456 28577
rect 33876 28568 33928 28620
rect 28540 28432 28592 28484
rect 28356 28364 28408 28416
rect 30012 28500 30064 28552
rect 30932 28500 30984 28552
rect 31760 28543 31812 28552
rect 31760 28509 31769 28543
rect 31769 28509 31803 28543
rect 31803 28509 31812 28543
rect 31760 28500 31812 28509
rect 35348 28500 35400 28552
rect 46940 28500 46992 28552
rect 32588 28432 32640 28484
rect 33140 28432 33192 28484
rect 34704 28475 34756 28484
rect 34704 28441 34713 28475
rect 34713 28441 34747 28475
rect 34747 28441 34756 28475
rect 34704 28432 34756 28441
rect 31852 28407 31904 28416
rect 31852 28373 31861 28407
rect 31861 28373 31895 28407
rect 31895 28373 31904 28407
rect 31852 28364 31904 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 16120 28160 16172 28212
rect 16764 28203 16816 28212
rect 16764 28169 16773 28203
rect 16773 28169 16807 28203
rect 16807 28169 16816 28203
rect 16764 28160 16816 28169
rect 17960 28203 18012 28212
rect 17960 28169 17969 28203
rect 17969 28169 18003 28203
rect 18003 28169 18012 28203
rect 17960 28160 18012 28169
rect 18972 28160 19024 28212
rect 8484 28024 8536 28076
rect 9220 28024 9272 28076
rect 9772 28024 9824 28076
rect 18052 28092 18104 28144
rect 11888 28067 11940 28076
rect 11888 28033 11897 28067
rect 11897 28033 11931 28067
rect 11931 28033 11940 28067
rect 11888 28024 11940 28033
rect 12164 28024 12216 28076
rect 13452 28067 13504 28076
rect 11980 27999 12032 28008
rect 11980 27965 11989 27999
rect 11989 27965 12023 27999
rect 12023 27965 12032 27999
rect 11980 27956 12032 27965
rect 13452 28033 13461 28067
rect 13461 28033 13495 28067
rect 13495 28033 13504 28067
rect 13452 28024 13504 28033
rect 15292 28024 15344 28076
rect 16028 28024 16080 28076
rect 17040 28024 17092 28076
rect 18236 28067 18288 28076
rect 18236 28033 18245 28067
rect 18245 28033 18279 28067
rect 18279 28033 18288 28067
rect 18236 28024 18288 28033
rect 19064 28024 19116 28076
rect 22652 28160 22704 28212
rect 23296 28160 23348 28212
rect 27252 28160 27304 28212
rect 28264 28203 28316 28212
rect 20536 28092 20588 28144
rect 21272 28092 21324 28144
rect 22376 28092 22428 28144
rect 22928 28135 22980 28144
rect 22928 28101 22937 28135
rect 22937 28101 22971 28135
rect 22971 28101 22980 28135
rect 22928 28092 22980 28101
rect 24492 28092 24544 28144
rect 28264 28169 28273 28203
rect 28273 28169 28307 28203
rect 28307 28169 28316 28203
rect 28264 28160 28316 28169
rect 32588 28203 32640 28212
rect 32588 28169 32597 28203
rect 32597 28169 32631 28203
rect 32631 28169 32640 28203
rect 32588 28160 32640 28169
rect 47032 28160 47084 28212
rect 22008 28067 22060 28076
rect 14188 27956 14240 28008
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 19524 27999 19576 28008
rect 19524 27965 19533 27999
rect 19533 27965 19567 27999
rect 19567 27965 19576 27999
rect 19524 27956 19576 27965
rect 18604 27888 18656 27940
rect 8300 27863 8352 27872
rect 8300 27829 8309 27863
rect 8309 27829 8343 27863
rect 8343 27829 8352 27863
rect 8300 27820 8352 27829
rect 9680 27820 9732 27872
rect 12164 27863 12216 27872
rect 12164 27829 12173 27863
rect 12173 27829 12207 27863
rect 12207 27829 12216 27863
rect 12164 27820 12216 27829
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 13544 27863 13596 27872
rect 13544 27829 13553 27863
rect 13553 27829 13587 27863
rect 13587 27829 13596 27863
rect 13544 27820 13596 27829
rect 17316 27820 17368 27872
rect 19064 27820 19116 27872
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 27068 28024 27120 28076
rect 21088 27956 21140 28008
rect 22652 27999 22704 28008
rect 22652 27965 22661 27999
rect 22661 27965 22695 27999
rect 22695 27965 22704 27999
rect 22652 27956 22704 27965
rect 25596 27999 25648 28008
rect 25596 27965 25605 27999
rect 25605 27965 25639 27999
rect 25639 27965 25648 27999
rect 25596 27956 25648 27965
rect 21732 27820 21784 27872
rect 27344 27888 27396 27940
rect 27620 28067 27672 28076
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 27988 28024 28040 28076
rect 28356 28024 28408 28076
rect 32772 28067 32824 28076
rect 28080 27956 28132 28008
rect 32772 28033 32781 28067
rect 32781 28033 32815 28067
rect 32815 28033 32824 28067
rect 32772 28024 32824 28033
rect 47676 28024 47728 28076
rect 28264 27888 28316 27940
rect 28540 27931 28592 27940
rect 28540 27897 28549 27931
rect 28549 27897 28583 27931
rect 28583 27897 28592 27931
rect 28540 27888 28592 27897
rect 29184 27888 29236 27940
rect 25136 27863 25188 27872
rect 25136 27829 25145 27863
rect 25145 27829 25179 27863
rect 25179 27829 25188 27863
rect 25136 27820 25188 27829
rect 28448 27820 28500 27872
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 12164 27616 12216 27668
rect 19524 27616 19576 27668
rect 25596 27659 25648 27668
rect 25596 27625 25605 27659
rect 25605 27625 25639 27659
rect 25639 27625 25648 27659
rect 25596 27616 25648 27625
rect 26332 27591 26384 27600
rect 26332 27557 26341 27591
rect 26341 27557 26375 27591
rect 26375 27557 26384 27591
rect 26332 27548 26384 27557
rect 8300 27480 8352 27532
rect 12716 27480 12768 27532
rect 15200 27480 15252 27532
rect 15844 27480 15896 27532
rect 17960 27480 18012 27532
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 14188 27455 14240 27464
rect 14188 27421 14197 27455
rect 14197 27421 14231 27455
rect 14231 27421 14240 27455
rect 14188 27412 14240 27421
rect 17040 27455 17092 27464
rect 17040 27421 17049 27455
rect 17049 27421 17083 27455
rect 17083 27421 17092 27455
rect 17040 27412 17092 27421
rect 18052 27412 18104 27464
rect 21180 27480 21232 27532
rect 21732 27480 21784 27532
rect 25320 27523 25372 27532
rect 25320 27489 25329 27523
rect 25329 27489 25363 27523
rect 25363 27489 25372 27523
rect 25320 27480 25372 27489
rect 26608 27616 26660 27668
rect 26700 27548 26752 27600
rect 27712 27591 27764 27600
rect 18604 27455 18656 27464
rect 9680 27344 9732 27396
rect 13544 27344 13596 27396
rect 14556 27344 14608 27396
rect 15200 27344 15252 27396
rect 18604 27421 18613 27455
rect 18613 27421 18647 27455
rect 18647 27421 18656 27455
rect 18604 27412 18656 27421
rect 19340 27455 19392 27464
rect 19340 27421 19349 27455
rect 19349 27421 19383 27455
rect 19383 27421 19392 27455
rect 19340 27412 19392 27421
rect 11336 27276 11388 27328
rect 11888 27276 11940 27328
rect 15844 27276 15896 27328
rect 16764 27276 16816 27328
rect 17960 27319 18012 27328
rect 17960 27285 17969 27319
rect 17969 27285 18003 27319
rect 18003 27285 18012 27319
rect 17960 27276 18012 27285
rect 18328 27276 18380 27328
rect 20076 27276 20128 27328
rect 22008 27412 22060 27464
rect 25136 27412 25188 27464
rect 27252 27480 27304 27532
rect 27712 27557 27721 27591
rect 27721 27557 27755 27591
rect 27755 27557 27764 27591
rect 27712 27548 27764 27557
rect 28724 27591 28776 27600
rect 28724 27557 28733 27591
rect 28733 27557 28767 27591
rect 28767 27557 28776 27591
rect 28724 27548 28776 27557
rect 33140 27548 33192 27600
rect 21548 27344 21600 27396
rect 21088 27276 21140 27328
rect 23848 27276 23900 27328
rect 25320 27344 25372 27396
rect 28356 27412 28408 27464
rect 28448 27412 28500 27464
rect 28908 27480 28960 27532
rect 31576 27480 31628 27532
rect 31852 27480 31904 27532
rect 30748 27455 30800 27464
rect 30748 27421 30757 27455
rect 30757 27421 30791 27455
rect 30791 27421 30800 27455
rect 30748 27412 30800 27421
rect 31668 27412 31720 27464
rect 33968 27523 34020 27532
rect 33968 27489 33977 27523
rect 33977 27489 34011 27523
rect 34011 27489 34020 27523
rect 33968 27480 34020 27489
rect 36176 27523 36228 27532
rect 36176 27489 36185 27523
rect 36185 27489 36219 27523
rect 36219 27489 36228 27523
rect 36176 27480 36228 27489
rect 40132 27480 40184 27532
rect 46940 27548 46992 27600
rect 47676 27480 47728 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 33876 27412 33928 27464
rect 35348 27455 35400 27464
rect 35348 27421 35357 27455
rect 35357 27421 35391 27455
rect 35391 27421 35400 27455
rect 35348 27412 35400 27421
rect 34060 27344 34112 27396
rect 34704 27344 34756 27396
rect 40040 27387 40092 27396
rect 40040 27353 40049 27387
rect 40049 27353 40083 27387
rect 40083 27353 40092 27387
rect 40040 27344 40092 27353
rect 27068 27276 27120 27328
rect 28080 27276 28132 27328
rect 31392 27276 31444 27328
rect 36176 27276 36228 27328
rect 47584 27276 47636 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8392 27072 8444 27124
rect 10784 27072 10836 27124
rect 10416 27047 10468 27056
rect 10416 27013 10425 27047
rect 10425 27013 10459 27047
rect 10459 27013 10468 27047
rect 10416 27004 10468 27013
rect 13452 27072 13504 27124
rect 15200 27072 15252 27124
rect 17960 27072 18012 27124
rect 25320 27115 25372 27124
rect 9220 26936 9272 26988
rect 9312 26911 9364 26920
rect 9312 26877 9321 26911
rect 9321 26877 9355 26911
rect 9355 26877 9364 26911
rect 9312 26868 9364 26877
rect 10324 26936 10376 26988
rect 10600 26979 10652 26988
rect 10600 26945 10609 26979
rect 10609 26945 10643 26979
rect 10643 26945 10652 26979
rect 10600 26936 10652 26945
rect 11336 26936 11388 26988
rect 11244 26868 11296 26920
rect 17040 27004 17092 27056
rect 17776 27004 17828 27056
rect 25320 27081 25329 27115
rect 25329 27081 25363 27115
rect 25363 27081 25372 27115
rect 25320 27072 25372 27081
rect 27620 27072 27672 27124
rect 23848 27047 23900 27056
rect 23848 27013 23857 27047
rect 23857 27013 23891 27047
rect 23891 27013 23900 27047
rect 23848 27004 23900 27013
rect 25228 27004 25280 27056
rect 27896 27004 27948 27056
rect 13820 26936 13872 26988
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 11612 26868 11664 26920
rect 15844 26936 15896 26988
rect 16120 26868 16172 26920
rect 18144 26800 18196 26852
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 13820 26732 13872 26784
rect 14648 26732 14700 26784
rect 22652 26936 22704 26988
rect 28264 26936 28316 26988
rect 30932 26936 30984 26988
rect 31024 26936 31076 26988
rect 31208 26979 31260 26988
rect 31208 26945 31249 26979
rect 31249 26945 31260 26979
rect 31208 26936 31260 26945
rect 33968 27072 34020 27124
rect 40040 27072 40092 27124
rect 28356 26868 28408 26920
rect 28816 26868 28868 26920
rect 29092 26868 29144 26920
rect 32496 26936 32548 26988
rect 33876 27004 33928 27056
rect 33968 26979 34020 26988
rect 33968 26945 33977 26979
rect 33977 26945 34011 26979
rect 34011 26945 34020 26979
rect 33968 26936 34020 26945
rect 34244 26936 34296 26988
rect 35532 26936 35584 26988
rect 39856 26979 39908 26988
rect 39856 26945 39865 26979
rect 39865 26945 39899 26979
rect 39899 26945 39908 26979
rect 39856 26936 39908 26945
rect 30380 26775 30432 26784
rect 30380 26741 30389 26775
rect 30389 26741 30423 26775
rect 30423 26741 30432 26775
rect 30380 26732 30432 26741
rect 30932 26775 30984 26784
rect 30932 26741 30941 26775
rect 30941 26741 30975 26775
rect 30975 26741 30984 26775
rect 30932 26732 30984 26741
rect 31392 26732 31444 26784
rect 33324 26732 33376 26784
rect 35348 26775 35400 26784
rect 35348 26741 35357 26775
rect 35357 26741 35391 26775
rect 35391 26741 35400 26775
rect 35348 26732 35400 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 20 26392 72 26444
rect 15476 26528 15528 26580
rect 10324 26503 10376 26512
rect 10324 26469 10333 26503
rect 10333 26469 10367 26503
rect 10367 26469 10376 26503
rect 10324 26460 10376 26469
rect 9312 26392 9364 26444
rect 8484 26324 8536 26376
rect 9128 26324 9180 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 10508 26324 10560 26376
rect 11520 26367 11572 26376
rect 9864 26256 9916 26308
rect 10692 26256 10744 26308
rect 11060 26333 11069 26354
rect 11069 26333 11103 26354
rect 11103 26333 11112 26354
rect 11060 26302 11112 26333
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 15292 26460 15344 26512
rect 22928 26528 22980 26580
rect 24308 26528 24360 26580
rect 25228 26571 25280 26580
rect 15844 26460 15896 26512
rect 15476 26435 15528 26444
rect 15476 26401 15485 26435
rect 15485 26401 15519 26435
rect 15519 26401 15528 26435
rect 15476 26392 15528 26401
rect 11612 26256 11664 26308
rect 15752 26324 15804 26376
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 24400 26367 24452 26376
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 25228 26537 25237 26571
rect 25237 26537 25271 26571
rect 25271 26537 25280 26571
rect 25228 26528 25280 26537
rect 31668 26528 31720 26580
rect 26516 26435 26568 26444
rect 26516 26401 26525 26435
rect 26525 26401 26559 26435
rect 26559 26401 26568 26435
rect 26516 26392 26568 26401
rect 25044 26324 25096 26376
rect 26608 26367 26660 26376
rect 26608 26333 26617 26367
rect 26617 26333 26651 26367
rect 26651 26333 26660 26367
rect 26608 26324 26660 26333
rect 27988 26392 28040 26444
rect 27620 26367 27672 26376
rect 27620 26333 27629 26367
rect 27629 26333 27663 26367
rect 27663 26333 27672 26367
rect 27620 26324 27672 26333
rect 28080 26367 28132 26376
rect 28080 26333 28089 26367
rect 28089 26333 28123 26367
rect 28123 26333 28132 26367
rect 28080 26324 28132 26333
rect 28264 26367 28316 26376
rect 28264 26333 28271 26367
rect 28271 26333 28316 26367
rect 28264 26324 28316 26333
rect 32404 26392 32456 26444
rect 32680 26528 32732 26580
rect 39856 26528 39908 26580
rect 26700 26256 26752 26308
rect 27160 26256 27212 26308
rect 27252 26256 27304 26308
rect 27896 26256 27948 26308
rect 28448 26299 28500 26308
rect 28448 26265 28457 26299
rect 28457 26265 28491 26299
rect 28491 26265 28500 26299
rect 28448 26256 28500 26265
rect 7932 26188 7984 26240
rect 8300 26188 8352 26240
rect 9680 26188 9732 26240
rect 11428 26188 11480 26240
rect 17040 26188 17092 26240
rect 26976 26188 27028 26240
rect 28724 26231 28776 26240
rect 28724 26197 28733 26231
rect 28733 26197 28767 26231
rect 28767 26197 28776 26231
rect 28724 26188 28776 26197
rect 28908 26188 28960 26240
rect 33324 26367 33376 26376
rect 30932 26299 30984 26308
rect 30932 26265 30941 26299
rect 30941 26265 30975 26299
rect 30975 26265 30984 26299
rect 30932 26256 30984 26265
rect 31944 26256 31996 26308
rect 31024 26188 31076 26240
rect 32496 26188 32548 26240
rect 32864 26231 32916 26240
rect 32864 26197 32873 26231
rect 32873 26197 32907 26231
rect 32907 26197 32916 26231
rect 32864 26188 32916 26197
rect 33324 26333 33333 26367
rect 33333 26333 33367 26367
rect 33367 26333 33376 26367
rect 33324 26324 33376 26333
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 47676 26367 47728 26376
rect 47676 26333 47685 26367
rect 47685 26333 47719 26367
rect 47719 26333 47728 26367
rect 47676 26324 47728 26333
rect 33600 26256 33652 26308
rect 33784 26256 33836 26308
rect 34244 26188 34296 26240
rect 45100 26231 45152 26240
rect 45100 26197 45109 26231
rect 45109 26197 45143 26231
rect 45143 26197 45152 26231
rect 45100 26188 45152 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9864 25984 9916 26036
rect 16120 26027 16172 26036
rect 16120 25993 16129 26027
rect 16129 25993 16163 26027
rect 16163 25993 16172 26027
rect 16120 25984 16172 25993
rect 16396 25984 16448 26036
rect 18604 25984 18656 26036
rect 8300 25916 8352 25968
rect 8760 25916 8812 25968
rect 10692 25916 10744 25968
rect 11520 25916 11572 25968
rect 15752 25959 15804 25968
rect 15752 25925 15761 25959
rect 15761 25925 15795 25959
rect 15795 25925 15804 25959
rect 15752 25916 15804 25925
rect 16764 25959 16816 25968
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 11336 25848 11388 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 14648 25891 14700 25900
rect 14648 25857 14657 25891
rect 14657 25857 14691 25891
rect 14691 25857 14700 25891
rect 14648 25848 14700 25857
rect 16764 25925 16773 25959
rect 16773 25925 16807 25959
rect 16807 25925 16816 25959
rect 16764 25916 16816 25925
rect 16672 25848 16724 25900
rect 15384 25780 15436 25832
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17408 25848 17460 25900
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 19248 25848 19300 25900
rect 20996 25848 21048 25900
rect 21548 25848 21600 25900
rect 17500 25780 17552 25832
rect 19984 25823 20036 25832
rect 9680 25755 9732 25764
rect 9680 25721 9689 25755
rect 9689 25721 9723 25755
rect 9723 25721 9732 25755
rect 9680 25712 9732 25721
rect 10784 25712 10836 25764
rect 10508 25644 10560 25696
rect 11612 25644 11664 25696
rect 15016 25644 15068 25696
rect 17040 25712 17092 25764
rect 16396 25644 16448 25696
rect 19616 25712 19668 25764
rect 19984 25789 19993 25823
rect 19993 25789 20027 25823
rect 20027 25789 20036 25823
rect 19984 25780 20036 25789
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22560 25848 22612 25900
rect 22928 25891 22980 25900
rect 22928 25857 22937 25891
rect 22937 25857 22971 25891
rect 22971 25857 22980 25891
rect 22928 25848 22980 25857
rect 23204 25891 23256 25900
rect 23204 25857 23213 25891
rect 23213 25857 23247 25891
rect 23247 25857 23256 25891
rect 25412 25916 25464 25968
rect 26608 25916 26660 25968
rect 23204 25848 23256 25857
rect 26976 25891 27028 25900
rect 26976 25857 26985 25891
rect 26985 25857 27019 25891
rect 27019 25857 27028 25891
rect 26976 25848 27028 25857
rect 27252 25891 27304 25900
rect 27252 25857 27261 25891
rect 27261 25857 27295 25891
rect 27295 25857 27304 25891
rect 27252 25848 27304 25857
rect 28448 25916 28500 25968
rect 27436 25891 27488 25900
rect 28908 25984 28960 26036
rect 29092 25984 29144 26036
rect 31944 25984 31996 26036
rect 34244 26027 34296 26036
rect 34244 25993 34253 26027
rect 34253 25993 34287 26027
rect 34287 25993 34296 26027
rect 34244 25984 34296 25993
rect 28724 25916 28776 25968
rect 30380 25916 30432 25968
rect 32864 25916 32916 25968
rect 33784 25916 33836 25968
rect 35440 25916 35492 25968
rect 45100 25916 45152 25968
rect 27436 25857 27450 25891
rect 27450 25857 27484 25891
rect 27484 25857 27488 25891
rect 27436 25848 27488 25857
rect 31668 25848 31720 25900
rect 32404 25848 32456 25900
rect 34796 25848 34848 25900
rect 35348 25848 35400 25900
rect 17408 25644 17460 25696
rect 19248 25644 19300 25696
rect 19524 25644 19576 25696
rect 24032 25780 24084 25832
rect 45100 25823 45152 25832
rect 26608 25712 26660 25764
rect 45100 25789 45109 25823
rect 45109 25789 45143 25823
rect 45143 25789 45152 25823
rect 45100 25780 45152 25789
rect 46848 25823 46900 25832
rect 46848 25789 46857 25823
rect 46857 25789 46891 25823
rect 46891 25789 46900 25823
rect 46848 25780 46900 25789
rect 27344 25644 27396 25696
rect 35900 25644 35952 25696
rect 47768 25687 47820 25696
rect 47768 25653 47777 25687
rect 47777 25653 47811 25687
rect 47811 25653 47820 25687
rect 47768 25644 47820 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10508 25440 10560 25492
rect 14648 25440 14700 25492
rect 16488 25440 16540 25492
rect 19984 25440 20036 25492
rect 22008 25483 22060 25492
rect 22008 25449 22017 25483
rect 22017 25449 22051 25483
rect 22051 25449 22060 25483
rect 22008 25440 22060 25449
rect 24032 25440 24084 25492
rect 25412 25440 25464 25492
rect 26792 25440 26844 25492
rect 33600 25483 33652 25492
rect 33600 25449 33609 25483
rect 33609 25449 33643 25483
rect 33643 25449 33652 25483
rect 33600 25440 33652 25449
rect 20996 25415 21048 25424
rect 10416 25347 10468 25356
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 10600 25304 10652 25356
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 20996 25381 21005 25415
rect 21005 25381 21039 25415
rect 21039 25381 21048 25415
rect 20996 25372 21048 25381
rect 22560 25372 22612 25424
rect 11244 25304 11296 25356
rect 11428 25347 11480 25356
rect 11428 25313 11437 25347
rect 11437 25313 11471 25347
rect 11471 25313 11480 25347
rect 11428 25304 11480 25313
rect 15016 25347 15068 25356
rect 15016 25313 15025 25347
rect 15025 25313 15059 25347
rect 15059 25313 15068 25347
rect 15016 25304 15068 25313
rect 16672 25304 16724 25356
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 18052 25304 18104 25356
rect 19524 25347 19576 25356
rect 19524 25313 19533 25347
rect 19533 25313 19567 25347
rect 19567 25313 19576 25347
rect 19524 25304 19576 25313
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 12624 25236 12676 25288
rect 16396 25236 16448 25288
rect 17040 25236 17092 25288
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17868 25236 17920 25288
rect 22284 25304 22336 25356
rect 27252 25372 27304 25424
rect 27436 25372 27488 25424
rect 28448 25304 28500 25356
rect 31576 25304 31628 25356
rect 35900 25347 35952 25356
rect 35900 25313 35909 25347
rect 35909 25313 35943 25347
rect 35943 25313 35952 25347
rect 35900 25304 35952 25313
rect 47676 25304 47728 25356
rect 25044 25279 25096 25288
rect 13360 25168 13412 25220
rect 15292 25211 15344 25220
rect 15292 25177 15301 25211
rect 15301 25177 15335 25211
rect 15335 25177 15344 25211
rect 15292 25168 15344 25177
rect 19432 25168 19484 25220
rect 19616 25168 19668 25220
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 29920 25236 29972 25288
rect 33416 25279 33468 25288
rect 33416 25245 33425 25279
rect 33425 25245 33459 25279
rect 33459 25245 33468 25279
rect 33416 25236 33468 25245
rect 34796 25236 34848 25288
rect 22376 25168 22428 25220
rect 22928 25168 22980 25220
rect 32128 25168 32180 25220
rect 45560 25168 45612 25220
rect 46940 25168 46992 25220
rect 48136 25211 48188 25220
rect 48136 25177 48145 25211
rect 48145 25177 48179 25211
rect 48179 25177 48188 25211
rect 48136 25168 48188 25177
rect 2044 25100 2096 25152
rect 10048 25100 10100 25152
rect 10784 25100 10836 25152
rect 12072 25100 12124 25152
rect 12532 25143 12584 25152
rect 12532 25109 12541 25143
rect 12541 25109 12575 25143
rect 12575 25109 12584 25143
rect 12532 25100 12584 25109
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 23204 25100 23256 25152
rect 33600 25100 33652 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 13360 24896 13412 24948
rect 15292 24896 15344 24948
rect 22928 24896 22980 24948
rect 23480 24896 23532 24948
rect 33416 24896 33468 24948
rect 42892 24896 42944 24948
rect 12072 24871 12124 24880
rect 12072 24837 12081 24871
rect 12081 24837 12115 24871
rect 12115 24837 12124 24871
rect 12072 24828 12124 24837
rect 18604 24828 18656 24880
rect 22560 24828 22612 24880
rect 13176 24760 13228 24812
rect 14924 24803 14976 24812
rect 12532 24692 12584 24744
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 15844 24803 15896 24812
rect 15844 24769 15853 24803
rect 15853 24769 15887 24803
rect 15887 24769 15896 24803
rect 15844 24760 15896 24769
rect 16120 24760 16172 24812
rect 20812 24760 20864 24812
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 14188 24692 14240 24744
rect 18052 24735 18104 24744
rect 14280 24556 14332 24608
rect 15108 24599 15160 24608
rect 15108 24565 15117 24599
rect 15117 24565 15151 24599
rect 15151 24565 15160 24599
rect 15108 24556 15160 24565
rect 18052 24701 18061 24735
rect 18061 24701 18095 24735
rect 18095 24701 18104 24735
rect 18052 24692 18104 24701
rect 21180 24692 21232 24744
rect 26700 24760 26752 24812
rect 28448 24760 28500 24812
rect 28724 24760 28776 24812
rect 33600 24803 33652 24812
rect 33600 24769 33609 24803
rect 33609 24769 33643 24803
rect 33643 24769 33652 24803
rect 33600 24760 33652 24769
rect 38660 24760 38712 24812
rect 25228 24692 25280 24744
rect 33968 24692 34020 24744
rect 34244 24735 34296 24744
rect 34244 24701 34253 24735
rect 34253 24701 34287 24735
rect 34287 24701 34296 24735
rect 34244 24692 34296 24701
rect 24676 24624 24728 24676
rect 46296 24760 46348 24812
rect 46388 24803 46440 24812
rect 46388 24769 46397 24803
rect 46397 24769 46431 24803
rect 46431 24769 46440 24803
rect 46848 24803 46900 24812
rect 46388 24760 46440 24769
rect 46848 24769 46857 24803
rect 46857 24769 46891 24803
rect 46891 24769 46900 24803
rect 46848 24760 46900 24769
rect 46940 24803 46992 24812
rect 46940 24769 46949 24803
rect 46949 24769 46983 24803
rect 46983 24769 46992 24803
rect 46940 24760 46992 24769
rect 47492 24760 47544 24812
rect 47952 24760 48004 24812
rect 45928 24692 45980 24744
rect 46480 24692 46532 24744
rect 47584 24624 47636 24676
rect 19524 24599 19576 24608
rect 19524 24565 19533 24599
rect 19533 24565 19567 24599
rect 19567 24565 19576 24599
rect 19524 24556 19576 24565
rect 20260 24556 20312 24608
rect 25136 24599 25188 24608
rect 25136 24565 25145 24599
rect 25145 24565 25179 24599
rect 25179 24565 25188 24599
rect 25136 24556 25188 24565
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 29552 24556 29604 24608
rect 31668 24556 31720 24608
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13176 24352 13228 24404
rect 19432 24395 19484 24404
rect 19432 24361 19441 24395
rect 19441 24361 19475 24395
rect 19475 24361 19484 24395
rect 19432 24352 19484 24361
rect 21180 24395 21232 24404
rect 21180 24361 21189 24395
rect 21189 24361 21223 24395
rect 21223 24361 21232 24395
rect 21180 24352 21232 24361
rect 21272 24352 21324 24404
rect 10048 24327 10100 24336
rect 10048 24293 10057 24327
rect 10057 24293 10091 24327
rect 10091 24293 10100 24327
rect 10048 24284 10100 24293
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 12440 24284 12492 24336
rect 13084 24216 13136 24268
rect 15384 24284 15436 24336
rect 17408 24284 17460 24336
rect 19524 24284 19576 24336
rect 9128 24148 9180 24157
rect 12532 24148 12584 24200
rect 14280 24259 14332 24268
rect 14280 24225 14289 24259
rect 14289 24225 14323 24259
rect 14323 24225 14332 24259
rect 14280 24216 14332 24225
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 24400 24284 24452 24336
rect 29092 24284 29144 24336
rect 34244 24352 34296 24404
rect 43076 24352 43128 24404
rect 43444 24352 43496 24404
rect 48228 24352 48280 24404
rect 40224 24284 40276 24336
rect 25136 24259 25188 24268
rect 25136 24225 25145 24259
rect 25145 24225 25179 24259
rect 25179 24225 25188 24259
rect 25136 24216 25188 24225
rect 46020 24216 46072 24268
rect 47768 24284 47820 24336
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 3884 24080 3936 24132
rect 9680 24123 9732 24132
rect 9036 24012 9088 24064
rect 9680 24089 9689 24123
rect 9689 24089 9723 24123
rect 9723 24089 9732 24123
rect 9680 24080 9732 24089
rect 14004 24080 14056 24132
rect 14740 24080 14792 24132
rect 20812 24148 20864 24200
rect 21732 24148 21784 24200
rect 22008 24191 22060 24200
rect 22008 24157 22017 24191
rect 22017 24157 22051 24191
rect 22051 24157 22060 24191
rect 22008 24148 22060 24157
rect 23204 24191 23256 24200
rect 23204 24157 23213 24191
rect 23213 24157 23247 24191
rect 23247 24157 23256 24191
rect 23204 24148 23256 24157
rect 23296 24191 23348 24200
rect 23296 24157 23305 24191
rect 23305 24157 23339 24191
rect 23339 24157 23348 24191
rect 23480 24191 23532 24200
rect 23296 24148 23348 24157
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 26884 24148 26936 24200
rect 16764 24080 16816 24132
rect 24400 24080 24452 24132
rect 28448 24080 28500 24132
rect 28724 24080 28776 24132
rect 30012 24148 30064 24200
rect 29276 24080 29328 24132
rect 30380 24148 30432 24200
rect 31668 24191 31720 24200
rect 31668 24157 31677 24191
rect 31677 24157 31711 24191
rect 31711 24157 31720 24191
rect 31668 24148 31720 24157
rect 35072 24191 35124 24200
rect 35072 24157 35081 24191
rect 35081 24157 35115 24191
rect 35115 24157 35124 24191
rect 35072 24148 35124 24157
rect 36912 24191 36964 24200
rect 36912 24157 36921 24191
rect 36921 24157 36955 24191
rect 36955 24157 36964 24191
rect 36912 24148 36964 24157
rect 43076 24191 43128 24200
rect 43076 24157 43085 24191
rect 43085 24157 43119 24191
rect 43119 24157 43128 24191
rect 43076 24148 43128 24157
rect 43260 24191 43312 24200
rect 43260 24157 43269 24191
rect 43269 24157 43303 24191
rect 43303 24157 43312 24191
rect 43260 24148 43312 24157
rect 43904 24191 43956 24200
rect 43904 24157 43913 24191
rect 43913 24157 43947 24191
rect 43947 24157 43956 24191
rect 43904 24148 43956 24157
rect 35808 24080 35860 24132
rect 45560 24148 45612 24200
rect 47400 24080 47452 24132
rect 10140 24055 10192 24064
rect 10140 24021 10149 24055
rect 10149 24021 10183 24055
rect 10183 24021 10192 24055
rect 10140 24012 10192 24021
rect 10692 24055 10744 24064
rect 10692 24021 10701 24055
rect 10701 24021 10735 24055
rect 10735 24021 10744 24055
rect 10692 24012 10744 24021
rect 29644 24012 29696 24064
rect 30656 24012 30708 24064
rect 31760 24055 31812 24064
rect 31760 24021 31769 24055
rect 31769 24021 31803 24055
rect 31803 24021 31812 24055
rect 43996 24055 44048 24064
rect 31760 24012 31812 24021
rect 43996 24021 44005 24055
rect 44005 24021 44039 24055
rect 44039 24021 44048 24055
rect 43996 24012 44048 24021
rect 47676 24012 47728 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 9772 23808 9824 23860
rect 16764 23851 16816 23860
rect 16764 23817 16773 23851
rect 16773 23817 16807 23851
rect 16807 23817 16816 23851
rect 16764 23808 16816 23817
rect 22560 23808 22612 23860
rect 29276 23808 29328 23860
rect 35072 23808 35124 23860
rect 35808 23851 35860 23860
rect 35808 23817 35817 23851
rect 35817 23817 35851 23851
rect 35851 23817 35860 23851
rect 35808 23808 35860 23817
rect 11704 23672 11756 23724
rect 15384 23740 15436 23792
rect 23296 23740 23348 23792
rect 23848 23740 23900 23792
rect 15108 23672 15160 23724
rect 17500 23715 17552 23724
rect 17500 23681 17509 23715
rect 17509 23681 17543 23715
rect 17543 23681 17552 23715
rect 17500 23672 17552 23681
rect 20352 23672 20404 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 23204 23672 23256 23724
rect 26884 23740 26936 23792
rect 29184 23740 29236 23792
rect 34704 23740 34756 23792
rect 41052 23740 41104 23792
rect 43904 23808 43956 23860
rect 45560 23808 45612 23860
rect 43076 23740 43128 23792
rect 45652 23740 45704 23792
rect 46112 23740 46164 23792
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 13912 23604 13964 23656
rect 14004 23647 14056 23656
rect 14004 23613 14013 23647
rect 14013 23613 14047 23647
rect 14047 23613 14056 23647
rect 17868 23647 17920 23656
rect 14004 23604 14056 23613
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 18788 23604 18840 23656
rect 23112 23604 23164 23656
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 28816 23672 28868 23724
rect 24032 23604 24084 23656
rect 28264 23604 28316 23656
rect 28724 23604 28776 23656
rect 25688 23536 25740 23588
rect 29000 23672 29052 23724
rect 19524 23468 19576 23520
rect 24676 23468 24728 23520
rect 24860 23468 24912 23520
rect 27804 23511 27856 23520
rect 27804 23477 27813 23511
rect 27813 23477 27847 23511
rect 27847 23477 27856 23511
rect 27804 23468 27856 23477
rect 31668 23672 31720 23724
rect 33508 23715 33560 23724
rect 33508 23681 33517 23715
rect 33517 23681 33551 23715
rect 33551 23681 33560 23715
rect 33508 23672 33560 23681
rect 35440 23672 35492 23724
rect 35808 23672 35860 23724
rect 39212 23715 39264 23724
rect 39212 23681 39221 23715
rect 39221 23681 39255 23715
rect 39255 23681 39264 23715
rect 39212 23672 39264 23681
rect 40040 23715 40092 23724
rect 40040 23681 40049 23715
rect 40049 23681 40083 23715
rect 40083 23681 40092 23715
rect 40040 23672 40092 23681
rect 43168 23672 43220 23724
rect 43996 23715 44048 23724
rect 43996 23681 44005 23715
rect 44005 23681 44039 23715
rect 44039 23681 44048 23715
rect 43996 23672 44048 23681
rect 38384 23604 38436 23656
rect 40224 23647 40276 23656
rect 40224 23613 40233 23647
rect 40233 23613 40267 23647
rect 40267 23613 40276 23647
rect 40224 23604 40276 23613
rect 41880 23647 41932 23656
rect 41880 23613 41889 23647
rect 41889 23613 41923 23647
rect 41923 23613 41932 23647
rect 41880 23604 41932 23613
rect 46112 23604 46164 23656
rect 47952 23672 48004 23724
rect 42892 23536 42944 23588
rect 30012 23468 30064 23520
rect 40040 23468 40092 23520
rect 41420 23468 41472 23520
rect 45560 23511 45612 23520
rect 45560 23477 45569 23511
rect 45569 23477 45603 23511
rect 45603 23477 45612 23511
rect 45560 23468 45612 23477
rect 47400 23468 47452 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 10416 23264 10468 23316
rect 13084 23307 13136 23316
rect 13084 23273 13093 23307
rect 13093 23273 13127 23307
rect 13127 23273 13136 23307
rect 13084 23264 13136 23273
rect 18512 23264 18564 23316
rect 9036 23171 9088 23180
rect 9036 23137 9045 23171
rect 9045 23137 9079 23171
rect 9079 23137 9088 23171
rect 9036 23128 9088 23137
rect 14924 23128 14976 23180
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 13820 23060 13872 23112
rect 15108 23060 15160 23112
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 25412 23264 25464 23316
rect 24216 23196 24268 23248
rect 25044 23196 25096 23248
rect 25596 23264 25648 23316
rect 28724 23307 28776 23316
rect 25688 23239 25740 23248
rect 25688 23205 25697 23239
rect 25697 23205 25731 23239
rect 25731 23205 25740 23239
rect 25688 23196 25740 23205
rect 19524 23171 19576 23180
rect 19524 23137 19533 23171
rect 19533 23137 19567 23171
rect 19567 23137 19576 23171
rect 19524 23128 19576 23137
rect 24676 23128 24728 23180
rect 27804 23128 27856 23180
rect 21824 23103 21876 23112
rect 9588 22992 9640 23044
rect 10692 22992 10744 23044
rect 15936 23035 15988 23044
rect 11704 22924 11756 22976
rect 13636 22924 13688 22976
rect 15936 23001 15945 23035
rect 15945 23001 15979 23035
rect 15979 23001 15988 23035
rect 15936 22992 15988 23001
rect 18696 22992 18748 23044
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 23388 23060 23440 23112
rect 26240 23103 26292 23112
rect 26240 23069 26249 23103
rect 26249 23069 26283 23103
rect 26283 23069 26292 23103
rect 26240 23060 26292 23069
rect 28724 23273 28733 23307
rect 28733 23273 28767 23307
rect 28767 23273 28776 23307
rect 28724 23264 28776 23273
rect 28816 23264 28868 23316
rect 28264 23196 28316 23248
rect 28908 23239 28960 23248
rect 28908 23205 28917 23239
rect 28917 23205 28951 23239
rect 28951 23205 28960 23239
rect 28908 23196 28960 23205
rect 30380 23264 30432 23316
rect 32128 23307 32180 23316
rect 32128 23273 32137 23307
rect 32137 23273 32171 23307
rect 32171 23273 32180 23307
rect 32128 23264 32180 23273
rect 33968 23196 34020 23248
rect 46756 23264 46808 23316
rect 43904 23196 43956 23248
rect 29552 23171 29604 23180
rect 29552 23137 29561 23171
rect 29561 23137 29595 23171
rect 29595 23137 29604 23171
rect 29552 23128 29604 23137
rect 30656 23171 30708 23180
rect 30656 23137 30665 23171
rect 30665 23137 30699 23171
rect 30699 23137 30708 23171
rect 30656 23128 30708 23137
rect 40040 23171 40092 23180
rect 40040 23137 40049 23171
rect 40049 23137 40083 23171
rect 40083 23137 40092 23171
rect 40040 23128 40092 23137
rect 40132 23128 40184 23180
rect 20076 22992 20128 23044
rect 22836 22992 22888 23044
rect 24952 22992 25004 23044
rect 26976 22992 27028 23044
rect 27804 22992 27856 23044
rect 29276 22992 29328 23044
rect 16672 22924 16724 22976
rect 17316 22924 17368 22976
rect 19156 22924 19208 22976
rect 23572 22967 23624 22976
rect 23572 22933 23581 22967
rect 23581 22933 23615 22967
rect 23615 22933 23624 22967
rect 23572 22924 23624 22933
rect 24492 22924 24544 22976
rect 25688 22924 25740 22976
rect 27344 22924 27396 22976
rect 27436 22924 27488 22976
rect 28448 22924 28500 22976
rect 29644 23060 29696 23112
rect 30104 23060 30156 23112
rect 31760 23060 31812 23112
rect 33968 23103 34020 23112
rect 33968 23069 33977 23103
rect 33977 23069 34011 23103
rect 34011 23069 34020 23103
rect 33968 23060 34020 23069
rect 33508 22992 33560 23044
rect 41420 23060 41472 23112
rect 35532 22992 35584 23044
rect 43260 23103 43312 23112
rect 43260 23069 43269 23103
rect 43269 23069 43303 23103
rect 43303 23069 43312 23103
rect 43260 23060 43312 23069
rect 43444 23103 43496 23112
rect 43444 23069 43453 23103
rect 43453 23069 43487 23103
rect 43487 23069 43496 23103
rect 43444 23060 43496 23069
rect 44456 23103 44508 23112
rect 44456 23069 44465 23103
rect 44465 23069 44499 23103
rect 44499 23069 44508 23103
rect 44456 23060 44508 23069
rect 45284 23035 45336 23044
rect 41604 22967 41656 22976
rect 41604 22933 41613 22967
rect 41613 22933 41647 22967
rect 41647 22933 41656 22967
rect 41604 22924 41656 22933
rect 45284 23001 45293 23035
rect 45293 23001 45327 23035
rect 45327 23001 45336 23035
rect 45284 22992 45336 23001
rect 45652 23128 45704 23180
rect 46940 23171 46992 23180
rect 46940 23137 46949 23171
rect 46949 23137 46983 23171
rect 46983 23137 46992 23171
rect 46940 23128 46992 23137
rect 47492 22992 47544 23044
rect 46572 22924 46624 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9588 22763 9640 22772
rect 9588 22729 9597 22763
rect 9597 22729 9631 22763
rect 9631 22729 9640 22763
rect 9588 22720 9640 22729
rect 13912 22763 13964 22772
rect 13912 22729 13921 22763
rect 13921 22729 13955 22763
rect 13955 22729 13964 22763
rect 13912 22720 13964 22729
rect 11704 22695 11756 22704
rect 11704 22661 11713 22695
rect 11713 22661 11747 22695
rect 11747 22661 11756 22695
rect 11704 22652 11756 22661
rect 10140 22584 10192 22636
rect 10784 22584 10836 22636
rect 11336 22448 11388 22500
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 14924 22584 14976 22636
rect 15108 22584 15160 22636
rect 18604 22652 18656 22704
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 19892 22627 19944 22636
rect 19892 22593 19901 22627
rect 19901 22593 19935 22627
rect 19935 22593 19944 22627
rect 19892 22584 19944 22593
rect 21824 22720 21876 22772
rect 22836 22763 22888 22772
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 24860 22720 24912 22772
rect 26976 22720 27028 22772
rect 24492 22695 24544 22704
rect 21824 22627 21876 22636
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 24492 22661 24501 22695
rect 24501 22661 24535 22695
rect 24535 22661 24544 22695
rect 24492 22652 24544 22661
rect 22284 22584 22336 22636
rect 22836 22584 22888 22636
rect 23572 22627 23624 22636
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 23848 22584 23900 22636
rect 26884 22652 26936 22704
rect 27436 22763 27488 22772
rect 27436 22729 27445 22763
rect 27445 22729 27479 22763
rect 27479 22729 27488 22763
rect 29184 22763 29236 22772
rect 27436 22720 27488 22729
rect 29184 22729 29193 22763
rect 29193 22729 29227 22763
rect 29227 22729 29236 22763
rect 29184 22720 29236 22729
rect 30104 22763 30156 22772
rect 30104 22729 30113 22763
rect 30113 22729 30147 22763
rect 30147 22729 30156 22763
rect 30104 22720 30156 22729
rect 40224 22720 40276 22772
rect 43076 22763 43128 22772
rect 43076 22729 43085 22763
rect 43085 22729 43119 22763
rect 43119 22729 43128 22763
rect 43076 22720 43128 22729
rect 44456 22720 44508 22772
rect 28908 22652 28960 22704
rect 25504 22627 25556 22636
rect 25504 22593 25513 22627
rect 25513 22593 25547 22627
rect 25547 22593 25556 22627
rect 25504 22584 25556 22593
rect 25688 22627 25740 22636
rect 25688 22593 25697 22627
rect 25697 22593 25731 22627
rect 25731 22593 25740 22627
rect 25688 22584 25740 22593
rect 26516 22584 26568 22636
rect 27160 22584 27212 22636
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 17224 22559 17276 22568
rect 17224 22525 17233 22559
rect 17233 22525 17267 22559
rect 17267 22525 17276 22559
rect 17224 22516 17276 22525
rect 15200 22491 15252 22500
rect 15200 22457 15209 22491
rect 15209 22457 15243 22491
rect 15243 22457 15252 22491
rect 15200 22448 15252 22457
rect 15384 22448 15436 22500
rect 21824 22448 21876 22500
rect 22744 22448 22796 22500
rect 24676 22516 24728 22568
rect 25780 22559 25832 22568
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 27068 22516 27120 22568
rect 29092 22627 29144 22636
rect 29092 22593 29101 22627
rect 29101 22593 29135 22627
rect 29135 22593 29144 22627
rect 29092 22584 29144 22593
rect 45560 22652 45612 22704
rect 29828 22584 29880 22636
rect 40224 22584 40276 22636
rect 27712 22559 27764 22568
rect 27712 22525 27721 22559
rect 27721 22525 27755 22559
rect 27755 22525 27764 22559
rect 27712 22516 27764 22525
rect 43444 22584 43496 22636
rect 45100 22584 45152 22636
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 43260 22516 43312 22568
rect 43720 22516 43772 22568
rect 44180 22559 44232 22568
rect 25044 22448 25096 22500
rect 25872 22448 25924 22500
rect 26148 22448 26200 22500
rect 41604 22448 41656 22500
rect 44180 22525 44189 22559
rect 44189 22525 44223 22559
rect 44223 22525 44232 22559
rect 44180 22516 44232 22525
rect 46940 22559 46992 22568
rect 46940 22525 46949 22559
rect 46949 22525 46983 22559
rect 46983 22525 46992 22559
rect 46940 22516 46992 22525
rect 47860 22559 47912 22568
rect 47860 22525 47869 22559
rect 47869 22525 47903 22559
rect 47903 22525 47912 22559
rect 47860 22516 47912 22525
rect 46848 22448 46900 22500
rect 16304 22380 16356 22432
rect 16488 22380 16540 22432
rect 20168 22380 20220 22432
rect 24400 22380 24452 22432
rect 24768 22380 24820 22432
rect 27252 22380 27304 22432
rect 27344 22380 27396 22432
rect 40040 22423 40092 22432
rect 40040 22389 40049 22423
rect 40049 22389 40083 22423
rect 40083 22389 40092 22423
rect 40040 22380 40092 22389
rect 41880 22380 41932 22432
rect 46940 22380 46992 22432
rect 47676 22423 47728 22432
rect 47676 22389 47685 22423
rect 47685 22389 47719 22423
rect 47719 22389 47728 22423
rect 47676 22380 47728 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 15936 22176 15988 22228
rect 17224 22176 17276 22228
rect 19892 22176 19944 22228
rect 26148 22176 26200 22228
rect 26240 22176 26292 22228
rect 27068 22176 27120 22228
rect 27528 22176 27580 22228
rect 28816 22176 28868 22228
rect 30012 22176 30064 22228
rect 13084 22108 13136 22160
rect 11888 22040 11940 22092
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 12532 21972 12584 22024
rect 9956 21904 10008 21956
rect 11060 21904 11112 21956
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 13820 21836 13872 21888
rect 14280 21879 14332 21888
rect 14280 21845 14289 21879
rect 14289 21845 14323 21879
rect 14323 21845 14332 21879
rect 14280 21836 14332 21845
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 15200 21972 15252 22024
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 17500 22108 17552 22160
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 26424 22108 26476 22160
rect 27620 22108 27672 22160
rect 16304 21904 16356 21956
rect 17684 21904 17736 21956
rect 19156 21972 19208 22024
rect 19984 22015 20036 22024
rect 19984 21981 19993 22015
rect 19993 21981 20027 22015
rect 20027 21981 20036 22015
rect 19984 21972 20036 21981
rect 23756 21972 23808 22024
rect 24676 22015 24728 22024
rect 20996 21904 21048 21956
rect 24216 21904 24268 21956
rect 24400 21947 24452 21956
rect 24400 21913 24409 21947
rect 24409 21913 24443 21947
rect 24443 21913 24452 21947
rect 24400 21904 24452 21913
rect 24676 21981 24685 22015
rect 24685 21981 24719 22015
rect 24719 21981 24728 22015
rect 24676 21972 24728 21981
rect 26148 22015 26200 22024
rect 26148 21981 26157 22015
rect 26157 21981 26191 22015
rect 26191 21981 26200 22015
rect 26148 21972 26200 21981
rect 26424 21972 26476 22024
rect 29644 21972 29696 22024
rect 24860 21904 24912 21956
rect 27436 21904 27488 21956
rect 27620 21904 27672 21956
rect 37280 21904 37332 21956
rect 40040 21972 40092 22024
rect 40224 21904 40276 21956
rect 40500 21904 40552 21956
rect 41696 22040 41748 22092
rect 42524 22015 42576 22024
rect 42524 21981 42533 22015
rect 42533 21981 42567 22015
rect 42567 21981 42576 22015
rect 42524 21972 42576 21981
rect 45560 22040 45612 22092
rect 44548 21972 44600 22024
rect 45284 21972 45336 22024
rect 47032 21972 47084 22024
rect 42248 21904 42300 21956
rect 42432 21904 42484 21956
rect 44180 21904 44232 21956
rect 44272 21947 44324 21956
rect 44272 21913 44281 21947
rect 44281 21913 44315 21947
rect 44315 21913 44324 21947
rect 44272 21904 44324 21913
rect 45928 21904 45980 21956
rect 46020 21904 46072 21956
rect 20076 21836 20128 21888
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 23848 21836 23900 21888
rect 27712 21879 27764 21888
rect 27712 21845 27737 21879
rect 27737 21845 27764 21879
rect 27896 21879 27948 21888
rect 27712 21836 27764 21845
rect 27896 21845 27905 21879
rect 27905 21845 27939 21879
rect 27939 21845 27948 21879
rect 27896 21836 27948 21845
rect 42340 21836 42392 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 11336 21564 11388 21616
rect 10416 21496 10468 21548
rect 12532 21564 12584 21616
rect 16948 21564 17000 21616
rect 20996 21607 21048 21616
rect 20996 21573 21005 21607
rect 21005 21573 21039 21607
rect 21039 21573 21048 21607
rect 20996 21564 21048 21573
rect 14280 21539 14332 21548
rect 2872 21428 2924 21480
rect 14280 21505 14289 21539
rect 14289 21505 14323 21539
rect 14323 21505 14332 21539
rect 14280 21496 14332 21505
rect 15660 21496 15712 21548
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 21824 21539 21876 21548
rect 11888 21471 11940 21480
rect 11888 21437 11897 21471
rect 11897 21437 11931 21471
rect 11931 21437 11940 21471
rect 11888 21428 11940 21437
rect 11980 21428 12032 21480
rect 14556 21471 14608 21480
rect 9312 21335 9364 21344
rect 9312 21301 9321 21335
rect 9321 21301 9355 21335
rect 9355 21301 9364 21335
rect 9312 21292 9364 21301
rect 9588 21292 9640 21344
rect 12532 21292 12584 21344
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 19432 21428 19484 21480
rect 20168 21428 20220 21480
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 22744 21539 22796 21548
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 23848 21564 23900 21616
rect 26976 21564 27028 21616
rect 27528 21675 27580 21684
rect 27528 21641 27553 21675
rect 27553 21641 27580 21675
rect 27712 21675 27764 21684
rect 27528 21632 27580 21641
rect 27712 21641 27721 21675
rect 27721 21641 27755 21675
rect 27755 21641 27764 21675
rect 27712 21632 27764 21641
rect 42432 21632 42484 21684
rect 43168 21632 43220 21684
rect 47492 21632 47544 21684
rect 24768 21496 24820 21548
rect 20352 21403 20404 21412
rect 20352 21369 20361 21403
rect 20361 21369 20395 21403
rect 20395 21369 20404 21403
rect 26148 21496 26200 21548
rect 29644 21496 29696 21548
rect 29828 21496 29880 21548
rect 20352 21360 20404 21369
rect 26056 21360 26108 21412
rect 29828 21360 29880 21412
rect 14740 21292 14792 21344
rect 16028 21335 16080 21344
rect 16028 21301 16037 21335
rect 16037 21301 16071 21335
rect 16071 21301 16080 21335
rect 16028 21292 16080 21301
rect 19984 21292 20036 21344
rect 21088 21292 21140 21344
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 23480 21292 23532 21344
rect 26884 21292 26936 21344
rect 27528 21335 27580 21344
rect 27528 21301 27537 21335
rect 27537 21301 27571 21335
rect 27571 21301 27580 21335
rect 27528 21292 27580 21301
rect 32036 21564 32088 21616
rect 41696 21539 41748 21548
rect 41696 21505 41705 21539
rect 41705 21505 41739 21539
rect 41739 21505 41748 21539
rect 41696 21496 41748 21505
rect 42524 21496 42576 21548
rect 42708 21496 42760 21548
rect 43260 21539 43312 21548
rect 43260 21505 43269 21539
rect 43269 21505 43303 21539
rect 43303 21505 43312 21539
rect 45744 21564 45796 21616
rect 47216 21564 47268 21616
rect 43260 21496 43312 21505
rect 44548 21539 44600 21548
rect 44548 21505 44557 21539
rect 44557 21505 44591 21539
rect 44591 21505 44600 21539
rect 44548 21496 44600 21505
rect 45376 21496 45428 21548
rect 47860 21539 47912 21548
rect 47860 21505 47869 21539
rect 47869 21505 47903 21539
rect 47903 21505 47912 21539
rect 47860 21496 47912 21505
rect 48044 21496 48096 21548
rect 32128 21471 32180 21480
rect 32128 21437 32137 21471
rect 32137 21437 32171 21471
rect 32171 21437 32180 21471
rect 32128 21428 32180 21437
rect 32588 21471 32640 21480
rect 30196 21360 30248 21412
rect 32588 21437 32597 21471
rect 32597 21437 32631 21471
rect 32631 21437 32640 21471
rect 32588 21428 32640 21437
rect 45008 21428 45060 21480
rect 46204 21471 46256 21480
rect 46204 21437 46213 21471
rect 46213 21437 46247 21471
rect 46247 21437 46256 21471
rect 46204 21428 46256 21437
rect 34796 21292 34848 21344
rect 40224 21292 40276 21344
rect 42248 21292 42300 21344
rect 46756 21292 46808 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 11888 21088 11940 21140
rect 3516 21020 3568 21072
rect 26056 21088 26108 21140
rect 9588 20995 9640 21004
rect 9588 20961 9597 20995
rect 9597 20961 9631 20995
rect 9631 20961 9640 20995
rect 9588 20952 9640 20961
rect 10140 20952 10192 21004
rect 14556 21020 14608 21072
rect 15660 21020 15712 21072
rect 9128 20884 9180 20936
rect 11980 20816 12032 20868
rect 12532 20884 12584 20936
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 23112 20952 23164 21004
rect 27252 21088 27304 21140
rect 29552 21088 29604 21140
rect 30104 20952 30156 21004
rect 30196 20952 30248 21004
rect 31208 21131 31260 21140
rect 31208 21097 31217 21131
rect 31217 21097 31251 21131
rect 31251 21097 31260 21131
rect 31208 21088 31260 21097
rect 32036 21131 32088 21140
rect 32036 21097 32045 21131
rect 32045 21097 32079 21131
rect 32079 21097 32088 21131
rect 32036 21088 32088 21097
rect 34796 21131 34848 21140
rect 34796 21097 34805 21131
rect 34805 21097 34839 21131
rect 34839 21097 34848 21131
rect 34796 21088 34848 21097
rect 14464 20927 14516 20936
rect 12716 20816 12768 20868
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 14464 20884 14516 20893
rect 16304 20884 16356 20936
rect 19432 20884 19484 20936
rect 26240 20884 26292 20936
rect 26884 20927 26936 20936
rect 26884 20893 26893 20927
rect 26893 20893 26927 20927
rect 26927 20893 26936 20927
rect 26884 20884 26936 20893
rect 14372 20816 14424 20868
rect 22100 20816 22152 20868
rect 27804 20816 27856 20868
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 22744 20748 22796 20800
rect 27528 20748 27580 20800
rect 29368 20748 29420 20800
rect 36360 20952 36412 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 35624 20884 35676 20936
rect 42340 20927 42392 20936
rect 34796 20816 34848 20868
rect 42340 20893 42349 20927
rect 42349 20893 42383 20927
rect 42383 20893 42392 20927
rect 42340 20884 42392 20893
rect 43260 20927 43312 20936
rect 43260 20893 43269 20927
rect 43269 20893 43303 20927
rect 43303 20893 43312 20927
rect 43260 20884 43312 20893
rect 43628 20884 43680 20936
rect 45376 20927 45428 20936
rect 45376 20893 45385 20927
rect 45385 20893 45419 20927
rect 45419 20893 45428 20927
rect 45376 20884 45428 20893
rect 42708 20816 42760 20868
rect 45744 20816 45796 20868
rect 46480 20859 46532 20868
rect 46480 20825 46489 20859
rect 46489 20825 46523 20859
rect 46523 20825 46532 20859
rect 46480 20816 46532 20825
rect 43904 20791 43956 20800
rect 43904 20757 43913 20791
rect 43913 20757 43947 20791
rect 43947 20757 43956 20791
rect 43904 20748 43956 20757
rect 47216 20748 47268 20800
rect 47860 20748 47912 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3424 20544 3476 20596
rect 9312 20519 9364 20528
rect 9312 20485 9321 20519
rect 9321 20485 9355 20519
rect 9355 20485 9364 20519
rect 9312 20476 9364 20485
rect 11980 20476 12032 20528
rect 12532 20519 12584 20528
rect 12532 20485 12557 20519
rect 12557 20485 12584 20519
rect 12716 20587 12768 20596
rect 12716 20553 12725 20587
rect 12725 20553 12759 20587
rect 12759 20553 12768 20587
rect 12716 20544 12768 20553
rect 14464 20544 14516 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 16580 20544 16632 20596
rect 22100 20587 22152 20596
rect 22100 20553 22109 20587
rect 22109 20553 22143 20587
rect 22143 20553 22152 20587
rect 22100 20544 22152 20553
rect 26240 20544 26292 20596
rect 27528 20544 27580 20596
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 12532 20476 12584 20485
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 12440 20408 12492 20460
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 15016 20408 15068 20460
rect 16120 20408 16172 20460
rect 3976 20272 4028 20324
rect 14556 20383 14608 20392
rect 14556 20349 14565 20383
rect 14565 20349 14599 20383
rect 14599 20349 14608 20383
rect 14832 20383 14884 20392
rect 14556 20340 14608 20349
rect 14832 20349 14841 20383
rect 14841 20349 14875 20383
rect 14875 20349 14884 20383
rect 14832 20340 14884 20349
rect 16672 20340 16724 20392
rect 17040 20417 17049 20426
rect 17049 20417 17083 20426
rect 17083 20417 17092 20426
rect 17040 20374 17092 20417
rect 15200 20272 15252 20324
rect 16028 20272 16080 20324
rect 16764 20315 16816 20324
rect 16764 20281 16773 20315
rect 16773 20281 16807 20315
rect 16807 20281 16816 20315
rect 16764 20272 16816 20281
rect 11428 20204 11480 20256
rect 12256 20204 12308 20256
rect 14372 20204 14424 20256
rect 19340 20476 19392 20528
rect 23480 20476 23532 20528
rect 23664 20476 23716 20528
rect 26516 20476 26568 20528
rect 26884 20476 26936 20528
rect 22836 20408 22888 20460
rect 25872 20451 25924 20460
rect 19248 20340 19300 20392
rect 22928 20383 22980 20392
rect 22928 20349 22937 20383
rect 22937 20349 22971 20383
rect 22971 20349 22980 20383
rect 22928 20340 22980 20349
rect 24400 20340 24452 20392
rect 25872 20417 25881 20451
rect 25881 20417 25915 20451
rect 25915 20417 25924 20451
rect 25872 20408 25924 20417
rect 26976 20451 27028 20460
rect 26976 20417 26985 20451
rect 26985 20417 27019 20451
rect 27019 20417 27028 20451
rect 26976 20408 27028 20417
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 28356 20476 28408 20528
rect 27252 20408 27304 20417
rect 30932 20408 30984 20460
rect 25688 20247 25740 20256
rect 25688 20213 25697 20247
rect 25697 20213 25731 20247
rect 25731 20213 25740 20247
rect 25688 20204 25740 20213
rect 32128 20408 32180 20460
rect 36360 20451 36412 20460
rect 36360 20417 36369 20451
rect 36369 20417 36403 20451
rect 36403 20417 36412 20451
rect 36360 20408 36412 20417
rect 41696 20408 41748 20460
rect 42800 20408 42852 20460
rect 43076 20408 43128 20460
rect 33140 20340 33192 20392
rect 34152 20383 34204 20392
rect 34152 20349 34161 20383
rect 34161 20349 34195 20383
rect 34195 20349 34204 20383
rect 34152 20340 34204 20349
rect 35716 20383 35768 20392
rect 35716 20349 35725 20383
rect 35725 20349 35759 20383
rect 35759 20349 35768 20383
rect 35716 20340 35768 20349
rect 43168 20340 43220 20392
rect 45560 20476 45612 20528
rect 47032 20544 47084 20596
rect 42708 20315 42760 20324
rect 42708 20281 42717 20315
rect 42717 20281 42751 20315
rect 42751 20281 42760 20315
rect 42708 20272 42760 20281
rect 42984 20272 43036 20324
rect 43904 20340 43956 20392
rect 47032 20383 47084 20392
rect 47032 20349 47041 20383
rect 47041 20349 47075 20383
rect 47075 20349 47084 20383
rect 47032 20340 47084 20349
rect 47676 20476 47728 20528
rect 47492 20408 47544 20460
rect 47952 20340 48004 20392
rect 43812 20272 43864 20324
rect 37280 20204 37332 20256
rect 44180 20204 44232 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 9128 20000 9180 20052
rect 12256 20000 12308 20052
rect 15016 20043 15068 20052
rect 15016 20009 15025 20043
rect 15025 20009 15059 20043
rect 15059 20009 15068 20043
rect 15016 20000 15068 20009
rect 17040 20000 17092 20052
rect 22928 20043 22980 20052
rect 22928 20009 22937 20043
rect 22937 20009 22971 20043
rect 22971 20009 22980 20043
rect 22928 20000 22980 20009
rect 23664 20000 23716 20052
rect 43628 20043 43680 20052
rect 15200 19932 15252 19984
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 18696 19932 18748 19984
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 18052 19864 18104 19916
rect 18512 19864 18564 19916
rect 1768 19796 1820 19848
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 11428 19728 11480 19780
rect 10416 19660 10468 19712
rect 12256 19796 12308 19848
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 16764 19796 16816 19848
rect 13820 19728 13872 19780
rect 14740 19771 14792 19780
rect 14740 19737 14749 19771
rect 14749 19737 14783 19771
rect 14783 19737 14792 19771
rect 14740 19728 14792 19737
rect 16120 19771 16172 19780
rect 16120 19737 16129 19771
rect 16129 19737 16163 19771
rect 16163 19737 16172 19771
rect 16120 19728 16172 19737
rect 16672 19728 16724 19780
rect 18328 19796 18380 19848
rect 20076 19796 20128 19848
rect 20996 19864 21048 19916
rect 25688 19907 25740 19916
rect 20904 19796 20956 19848
rect 22836 19796 22888 19848
rect 25688 19873 25697 19907
rect 25697 19873 25731 19907
rect 25731 19873 25740 19907
rect 25688 19864 25740 19873
rect 24860 19796 24912 19848
rect 29644 19796 29696 19848
rect 30196 19932 30248 19984
rect 30932 19975 30984 19984
rect 30932 19941 30941 19975
rect 30941 19941 30975 19975
rect 30975 19941 30984 19975
rect 30932 19932 30984 19941
rect 43628 20009 43637 20043
rect 43637 20009 43671 20043
rect 43671 20009 43680 20043
rect 43628 20000 43680 20009
rect 46480 20000 46532 20052
rect 34152 19932 34204 19984
rect 34796 19932 34848 19984
rect 46664 19932 46716 19984
rect 30012 19796 30064 19848
rect 35716 19864 35768 19916
rect 47032 19907 47084 19916
rect 33600 19796 33652 19848
rect 47032 19873 47041 19907
rect 47041 19873 47075 19907
rect 47075 19873 47084 19907
rect 47032 19864 47084 19873
rect 42984 19839 43036 19848
rect 42984 19805 42993 19839
rect 42993 19805 43027 19839
rect 43027 19805 43036 19839
rect 42984 19796 43036 19805
rect 43168 19839 43220 19848
rect 43168 19805 43177 19839
rect 43177 19805 43211 19839
rect 43211 19805 43220 19839
rect 43168 19796 43220 19805
rect 43812 19839 43864 19848
rect 43812 19805 43821 19839
rect 43821 19805 43855 19839
rect 43855 19805 43864 19839
rect 43812 19796 43864 19805
rect 44548 19796 44600 19848
rect 45008 19796 45060 19848
rect 45652 19796 45704 19848
rect 19248 19728 19300 19780
rect 27068 19728 27120 19780
rect 29828 19728 29880 19780
rect 35624 19728 35676 19780
rect 46112 19771 46164 19780
rect 46112 19737 46121 19771
rect 46121 19737 46155 19771
rect 46155 19737 46164 19771
rect 46112 19728 46164 19737
rect 11704 19660 11756 19712
rect 13452 19660 13504 19712
rect 14556 19660 14608 19712
rect 17776 19660 17828 19712
rect 20812 19703 20864 19712
rect 20812 19669 20821 19703
rect 20821 19669 20855 19703
rect 20855 19669 20864 19703
rect 20812 19660 20864 19669
rect 26516 19660 26568 19712
rect 26976 19660 27028 19712
rect 33876 19703 33928 19712
rect 33876 19669 33885 19703
rect 33885 19669 33919 19703
rect 33919 19669 33928 19703
rect 33876 19660 33928 19669
rect 33968 19660 34020 19712
rect 38292 19660 38344 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 9864 19456 9916 19508
rect 27068 19499 27120 19508
rect 4896 19388 4948 19440
rect 12440 19388 12492 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 15752 19388 15804 19440
rect 16120 19431 16172 19440
rect 16120 19397 16129 19431
rect 16129 19397 16163 19431
rect 16163 19397 16172 19431
rect 16120 19388 16172 19397
rect 19340 19388 19392 19440
rect 23112 19388 23164 19440
rect 27068 19465 27077 19499
rect 27077 19465 27111 19499
rect 27111 19465 27120 19499
rect 27068 19456 27120 19465
rect 30012 19456 30064 19508
rect 29000 19388 29052 19440
rect 29828 19388 29880 19440
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 12716 19252 12768 19304
rect 16672 19320 16724 19372
rect 13452 19252 13504 19304
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 16764 19252 16816 19304
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 17776 19363 17828 19372
rect 16948 19320 17000 19329
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 20076 19320 20128 19372
rect 24400 19320 24452 19372
rect 24768 19320 24820 19372
rect 26884 19320 26936 19372
rect 29644 19320 29696 19372
rect 33140 19320 33192 19372
rect 33876 19431 33928 19440
rect 33876 19397 33885 19431
rect 33885 19397 33919 19431
rect 33919 19397 33928 19431
rect 33876 19388 33928 19397
rect 38292 19456 38344 19508
rect 45928 19456 45980 19508
rect 43904 19388 43956 19440
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 18052 19295 18104 19304
rect 17132 19252 17184 19261
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 19248 19252 19300 19304
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 35532 19363 35584 19372
rect 35532 19329 35541 19363
rect 35541 19329 35575 19363
rect 35575 19329 35584 19363
rect 35532 19320 35584 19329
rect 37280 19363 37332 19372
rect 37280 19329 37289 19363
rect 37289 19329 37323 19363
rect 37323 19329 37332 19363
rect 37280 19320 37332 19329
rect 39120 19363 39172 19372
rect 39120 19329 39129 19363
rect 39129 19329 39163 19363
rect 39163 19329 39172 19363
rect 39120 19320 39172 19329
rect 44548 19363 44600 19372
rect 44548 19329 44557 19363
rect 44557 19329 44591 19363
rect 44591 19329 44600 19363
rect 44548 19320 44600 19329
rect 22100 19252 22152 19261
rect 33968 19252 34020 19304
rect 37464 19295 37516 19304
rect 37464 19261 37473 19295
rect 37473 19261 37507 19295
rect 37507 19261 37516 19295
rect 37464 19252 37516 19261
rect 44088 19252 44140 19304
rect 45100 19295 45152 19304
rect 45100 19261 45109 19295
rect 45109 19261 45143 19295
rect 45143 19261 45152 19295
rect 45100 19252 45152 19261
rect 47124 19456 47176 19508
rect 46112 19388 46164 19440
rect 46388 19363 46440 19372
rect 46388 19329 46397 19363
rect 46397 19329 46431 19363
rect 46431 19329 46440 19363
rect 46388 19320 46440 19329
rect 3976 19184 4028 19236
rect 11980 19116 12032 19168
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 14740 19159 14792 19168
rect 14740 19125 14749 19159
rect 14749 19125 14783 19159
rect 14783 19125 14792 19159
rect 14740 19116 14792 19125
rect 17316 19116 17368 19168
rect 20904 19159 20956 19168
rect 20904 19125 20913 19159
rect 20913 19125 20947 19159
rect 20947 19125 20956 19159
rect 20904 19116 20956 19125
rect 23388 19184 23440 19236
rect 31024 19184 31076 19236
rect 33140 19184 33192 19236
rect 24308 19159 24360 19168
rect 24308 19125 24317 19159
rect 24317 19125 24351 19159
rect 24351 19125 24360 19159
rect 24308 19116 24360 19125
rect 32312 19116 32364 19168
rect 33048 19159 33100 19168
rect 33048 19125 33057 19159
rect 33057 19125 33091 19159
rect 33091 19125 33100 19159
rect 33048 19116 33100 19125
rect 43628 19159 43680 19168
rect 43628 19125 43637 19159
rect 43637 19125 43671 19159
rect 43671 19125 43680 19159
rect 43628 19116 43680 19125
rect 45928 19184 45980 19236
rect 47676 19320 47728 19372
rect 48044 19252 48096 19304
rect 47768 19184 47820 19236
rect 46388 19116 46440 19168
rect 47400 19116 47452 19168
rect 47676 19116 47728 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 2136 18844 2188 18896
rect 6644 18912 6696 18964
rect 46020 18912 46072 18964
rect 15752 18844 15804 18896
rect 17040 18844 17092 18896
rect 17316 18887 17368 18896
rect 17316 18853 17325 18887
rect 17325 18853 17359 18887
rect 17359 18853 17368 18887
rect 17316 18844 17368 18853
rect 17684 18844 17736 18896
rect 17868 18844 17920 18896
rect 19340 18887 19392 18896
rect 19340 18853 19349 18887
rect 19349 18853 19383 18887
rect 19383 18853 19392 18887
rect 19340 18844 19392 18853
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 11980 18819 12032 18828
rect 11980 18785 11989 18819
rect 11989 18785 12023 18819
rect 12023 18785 12032 18819
rect 11980 18776 12032 18785
rect 14740 18819 14792 18828
rect 14740 18785 14749 18819
rect 14749 18785 14783 18819
rect 14783 18785 14792 18819
rect 14740 18776 14792 18785
rect 16764 18776 16816 18828
rect 17132 18776 17184 18828
rect 20076 18776 20128 18828
rect 20812 18819 20864 18828
rect 20812 18785 20821 18819
rect 20821 18785 20855 18819
rect 20855 18785 20864 18819
rect 20812 18776 20864 18785
rect 23112 18844 23164 18896
rect 24400 18844 24452 18896
rect 37464 18844 37516 18896
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 13084 18708 13136 18760
rect 14096 18708 14148 18760
rect 15844 18708 15896 18760
rect 17224 18708 17276 18760
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 22836 18708 22888 18760
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 16304 18572 16356 18624
rect 22376 18640 22428 18692
rect 25044 18776 25096 18828
rect 26516 18819 26568 18828
rect 24400 18640 24452 18692
rect 25780 18708 25832 18760
rect 26516 18785 26525 18819
rect 26525 18785 26559 18819
rect 26559 18785 26568 18819
rect 26516 18776 26568 18785
rect 31024 18819 31076 18828
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 30012 18708 30064 18760
rect 31024 18785 31033 18819
rect 31033 18785 31067 18819
rect 31067 18785 31076 18819
rect 31024 18776 31076 18785
rect 33048 18776 33100 18828
rect 47768 18844 47820 18896
rect 30564 18751 30616 18760
rect 30564 18717 30573 18751
rect 30573 18717 30607 18751
rect 30607 18717 30616 18751
rect 30564 18708 30616 18717
rect 33140 18751 33192 18760
rect 17592 18572 17644 18624
rect 18052 18572 18104 18624
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 23296 18572 23348 18624
rect 24584 18572 24636 18624
rect 28356 18683 28408 18692
rect 28356 18649 28365 18683
rect 28365 18649 28399 18683
rect 28399 18649 28408 18683
rect 28356 18640 28408 18649
rect 31024 18640 31076 18692
rect 26240 18572 26292 18624
rect 26884 18572 26936 18624
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 43628 18776 43680 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 33968 18708 34020 18760
rect 37096 18751 37148 18760
rect 37096 18717 37105 18751
rect 37105 18717 37139 18751
rect 37139 18717 37148 18751
rect 37096 18708 37148 18717
rect 43812 18708 43864 18760
rect 44180 18751 44232 18760
rect 44180 18717 44189 18751
rect 44189 18717 44223 18751
rect 44223 18717 44232 18751
rect 44180 18708 44232 18717
rect 45192 18751 45244 18760
rect 45192 18717 45201 18751
rect 45201 18717 45235 18751
rect 45235 18717 45244 18751
rect 45192 18708 45244 18717
rect 45376 18751 45428 18760
rect 45376 18717 45385 18751
rect 45385 18717 45419 18751
rect 45419 18717 45428 18751
rect 45376 18708 45428 18717
rect 34612 18640 34664 18692
rect 44088 18683 44140 18692
rect 44088 18649 44097 18683
rect 44097 18649 44131 18683
rect 44131 18649 44140 18683
rect 44088 18640 44140 18649
rect 47676 18640 47728 18692
rect 37096 18572 37148 18624
rect 45008 18572 45060 18624
rect 45284 18615 45336 18624
rect 45284 18581 45293 18615
rect 45293 18581 45327 18615
rect 45327 18581 45336 18615
rect 45284 18572 45336 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1584 18368 1636 18420
rect 14096 18411 14148 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 14096 18377 14105 18411
rect 14105 18377 14139 18411
rect 14139 18377 14148 18411
rect 14096 18368 14148 18377
rect 15844 18411 15896 18420
rect 15844 18377 15853 18411
rect 15853 18377 15887 18411
rect 15887 18377 15896 18411
rect 15844 18368 15896 18377
rect 3332 18300 3384 18352
rect 18420 18368 18472 18420
rect 13820 18232 13872 18284
rect 16304 18232 16356 18284
rect 19984 18300 20036 18352
rect 21824 18368 21876 18420
rect 26884 18368 26936 18420
rect 28816 18368 28868 18420
rect 31024 18411 31076 18420
rect 31024 18377 31033 18411
rect 31033 18377 31067 18411
rect 31067 18377 31076 18411
rect 31024 18368 31076 18377
rect 44456 18368 44508 18420
rect 47676 18411 47728 18420
rect 23296 18343 23348 18352
rect 23296 18309 23305 18343
rect 23305 18309 23339 18343
rect 23339 18309 23348 18343
rect 23296 18300 23348 18309
rect 28540 18300 28592 18352
rect 30564 18300 30616 18352
rect 32312 18343 32364 18352
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 20904 18232 20956 18284
rect 24860 18232 24912 18284
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 28816 18232 28868 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 32312 18309 32321 18343
rect 32321 18309 32355 18343
rect 32355 18309 32364 18343
rect 32312 18300 32364 18309
rect 34612 18343 34664 18352
rect 34612 18309 34621 18343
rect 34621 18309 34655 18343
rect 34655 18309 34664 18343
rect 34612 18300 34664 18309
rect 33600 18232 33652 18284
rect 45928 18300 45980 18352
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 44732 18275 44784 18284
rect 44732 18241 44741 18275
rect 44741 18241 44775 18275
rect 44775 18241 44784 18275
rect 44732 18232 44784 18241
rect 45284 18232 45336 18284
rect 18420 18164 18472 18216
rect 23388 18164 23440 18216
rect 28908 18164 28960 18216
rect 29552 18164 29604 18216
rect 33692 18164 33744 18216
rect 34152 18164 34204 18216
rect 41880 18164 41932 18216
rect 45652 18207 45704 18216
rect 45652 18173 45661 18207
rect 45661 18173 45695 18207
rect 45695 18173 45704 18207
rect 45652 18164 45704 18173
rect 45928 18164 45980 18216
rect 47492 18232 47544 18284
rect 19892 18028 19944 18080
rect 27988 18096 28040 18148
rect 29644 18096 29696 18148
rect 30196 18096 30248 18148
rect 37096 18096 37148 18148
rect 45192 18096 45244 18148
rect 25412 18071 25464 18080
rect 25412 18037 25421 18071
rect 25421 18037 25455 18071
rect 25455 18037 25464 18071
rect 25412 18028 25464 18037
rect 26332 18028 26384 18080
rect 28540 18028 28592 18080
rect 29092 18071 29144 18080
rect 29092 18037 29101 18071
rect 29101 18037 29135 18071
rect 29135 18037 29144 18071
rect 29092 18028 29144 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 22100 17824 22152 17876
rect 24032 17824 24084 17876
rect 44548 17824 44600 17876
rect 20260 17688 20312 17740
rect 23756 17756 23808 17808
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 24768 17620 24820 17672
rect 27712 17756 27764 17808
rect 44732 17756 44784 17808
rect 25780 17688 25832 17740
rect 26240 17688 26292 17740
rect 3516 17552 3568 17604
rect 11060 17552 11112 17604
rect 20168 17595 20220 17604
rect 20168 17561 20177 17595
rect 20177 17561 20211 17595
rect 20211 17561 20220 17595
rect 20168 17552 20220 17561
rect 21916 17552 21968 17604
rect 24676 17595 24728 17604
rect 24676 17561 24685 17595
rect 24685 17561 24719 17595
rect 24719 17561 24728 17595
rect 24676 17552 24728 17561
rect 22192 17484 22244 17536
rect 24400 17484 24452 17536
rect 27896 17688 27948 17740
rect 45376 17731 45428 17740
rect 45376 17697 45385 17731
rect 45385 17697 45419 17731
rect 45419 17697 45428 17731
rect 45376 17688 45428 17697
rect 26976 17620 27028 17672
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 29092 17620 29144 17672
rect 29552 17620 29604 17672
rect 29828 17663 29880 17672
rect 29828 17629 29837 17663
rect 29837 17629 29871 17663
rect 29871 17629 29880 17663
rect 29828 17620 29880 17629
rect 44456 17663 44508 17672
rect 28080 17552 28132 17604
rect 26516 17527 26568 17536
rect 26516 17493 26525 17527
rect 26525 17493 26559 17527
rect 26559 17493 26568 17527
rect 26516 17484 26568 17493
rect 27252 17484 27304 17536
rect 28632 17484 28684 17536
rect 29184 17552 29236 17604
rect 44456 17629 44465 17663
rect 44465 17629 44499 17663
rect 44499 17629 44508 17663
rect 44456 17620 44508 17629
rect 45192 17620 45244 17672
rect 46296 17663 46348 17672
rect 46296 17629 46305 17663
rect 46305 17629 46339 17663
rect 46339 17629 46348 17663
rect 46296 17620 46348 17629
rect 45928 17552 45980 17604
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 33600 17484 33652 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 5448 17212 5500 17264
rect 27804 17280 27856 17332
rect 24308 17212 24360 17264
rect 26516 17212 26568 17264
rect 20996 17144 21048 17196
rect 28632 17280 28684 17332
rect 29000 17280 29052 17332
rect 29828 17280 29880 17332
rect 27988 17144 28040 17196
rect 28540 17144 28592 17196
rect 28816 17187 28868 17196
rect 28816 17153 28825 17187
rect 28825 17153 28859 17187
rect 28859 17153 28868 17187
rect 28816 17144 28868 17153
rect 29092 17144 29144 17196
rect 30104 17280 30156 17332
rect 47676 17323 47728 17332
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 35808 17212 35860 17264
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 22192 17076 22244 17128
rect 13820 17008 13872 17060
rect 25412 17076 25464 17128
rect 29000 17076 29052 17128
rect 30012 17076 30064 17128
rect 33784 17119 33836 17128
rect 33784 17085 33793 17119
rect 33793 17085 33827 17119
rect 33827 17085 33836 17119
rect 33784 17076 33836 17085
rect 35440 17119 35492 17128
rect 35440 17085 35449 17119
rect 35449 17085 35483 17119
rect 35483 17085 35492 17119
rect 35440 17076 35492 17085
rect 29184 17008 29236 17060
rect 46664 17076 46716 17128
rect 46848 17119 46900 17128
rect 46848 17085 46857 17119
rect 46857 17085 46891 17119
rect 46891 17085 46900 17119
rect 46848 17076 46900 17085
rect 46756 17008 46808 17060
rect 1400 16940 1452 16992
rect 24400 16940 24452 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 19984 16600 20036 16652
rect 20996 16600 21048 16652
rect 26332 16736 26384 16788
rect 29552 16779 29604 16788
rect 29552 16745 29561 16779
rect 29561 16745 29595 16779
rect 29595 16745 29604 16779
rect 29552 16736 29604 16745
rect 33784 16779 33836 16788
rect 33784 16745 33793 16779
rect 33793 16745 33827 16779
rect 33827 16745 33836 16779
rect 33784 16736 33836 16745
rect 46296 16736 46348 16788
rect 19432 16532 19484 16584
rect 26240 16643 26292 16652
rect 26240 16609 26249 16643
rect 26249 16609 26283 16643
rect 26283 16609 26292 16643
rect 26240 16600 26292 16609
rect 29184 16600 29236 16652
rect 29644 16600 29696 16652
rect 45652 16668 45704 16720
rect 45468 16643 45520 16652
rect 45468 16609 45477 16643
rect 45477 16609 45511 16643
rect 45511 16609 45520 16643
rect 45468 16600 45520 16609
rect 46940 16600 46992 16652
rect 33692 16575 33744 16584
rect 33692 16541 33701 16575
rect 33701 16541 33735 16575
rect 33735 16541 33744 16575
rect 33692 16532 33744 16541
rect 47308 16575 47360 16584
rect 47308 16541 47317 16575
rect 47317 16541 47351 16575
rect 47351 16541 47360 16575
rect 47308 16532 47360 16541
rect 2136 16464 2188 16516
rect 22008 16507 22060 16516
rect 22008 16473 22017 16507
rect 22017 16473 22051 16507
rect 22051 16473 22060 16507
rect 22008 16464 22060 16473
rect 24400 16507 24452 16516
rect 24400 16473 24409 16507
rect 24409 16473 24443 16507
rect 24443 16473 24452 16507
rect 24400 16464 24452 16473
rect 25780 16464 25832 16516
rect 27252 16464 27304 16516
rect 45192 16507 45244 16516
rect 45192 16473 45201 16507
rect 45201 16473 45235 16507
rect 45235 16473 45244 16507
rect 45192 16464 45244 16473
rect 46664 16464 46716 16516
rect 22928 16396 22980 16448
rect 27712 16439 27764 16448
rect 27712 16405 27721 16439
rect 27721 16405 27755 16439
rect 27755 16405 27764 16439
rect 27712 16396 27764 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 17408 16192 17460 16244
rect 45192 16235 45244 16244
rect 45192 16201 45201 16235
rect 45201 16201 45235 16235
rect 45235 16201 45244 16235
rect 45192 16192 45244 16201
rect 45468 16124 45520 16176
rect 13452 16056 13504 16108
rect 22744 16099 22796 16108
rect 22744 16065 22753 16099
rect 22753 16065 22787 16099
rect 22787 16065 22796 16099
rect 22744 16056 22796 16065
rect 27712 16056 27764 16108
rect 45744 16056 45796 16108
rect 46664 16056 46716 16108
rect 46756 16056 46808 16108
rect 19340 15988 19392 16040
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 22928 15988 22980 15997
rect 29920 16031 29972 16040
rect 29920 15997 29929 16031
rect 29929 15997 29963 16031
rect 29963 15997 29972 16031
rect 29920 15988 29972 15997
rect 31392 16031 31444 16040
rect 31392 15997 31401 16031
rect 31401 15997 31435 16031
rect 31435 15997 31444 16031
rect 31392 15988 31444 15997
rect 45560 15988 45612 16040
rect 2872 15852 2924 15904
rect 17776 15852 17828 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 29920 15691 29972 15700
rect 29920 15657 29929 15691
rect 29929 15657 29963 15691
rect 29963 15657 29972 15691
rect 29920 15648 29972 15657
rect 1768 15444 1820 15496
rect 19340 15444 19392 15496
rect 29828 15487 29880 15496
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 30196 15444 30248 15496
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 19340 14968 19392 15020
rect 2320 14900 2372 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 21732 14764 21784 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 21732 14467 21784 14476
rect 21732 14433 21741 14467
rect 21741 14433 21775 14467
rect 21775 14433 21784 14467
rect 21732 14424 21784 14433
rect 22652 14467 22704 14476
rect 22652 14433 22661 14467
rect 22661 14433 22695 14467
rect 22695 14433 22704 14467
rect 22652 14424 22704 14433
rect 27436 14424 27488 14476
rect 2136 14356 2188 14408
rect 27068 14288 27120 14340
rect 28448 14288 28500 14340
rect 34704 14220 34756 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 29828 13880 29880 13932
rect 46664 13923 46716 13932
rect 46664 13889 46673 13923
rect 46673 13889 46707 13923
rect 46707 13889 46716 13923
rect 46664 13880 46716 13889
rect 8116 13812 8168 13864
rect 3976 13676 4028 13728
rect 10876 13676 10928 13728
rect 46480 13676 46532 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 46480 13379 46532 13388
rect 46480 13345 46489 13379
rect 46489 13345 46523 13379
rect 46523 13345 46532 13379
rect 46480 13336 46532 13345
rect 46296 13311 46348 13320
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 46296 12792 46348 12844
rect 32956 12588 33008 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 47676 11024 47728 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 3148 10956 3200 11008
rect 15568 10956 15620 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 47676 10795 47728 10804
rect 47676 10761 47685 10795
rect 47685 10761 47719 10795
rect 47719 10761 47728 10795
rect 47676 10752 47728 10761
rect 34704 10616 34756 10668
rect 46296 10412 46348 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 46940 9936 46992 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 46940 9639 46992 9648
rect 46940 9605 46949 9639
rect 46949 9605 46983 9639
rect 46983 9605 46992 9639
rect 46940 9596 46992 9605
rect 45652 9528 45704 9580
rect 47308 9528 47360 9580
rect 47860 9571 47912 9580
rect 47860 9537 47869 9571
rect 47869 9537 47903 9571
rect 47903 9537 47912 9571
rect 47860 9528 47912 9537
rect 45836 9392 45888 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47860 8959 47912 8968
rect 47860 8925 47869 8959
rect 47869 8925 47903 8959
rect 47903 8925 47912 8959
rect 47860 8916 47912 8925
rect 32220 8780 32272 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 46112 8483 46164 8492
rect 46112 8449 46121 8483
rect 46121 8449 46155 8483
rect 46155 8449 46164 8483
rect 46112 8440 46164 8449
rect 2044 8304 2096 8356
rect 39120 8236 39172 8288
rect 45744 8236 45796 8288
rect 46388 8236 46440 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 45928 7896 45980 7948
rect 46388 7871 46440 7880
rect 46388 7837 46397 7871
rect 46397 7837 46431 7871
rect 46431 7837 46440 7871
rect 46388 7828 46440 7837
rect 46940 7803 46992 7812
rect 46940 7769 46949 7803
rect 46949 7769 46983 7803
rect 46983 7769 46992 7803
rect 46940 7760 46992 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 46940 7488 46992 7540
rect 46112 7463 46164 7472
rect 46112 7429 46121 7463
rect 46121 7429 46155 7463
rect 46155 7429 46164 7463
rect 46112 7420 46164 7429
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 46020 7327 46072 7336
rect 46020 7293 46029 7327
rect 46029 7293 46063 7327
rect 46063 7293 46072 7327
rect 46020 7284 46072 7293
rect 45928 7216 45980 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3424 6808 3476 6860
rect 28356 6808 28408 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47216 6740 47268 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 48044 6443 48096 6452
rect 48044 6409 48053 6443
rect 48053 6409 48087 6443
rect 48087 6409 48096 6443
rect 48044 6400 48096 6409
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 40132 5652 40184 5704
rect 40040 5516 40092 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3976 5244 4028 5296
rect 37280 5312 37332 5364
rect 37372 5312 37424 5364
rect 37556 5244 37608 5296
rect 20260 5176 20312 5228
rect 23020 5176 23072 5228
rect 23480 5219 23532 5228
rect 23480 5185 23489 5219
rect 23489 5185 23523 5219
rect 23523 5185 23532 5219
rect 23480 5176 23532 5185
rect 37372 5151 37424 5160
rect 37372 5117 37381 5151
rect 37381 5117 37415 5151
rect 37415 5117 37424 5151
rect 37372 5108 37424 5117
rect 38292 5151 38344 5160
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 23756 5040 23808 5092
rect 30104 5040 30156 5092
rect 42340 5244 42392 5296
rect 40040 5219 40092 5228
rect 40040 5185 40049 5219
rect 40049 5185 40083 5219
rect 40083 5185 40092 5219
rect 40040 5176 40092 5185
rect 40224 5151 40276 5160
rect 40224 5117 40233 5151
rect 40233 5117 40267 5151
rect 40267 5117 40276 5151
rect 40224 5108 40276 5117
rect 41880 5151 41932 5160
rect 41880 5117 41889 5151
rect 41889 5117 41923 5151
rect 41923 5117 41932 5151
rect 41880 5108 41932 5117
rect 20076 4972 20128 5024
rect 24768 4972 24820 5024
rect 37372 4972 37424 5024
rect 46756 5176 46808 5228
rect 43720 5108 43772 5160
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 40224 4811 40276 4820
rect 40224 4777 40233 4811
rect 40233 4777 40267 4811
rect 40267 4777 40276 4811
rect 40224 4768 40276 4777
rect 42340 4811 42392 4820
rect 42340 4777 42349 4811
rect 42349 4777 42383 4811
rect 42383 4777 42392 4811
rect 42340 4768 42392 4777
rect 40132 4700 40184 4752
rect 46112 4700 46164 4752
rect 21272 4632 21324 4684
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 22560 4564 22612 4616
rect 23204 4564 23256 4616
rect 40408 4607 40460 4616
rect 22192 4496 22244 4548
rect 40408 4573 40417 4607
rect 40417 4573 40451 4607
rect 40451 4573 40460 4607
rect 40408 4564 40460 4573
rect 40776 4564 40828 4616
rect 42892 4564 42944 4616
rect 47492 4632 47544 4684
rect 46848 4564 46900 4616
rect 19432 4471 19484 4480
rect 19432 4437 19441 4471
rect 19441 4437 19475 4471
rect 19475 4437 19484 4471
rect 19432 4428 19484 4437
rect 20628 4428 20680 4480
rect 21088 4471 21140 4480
rect 21088 4437 21097 4471
rect 21097 4437 21131 4471
rect 21131 4437 21140 4471
rect 21088 4428 21140 4437
rect 22284 4428 22336 4480
rect 22468 4428 22520 4480
rect 23296 4428 23348 4480
rect 46480 4428 46532 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 3424 4020 3476 4072
rect 17868 4088 17920 4140
rect 18328 4088 18380 4140
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19800 4156 19852 4208
rect 20996 4224 21048 4276
rect 21640 4224 21692 4276
rect 22560 4267 22612 4276
rect 22560 4233 22569 4267
rect 22569 4233 22603 4267
rect 22603 4233 22612 4267
rect 22560 4224 22612 4233
rect 37556 4224 37608 4276
rect 40408 4224 40460 4276
rect 22376 4156 22428 4208
rect 25596 4156 25648 4208
rect 40776 4156 40828 4208
rect 43260 4156 43312 4208
rect 43720 4199 43772 4208
rect 43720 4165 43729 4199
rect 43729 4165 43763 4199
rect 43763 4165 43772 4199
rect 43720 4156 43772 4165
rect 46664 4199 46716 4208
rect 46664 4165 46673 4199
rect 46673 4165 46707 4199
rect 46707 4165 46716 4199
rect 46664 4156 46716 4165
rect 47860 4156 47912 4208
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 21088 4088 21140 4140
rect 22284 4088 22336 4140
rect 22560 4088 22612 4140
rect 23388 4088 23440 4140
rect 20904 4020 20956 4072
rect 24400 4020 24452 4072
rect 25228 4088 25280 4140
rect 28816 4088 28868 4140
rect 30932 4088 30984 4140
rect 37740 4088 37792 4140
rect 40500 4131 40552 4140
rect 24676 3952 24728 4004
rect 26608 4020 26660 4072
rect 28540 4020 28592 4072
rect 39396 4063 39448 4072
rect 39396 4029 39405 4063
rect 39405 4029 39439 4063
rect 39439 4029 39448 4063
rect 39396 4020 39448 4029
rect 39580 4063 39632 4072
rect 39580 4029 39589 4063
rect 39589 4029 39623 4063
rect 39623 4029 39632 4063
rect 39580 4020 39632 4029
rect 40224 4020 40276 4072
rect 40500 4097 40509 4131
rect 40509 4097 40543 4131
rect 40543 4097 40552 4131
rect 40500 4088 40552 4097
rect 40776 4020 40828 4072
rect 46020 4088 46072 4140
rect 43720 4020 43772 4072
rect 1952 3884 2004 3936
rect 2780 3884 2832 3936
rect 6552 3884 6604 3936
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 7932 3884 7984 3936
rect 9312 3884 9364 3936
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 11520 3884 11572 3936
rect 17592 3884 17644 3936
rect 18880 3884 18932 3936
rect 23112 3884 23164 3936
rect 23848 3927 23900 3936
rect 23848 3893 23857 3927
rect 23857 3893 23891 3927
rect 23891 3893 23900 3927
rect 23848 3884 23900 3893
rect 24584 3884 24636 3936
rect 25320 3884 25372 3936
rect 30380 3884 30432 3936
rect 40316 3884 40368 3936
rect 43536 3884 43588 3936
rect 46296 3884 46348 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19248 3680 19300 3732
rect 20352 3680 20404 3732
rect 3884 3612 3936 3664
rect 35532 3680 35584 3732
rect 22560 3655 22612 3664
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 23204 3655 23256 3664
rect 23204 3621 23213 3655
rect 23213 3621 23247 3655
rect 23247 3621 23256 3655
rect 23204 3612 23256 3621
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 10140 3544 10192 3596
rect 1768 3476 1820 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 1308 3408 1360 3460
rect 6736 3451 6788 3460
rect 6736 3417 6745 3451
rect 6745 3417 6779 3451
rect 6779 3417 6788 3451
rect 6736 3408 6788 3417
rect 9036 3408 9088 3460
rect 20444 3544 20496 3596
rect 20812 3544 20864 3596
rect 30380 3612 30432 3664
rect 24768 3544 24820 3596
rect 26608 3587 26660 3596
rect 26608 3553 26617 3587
rect 26617 3553 26651 3587
rect 26651 3553 26660 3587
rect 26608 3544 26660 3553
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 13820 3476 13872 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 17776 3476 17828 3528
rect 19800 3476 19852 3528
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 26700 3476 26752 3528
rect 27344 3476 27396 3528
rect 35440 3544 35492 3596
rect 37280 3544 37332 3596
rect 39396 3612 39448 3664
rect 40500 3680 40552 3732
rect 44272 3612 44324 3664
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 33784 3519 33836 3528
rect 33784 3485 33793 3519
rect 33793 3485 33827 3519
rect 33827 3485 33836 3519
rect 33784 3476 33836 3485
rect 20352 3451 20404 3460
rect 11704 3340 11756 3392
rect 14004 3340 14056 3392
rect 18236 3340 18288 3392
rect 20352 3417 20361 3451
rect 20361 3417 20395 3451
rect 20395 3417 20404 3451
rect 20352 3408 20404 3417
rect 20904 3340 20956 3392
rect 21916 3340 21968 3392
rect 24492 3340 24544 3392
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 30012 3408 30064 3460
rect 38292 3587 38344 3596
rect 38292 3553 38301 3587
rect 38301 3553 38335 3587
rect 38335 3553 38344 3587
rect 38292 3544 38344 3553
rect 41696 3544 41748 3596
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 42800 3544 42852 3596
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 39120 3476 39172 3528
rect 39580 3476 39632 3528
rect 40960 3519 41012 3528
rect 40960 3485 40969 3519
rect 40969 3485 41003 3519
rect 41003 3485 41012 3519
rect 40960 3476 41012 3485
rect 42708 3476 42760 3528
rect 45192 3519 45244 3528
rect 38660 3408 38712 3460
rect 39764 3408 39816 3460
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 45652 3519 45704 3528
rect 45652 3485 45661 3519
rect 45661 3485 45695 3519
rect 45695 3485 45704 3519
rect 45652 3476 45704 3485
rect 46204 3408 46256 3460
rect 48964 3408 49016 3460
rect 33140 3340 33192 3392
rect 39948 3340 40000 3392
rect 42984 3340 43036 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 6736 3179 6788 3188
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 14096 3136 14148 3188
rect 18328 3179 18380 3188
rect 18328 3145 18337 3179
rect 18337 3145 18371 3179
rect 18371 3145 18380 3179
rect 18328 3136 18380 3145
rect 19340 3136 19392 3188
rect 20352 3136 20404 3188
rect 24400 3136 24452 3188
rect 24492 3136 24544 3188
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 7932 3043 7984 3052
rect 6644 3000 6696 3009
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 18696 3068 18748 3120
rect 23388 3068 23440 3120
rect 24768 3111 24820 3120
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 24860 3068 24912 3120
rect 25228 3068 25280 3120
rect 30012 3068 30064 3120
rect 32220 3068 32272 3120
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 664 2932 716 2984
rect 7748 2932 7800 2984
rect 10968 2932 11020 2984
rect 14188 2932 14240 2984
rect 15200 2932 15252 2984
rect 17776 2975 17828 2984
rect 17776 2941 17785 2975
rect 17785 2941 17819 2975
rect 17819 2941 17828 2975
rect 17776 2932 17828 2941
rect 20168 3000 20220 3052
rect 22192 3000 22244 3052
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 23296 3000 23348 3052
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 27068 3000 27120 3052
rect 33784 3136 33836 3188
rect 37740 3179 37792 3188
rect 37740 3145 37749 3179
rect 37749 3145 37783 3179
rect 37783 3145 37792 3179
rect 37740 3136 37792 3145
rect 39764 3179 39816 3188
rect 39764 3145 39773 3179
rect 39773 3145 39807 3179
rect 39807 3145 39816 3179
rect 39764 3136 39816 3145
rect 40960 3136 41012 3188
rect 47768 3136 47820 3188
rect 33140 3111 33192 3120
rect 33140 3077 33149 3111
rect 33149 3077 33183 3111
rect 33183 3077 33192 3111
rect 33140 3068 33192 3077
rect 22008 2932 22060 2984
rect 24860 2932 24912 2984
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 12072 2864 12124 2916
rect 13360 2796 13412 2848
rect 18696 2796 18748 2848
rect 21272 2796 21324 2848
rect 23572 2796 23624 2848
rect 31300 2796 31352 2848
rect 32956 2796 33008 2848
rect 42708 3068 42760 3120
rect 42984 3111 43036 3120
rect 42984 3077 42993 3111
rect 42993 3077 43027 3111
rect 43027 3077 43036 3111
rect 42984 3068 43036 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 38660 3000 38712 3052
rect 39948 3043 40000 3052
rect 39948 3009 39957 3043
rect 39957 3009 39991 3043
rect 39991 3009 40000 3043
rect 39948 3000 40000 3009
rect 39396 2932 39448 2984
rect 40776 3000 40828 3052
rect 42800 3043 42852 3052
rect 42800 3009 42809 3043
rect 42809 3009 42843 3043
rect 42843 3009 42852 3043
rect 42800 3000 42852 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 48320 3000 48372 3052
rect 41696 2932 41748 2984
rect 43168 2932 43220 2984
rect 47676 2932 47728 2984
rect 37280 2864 37332 2916
rect 45100 2864 45152 2916
rect 37372 2839 37424 2848
rect 37372 2805 37381 2839
rect 37381 2805 37415 2839
rect 37415 2805 37424 2839
rect 37372 2796 37424 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20536 2592 20588 2644
rect 22376 2635 22428 2644
rect 22376 2601 22385 2635
rect 22385 2601 22419 2635
rect 22419 2601 22428 2635
rect 22376 2592 22428 2601
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 28080 2592 28132 2644
rect 28172 2592 28224 2644
rect 30288 2592 30340 2644
rect 3976 2524 4028 2576
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 15200 2524 15252 2576
rect 20260 2524 20312 2576
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 5172 2388 5224 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 16120 2388 16172 2440
rect 19432 2388 19484 2440
rect 20076 2388 20128 2440
rect 20628 2388 20680 2440
rect 21180 2388 21232 2440
rect 23848 2456 23900 2508
rect 26700 2524 26752 2576
rect 35624 2592 35676 2644
rect 39120 2635 39172 2644
rect 39120 2601 39129 2635
rect 39129 2601 39163 2635
rect 39163 2601 39172 2635
rect 39120 2592 39172 2601
rect 41696 2635 41748 2644
rect 41696 2601 41705 2635
rect 41705 2601 41739 2635
rect 41739 2601 41748 2635
rect 41696 2592 41748 2601
rect 42524 2635 42576 2644
rect 42524 2601 42533 2635
rect 42533 2601 42567 2635
rect 42567 2601 42576 2635
rect 42524 2592 42576 2601
rect 42892 2635 42944 2644
rect 42892 2601 42901 2635
rect 42901 2601 42935 2635
rect 42935 2601 42944 2635
rect 42892 2592 42944 2601
rect 43076 2524 43128 2576
rect 2780 2320 2832 2372
rect 2596 2252 2648 2304
rect 7564 2320 7616 2372
rect 8392 2320 8444 2372
rect 15476 2320 15528 2372
rect 21916 2320 21968 2372
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 25504 2388 25556 2440
rect 26424 2388 26476 2440
rect 27988 2456 28040 2508
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 6460 2252 6512 2304
rect 7012 2252 7064 2304
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 22008 2252 22060 2304
rect 24492 2320 24544 2372
rect 28080 2320 28132 2372
rect 31208 2456 31260 2508
rect 35440 2388 35492 2440
rect 37372 2388 37424 2440
rect 38016 2388 38068 2440
rect 39948 2388 40000 2440
rect 41236 2388 41288 2440
rect 43260 2456 43312 2508
rect 47400 2456 47452 2508
rect 43812 2388 43864 2440
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 36084 2320 36136 2372
rect 39396 2320 39448 2372
rect 40592 2320 40644 2372
rect 38660 2252 38712 2304
rect 47032 2388 47084 2440
rect 48044 2388 48096 2440
rect 46388 2320 46440 2372
rect 45468 2295 45520 2304
rect 45468 2261 45477 2295
rect 45477 2261 45511 2295
rect 45511 2261 45520 2295
rect 45468 2252 45520 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 9680 2048 9732 2100
rect 23940 2048 23992 2100
rect 4436 1980 4488 2032
rect 29552 1980 29604 2032
rect 3516 1912 3568 1964
rect 16856 1912 16908 1964
rect 26792 1912 26844 1964
rect 28724 1912 28776 1964
rect 45468 1912 45520 1964
rect 28448 1844 28500 1896
rect 29736 1844 29788 1896
rect 42524 1844 42576 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4844 49314
rect 4498 49200 4610 49286
rect 32 26450 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 1964 47054 1992 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2504 46980 2556 46986
rect 2504 46922 2556 46928
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2412 46368 2464 46374
rect 2412 46310 2464 46316
rect 2228 45892 2280 45898
rect 2228 45834 2280 45840
rect 2240 45626 2268 45834
rect 2228 45620 2280 45626
rect 2228 45562 2280 45568
rect 1952 45484 2004 45490
rect 1952 45426 2004 45432
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 20 26444 72 26450
rect 20 26386 72 26392
rect 1504 26234 1532 43182
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1584 41540 1636 41546
rect 1858 41511 1914 41520
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1964 35894 1992 45426
rect 2044 40452 2096 40458
rect 2044 40394 2096 40400
rect 2056 36310 2084 40394
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2044 36304 2096 36310
rect 2044 36246 2096 36252
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 1964 35866 2084 35894
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35465 1624 35634
rect 1860 35488 1912 35494
rect 1582 35456 1638 35465
rect 1860 35430 1912 35436
rect 1582 35391 1638 35400
rect 1584 33992 1636 33998
rect 1584 33934 1636 33940
rect 1596 32745 1624 33934
rect 1676 33448 1728 33454
rect 1676 33390 1728 33396
rect 1688 32910 1716 33390
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1872 32434 1900 35430
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1964 33114 1992 33798
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1860 32428 1912 32434
rect 1860 32370 1912 32376
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1964 31958 1992 32846
rect 1952 31952 2004 31958
rect 1952 31894 2004 31900
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 2056 31346 2084 35866
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1504 26206 1624 26234
rect 1596 18426 1624 26206
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 12345 1900 12786
rect 1858 12336 1914 12345
rect 1858 12271 1914 12280
rect 2056 8362 2084 25094
rect 2148 18902 2176 36110
rect 2228 32768 2280 32774
rect 2228 32710 2280 32716
rect 2240 32502 2268 32710
rect 2228 32496 2280 32502
rect 2228 32438 2280 32444
rect 2332 27577 2360 46310
rect 2424 46034 2452 46310
rect 2412 46028 2464 46034
rect 2412 45970 2464 45976
rect 2516 45554 2544 46922
rect 2608 46918 2636 49200
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 3422 46951 3478 46960
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 2872 46912 2924 46918
rect 2872 46854 2924 46860
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2792 46034 2820 46271
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2424 45526 2544 45554
rect 2318 27568 2374 27577
rect 2318 27503 2374 27512
rect 2424 22545 2452 45526
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2410 22536 2466 22545
rect 2410 22471 2466 22480
rect 2884 21486 2912 46854
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 3436 20602 3464 46951
rect 3896 46646 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4816 47054 4844 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7420 49314
rect 7074 49200 7186 49286
rect 5828 47054 5856 49200
rect 7392 47054 7420 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7380 47048 7432 47054
rect 7380 46990 7432 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 7472 46980 7524 46986
rect 7472 46922 7524 46928
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3514 44976 3570 44985
rect 3514 44911 3570 44920
rect 3528 21078 3556 44911
rect 3698 43616 3754 43625
rect 3698 43551 3754 43560
rect 3712 31770 3740 43551
rect 3882 39536 3938 39545
rect 3882 39471 3938 39480
rect 3792 32564 3844 32570
rect 3792 32506 3844 32512
rect 3804 31890 3832 32506
rect 3896 32026 3924 39471
rect 3884 32020 3936 32026
rect 3884 31962 3936 31968
rect 3792 31884 3844 31890
rect 3792 31826 3844 31832
rect 3712 31742 3832 31770
rect 3804 28694 3832 31742
rect 3882 31376 3938 31385
rect 3882 31311 3938 31320
rect 3792 28688 3844 28694
rect 3792 28630 3844 28636
rect 3896 24138 3924 31311
rect 3974 28656 4030 28665
rect 3974 28591 3976 28600
rect 4028 28591 4030 28600
rect 3976 28562 4028 28568
rect 3884 24132 3936 24138
rect 3884 24074 3936 24080
rect 3516 21072 3568 21078
rect 3516 21014 3568 21020
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3988 19825 4016 20266
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 3976 19236 4028 19242
rect 3976 19178 4028 19184
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2148 18766 2176 18838
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 3988 18465 4016 19178
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3332 18352 3384 18358
rect 3332 18294 3384 18300
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2332 14618 2360 14894
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2148 4146 2176 14350
rect 2884 6914 2912 15846
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10305 3188 10950
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 3344 7585 3372 18294
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3528 17105 3556 17546
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3976 13728 4028 13734
rect 3974 13696 3976 13705
rect 4028 13696 4030 13705
rect 3974 13631 4030 13640
rect 3330 7576 3386 7585
rect 3330 7511 3386 7520
rect 4080 6914 4108 46922
rect 4896 46912 4948 46918
rect 4896 46854 4948 46860
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4632 31890 4660 32302
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4908 19446 4936 46854
rect 7484 32230 7512 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 8312 31958 8340 45526
rect 9508 34134 9536 46922
rect 10980 46374 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 12912 47054 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 13740 47110 13860 47138
rect 13832 47054 13860 47110
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 13820 47048 13872 47054
rect 13820 46990 13872 46996
rect 11704 46980 11756 46986
rect 11704 46922 11756 46928
rect 12440 46980 12492 46986
rect 12440 46922 12492 46928
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 11716 38010 11744 46922
rect 12072 46504 12124 46510
rect 12072 46446 12124 46452
rect 12084 46170 12112 46446
rect 12072 46164 12124 46170
rect 12072 46106 12124 46112
rect 11980 45960 12032 45966
rect 11980 45902 12032 45908
rect 11992 45626 12020 45902
rect 11980 45620 12032 45626
rect 11980 45562 12032 45568
rect 11704 38004 11756 38010
rect 11704 37946 11756 37952
rect 12452 36650 12480 46922
rect 14200 46594 14228 49200
rect 14372 47048 14424 47054
rect 14372 46990 14424 46996
rect 14200 46566 14320 46594
rect 14292 46510 14320 46566
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 13556 46170 13584 46446
rect 14200 46170 14228 46446
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 12440 36644 12492 36650
rect 12440 36586 12492 36592
rect 9496 34128 9548 34134
rect 9496 34070 9548 34076
rect 14384 33522 14412 46990
rect 15488 45554 15516 49200
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49314 17490 50000
rect 17378 49286 17908 49314
rect 17378 49200 17490 49286
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 17776 47048 17828 47054
rect 17776 46990 17828 46996
rect 15488 45526 15884 45554
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 8300 31952 8352 31958
rect 8300 31894 8352 31900
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 5460 17270 5488 31826
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9220 30184 9272 30190
rect 9220 30126 9272 30132
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8496 28082 8524 29106
rect 9232 28082 9260 30126
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9692 29714 9720 29990
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9324 29306 9352 29582
rect 9784 29306 9812 30194
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10336 29578 10364 29990
rect 11716 29714 11744 31758
rect 12900 31748 12952 31754
rect 12900 31690 12952 31696
rect 15016 31748 15068 31754
rect 15016 31690 15068 31696
rect 12912 31482 12940 31690
rect 15028 31482 15056 31690
rect 12900 31476 12952 31482
rect 12900 31418 12952 31424
rect 15016 31476 15068 31482
rect 15016 31418 15068 31424
rect 14740 31340 14792 31346
rect 14740 31282 14792 31288
rect 12532 30728 12584 30734
rect 12532 30670 12584 30676
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 12440 30592 12492 30598
rect 12440 30534 12492 30540
rect 12452 30326 12480 30534
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 11888 29776 11940 29782
rect 11888 29718 11940 29724
rect 11704 29708 11756 29714
rect 11704 29650 11756 29656
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8312 27538 8340 27814
rect 8300 27532 8352 27538
rect 8300 27474 8352 27480
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8404 27130 8432 27406
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8496 26382 8524 28018
rect 9232 26994 9260 28018
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 27402 9720 27814
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9312 26920 9364 26926
rect 9312 26862 9364 26868
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 7932 26240 7984 26246
rect 7932 26182 7984 26188
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 7944 25906 7972 26182
rect 8312 25974 8340 26182
rect 8772 25974 8800 26726
rect 9324 26450 9352 26862
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8760 25968 8812 25974
rect 8760 25910 8812 25916
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 9140 24206 9168 26318
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9692 25770 9720 26182
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23186 9076 24006
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9600 22778 9628 22986
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 9588 21344 9640 21350
rect 9692 21332 9720 24074
rect 9784 23866 9812 28018
rect 9968 26382 9996 29038
rect 11256 29034 11284 29446
rect 11716 29238 11744 29650
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11900 29170 11928 29718
rect 12084 29170 12112 29786
rect 12164 29640 12216 29646
rect 12544 29594 12572 30670
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 13096 30326 13124 30534
rect 13084 30320 13136 30326
rect 13084 30262 13136 30268
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12164 29582 12216 29588
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11900 28914 11928 29106
rect 12176 29102 12204 29582
rect 12452 29566 12572 29594
rect 12452 29306 12480 29566
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 11900 28886 12020 28914
rect 10048 28484 10100 28490
rect 10048 28426 10100 28432
rect 10060 28218 10088 28426
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10428 27062 10456 28358
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 11900 27334 11928 28018
rect 11992 28014 12020 28886
rect 12176 28082 12204 29038
rect 12636 28762 12664 29990
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 13004 29238 13032 29514
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 13096 29306 13124 29446
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 12992 29232 13044 29238
rect 12992 29174 13044 29180
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12176 27674 12204 27814
rect 12164 27668 12216 27674
rect 12164 27610 12216 27616
rect 12728 27538 12756 27814
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10416 27056 10468 27062
rect 10416 26998 10468 27004
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10336 26518 10364 26930
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9876 26042 9904 26250
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 10428 25362 10456 26998
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10520 25702 10548 26318
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10520 25498 10548 25638
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10612 25362 10640 26930
rect 10796 26330 10824 27066
rect 11348 26994 11376 27270
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11060 26354 11112 26360
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10796 26302 11060 26330
rect 10704 25974 10732 26250
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10796 25770 10824 26302
rect 11060 26296 11112 26302
rect 10784 25764 10836 25770
rect 10784 25706 10836 25712
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 24342 10088 25094
rect 10048 24336 10100 24342
rect 10048 24278 10100 24284
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 10152 22642 10180 24006
rect 10428 23322 10456 25298
rect 10796 25158 10824 25706
rect 11256 25362 11284 26862
rect 11348 25906 11376 26930
rect 11612 26920 11664 26926
rect 11532 26880 11612 26908
rect 11532 26382 11560 26880
rect 11612 26862 11664 26868
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11440 25362 11468 26182
rect 11532 25974 11560 26318
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11624 25702 11652 26250
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11612 25696 11664 25702
rect 11612 25638 11664 25644
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10704 23050 10732 24006
rect 10692 23044 10744 23050
rect 10692 22986 10744 22992
rect 10796 22642 10824 25094
rect 11716 23730 11744 25842
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9968 21690 9996 21898
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 9640 21304 9720 21332
rect 9588 21286 9640 21292
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 20466 9168 20878
rect 9324 20534 9352 21286
rect 9600 21010 9628 21286
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 10140 21004 10192 21010
rect 10140 20946 10192 20952
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9140 20058 9168 20402
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 10152 19922 10180 20946
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 19514 9904 19790
rect 10428 19718 10456 21490
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 10428 19378 10456 19654
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 2792 6886 2912 6914
rect 3422 6896 3478 6905
rect 2792 4146 2820 6886
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3988 6886 4108 6914
rect 3424 6802 3476 6808
rect 3988 5302 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3402
rect 1780 3058 1808 3470
rect 1964 3126 1992 3878
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2792 2378 2820 3878
rect 3436 3505 3464 4014
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 3528 1465 3556 1906
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3896 800 3924 3606
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 2582 4016 3470
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 6564 2446 6592 3878
rect 6656 3058 6684 18906
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6748 3194 6776 3402
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4448 2038 4476 2246
rect 4436 2032 4488 2038
rect 4436 1974 4488 1980
rect 5184 800 5212 2382
rect 7024 2310 7052 2450
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6472 800 6500 2246
rect 7116 800 7144 3538
rect 7576 2378 7604 3878
rect 7944 3058 7972 3878
rect 8128 3126 8156 13806
rect 10888 13734 10916 23598
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 22506 11376 23054
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11716 22710 11744 22918
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 11072 17610 11100 21898
rect 11348 21622 11376 22442
rect 11900 22098 11928 27270
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12084 24886 12112 25094
rect 12072 24880 12124 24886
rect 12072 24822 12124 24828
rect 12452 24342 12480 25230
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24750 12572 25094
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12636 24562 12664 25230
rect 13372 25226 13400 29038
rect 13464 28082 13492 30670
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13464 27130 13492 28018
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13556 27402 13584 27814
rect 13544 27396 13596 27402
rect 13544 27338 13596 27344
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 26790 13860 26930
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13372 24954 13400 25162
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 12544 24534 12664 24562
rect 12440 24336 12492 24342
rect 12440 24278 12492 24284
rect 12544 24206 12572 24534
rect 13188 24410 13216 24754
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 12544 22030 12572 24142
rect 13096 23322 13124 24210
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13096 22166 13124 23258
rect 13832 23118 13860 26726
rect 14108 26234 14136 30262
rect 14200 28558 14228 30670
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14292 29646 14320 30194
rect 14384 29646 14412 30330
rect 14752 30326 14780 31282
rect 15016 30660 15068 30666
rect 15016 30602 15068 30608
rect 14740 30320 14792 30326
rect 14740 30262 14792 30268
rect 15028 29714 15056 30602
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14292 29306 14320 29582
rect 14384 29306 14412 29582
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14200 28014 14228 28494
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 14188 28008 14240 28014
rect 14188 27950 14240 27956
rect 14200 27470 14228 27950
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14556 27396 14608 27402
rect 14556 27338 14608 27344
rect 14568 26234 14596 27338
rect 14660 26790 14688 28358
rect 15212 27538 15240 31826
rect 15476 30116 15528 30122
rect 15476 30058 15528 30064
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15396 29714 15424 29990
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15488 29578 15516 30058
rect 15856 30054 15884 45526
rect 17500 37800 17552 37806
rect 17500 37742 17552 37748
rect 17512 35834 17540 37742
rect 17500 35828 17552 35834
rect 17500 35770 17552 35776
rect 16672 35556 16724 35562
rect 16672 35498 16724 35504
rect 16684 35086 16712 35498
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16960 35086 16988 35430
rect 16672 35080 16724 35086
rect 16672 35022 16724 35028
rect 16948 35080 17000 35086
rect 16948 35022 17000 35028
rect 17512 34610 17540 35770
rect 17788 35086 17816 46990
rect 17592 35080 17644 35086
rect 17592 35022 17644 35028
rect 17776 35080 17828 35086
rect 17776 35022 17828 35028
rect 17604 34746 17632 35022
rect 17592 34740 17644 34746
rect 17644 34700 17816 34728
rect 17592 34682 17644 34688
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17696 31890 17724 32166
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17788 31822 17816 34700
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 17880 30802 17908 49286
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49314 20710 50000
rect 20456 49286 20710 49314
rect 18708 46918 18736 49200
rect 19996 46918 20024 49200
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 20456 46510 20484 49286
rect 20598 49200 20710 49286
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26712 49286 27150 49314
rect 20536 47184 20588 47190
rect 20536 47126 20588 47132
rect 19248 46504 19300 46510
rect 19248 46446 19300 46452
rect 20444 46504 20496 46510
rect 20444 46446 20496 46452
rect 18604 46436 18656 46442
rect 18604 46378 18656 46384
rect 18616 46170 18644 46378
rect 19260 46170 19288 46446
rect 18604 46164 18656 46170
rect 18604 46106 18656 46112
rect 19248 46164 19300 46170
rect 19248 46106 19300 46112
rect 18696 45960 18748 45966
rect 18696 45902 18748 45908
rect 18708 41414 18736 45902
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 18708 41386 18828 41414
rect 18144 39432 18196 39438
rect 18144 39374 18196 39380
rect 18156 37942 18184 39374
rect 18512 38344 18564 38350
rect 18512 38286 18564 38292
rect 18144 37936 18196 37942
rect 18144 37878 18196 37884
rect 18236 37800 18288 37806
rect 18236 37742 18288 37748
rect 18248 37466 18276 37742
rect 18236 37460 18288 37466
rect 18236 37402 18288 37408
rect 18524 36174 18552 38286
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 35222 18000 35634
rect 17960 35216 18012 35222
rect 17960 35158 18012 35164
rect 18236 35080 18288 35086
rect 18236 35022 18288 35028
rect 18052 34944 18104 34950
rect 18052 34886 18104 34892
rect 18064 34678 18092 34886
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18248 32978 18276 35022
rect 18524 34678 18552 35974
rect 18512 34672 18564 34678
rect 18512 34614 18564 34620
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 18156 32502 18184 32710
rect 18144 32496 18196 32502
rect 18144 32438 18196 32444
rect 18248 31822 18276 32914
rect 18236 31816 18288 31822
rect 18236 31758 18288 31764
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 18340 31278 18368 31622
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 17868 30796 17920 30802
rect 17868 30738 17920 30744
rect 16304 30728 16356 30734
rect 16304 30670 16356 30676
rect 16316 30394 16344 30670
rect 16580 30660 16632 30666
rect 16580 30602 16632 30608
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15476 29572 15528 29578
rect 15476 29514 15528 29520
rect 15488 28762 15516 29514
rect 15764 29238 15792 29990
rect 16592 29306 16620 30602
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 16684 29850 16712 30126
rect 17512 29850 17540 30126
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 15476 28756 15528 28762
rect 15476 28698 15528 28704
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15212 27130 15240 27338
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 15304 26518 15332 28018
rect 15488 26994 15516 28698
rect 16040 28082 16068 29106
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16120 28484 16172 28490
rect 16120 28426 16172 28432
rect 16132 28218 16160 28426
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15856 27334 15884 27474
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15856 26994 15884 27270
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 15488 26450 15516 26522
rect 15844 26512 15896 26518
rect 15844 26454 15896 26460
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 14108 26206 14228 26234
rect 14568 26206 14688 26234
rect 14200 24750 14228 26206
rect 14660 25906 14688 26206
rect 15764 25974 15792 26318
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14660 25498 14688 25842
rect 15384 25832 15436 25838
rect 15384 25774 15436 25780
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 15028 25362 15056 25638
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15304 24954 15332 25162
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14292 24274 14320 24550
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14016 23662 14044 24074
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 14004 23656 14056 23662
rect 14004 23598 14056 23604
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 11336 21616 11388 21622
rect 11336 21558 11388 21564
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11900 21146 11928 21422
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11992 20874 12020 21422
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11992 20534 12020 20810
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 12268 20262 12296 20742
rect 12452 20466 12480 21966
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12544 21622 12572 21830
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 20942 12572 21286
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12544 20534 12572 20878
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12728 20602 12756 20810
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11440 19786 11468 20198
rect 12268 20058 12296 20198
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12268 19854 12296 19994
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 18834 11744 19654
rect 12452 19446 12480 20402
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12728 19310 12756 20538
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 11992 18834 12020 19110
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 13096 18766 13124 19110
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 9324 3602 9352 3878
rect 10152 3602 10180 3878
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7760 800 7788 2926
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 3402
rect 11532 3058 11560 3878
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3126 11744 3334
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2106 9720 2246
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 10980 800 11008 2926
rect 12084 2922 12112 3470
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 13372 2854 13400 22510
rect 13648 20466 13676 22918
rect 13924 22778 13952 23598
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13832 19786 13860 21830
rect 14292 21554 14320 21830
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14568 21078 14596 21422
rect 14752 21350 14780 24074
rect 14936 23186 14964 24754
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 23730 15148 24550
rect 15396 24342 15424 25774
rect 15856 24818 15884 26454
rect 16132 26042 16160 26862
rect 16408 26382 16436 28562
rect 16776 28218 16804 29514
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 17972 28218 18000 28970
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17052 27470 17080 28018
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16408 26042 16436 26318
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16132 24818 16160 25978
rect 16408 25786 16436 25978
rect 16684 25906 16712 26318
rect 16776 25974 16804 27270
rect 17052 27062 17080 27406
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 17052 25906 17080 26182
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16408 25758 16528 25786
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16408 25294 16436 25638
rect 16500 25498 16528 25758
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16684 25362 16712 25842
rect 17052 25770 17080 25842
rect 17040 25764 17092 25770
rect 17040 25706 17092 25712
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 17052 25294 17080 25706
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15108 23724 15160 23730
rect 15108 23666 15160 23672
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 14936 22642 14964 23122
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15120 22642 15148 23054
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15396 22506 15424 23734
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15212 22030 15240 22442
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14556 21072 14608 21078
rect 14556 21014 14608 21020
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 20262 14412 20810
rect 14476 20602 14504 20878
rect 14752 20602 14780 21286
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 19310 13492 19654
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13464 18630 13492 19246
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 16114 13492 18566
rect 13832 18290 13860 19722
rect 14384 19310 14412 20198
rect 14568 19718 14596 20334
rect 14752 19786 14780 20538
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14844 19854 14872 20334
rect 15028 20058 15056 20402
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15212 19990 15240 20266
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 18834 14780 19110
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14108 18426 14136 18702
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16574 13860 17002
rect 13832 16546 14872 16574
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13832 3058 13860 3470
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 3126 14044 3334
rect 14108 3194 14136 3470
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 14200 800 14228 2926
rect 14844 800 14872 16546
rect 15580 11014 15608 24210
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16776 23866 16804 24074
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15672 21078 15700 21490
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15764 19446 15792 23054
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15948 22234 15976 22986
rect 17328 22982 17356 27814
rect 17972 27538 18000 28154
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 18064 27470 18092 28086
rect 18248 28082 18276 28426
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 17972 27130 18000 27270
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 17776 27056 17828 27062
rect 17776 26998 17828 27004
rect 17788 25906 17816 26998
rect 18156 26858 18184 27950
rect 18340 27334 18368 28698
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 18144 26852 18196 26858
rect 18144 26794 18196 26800
rect 18432 26234 18460 29582
rect 18696 29028 18748 29034
rect 18696 28970 18748 28976
rect 18708 28626 18736 28970
rect 18696 28620 18748 28626
rect 18696 28562 18748 28568
rect 18512 28552 18564 28558
rect 18564 28512 18644 28540
rect 18512 28494 18564 28500
rect 18616 27946 18644 28512
rect 18604 27940 18656 27946
rect 18604 27882 18656 27888
rect 18616 27470 18644 27882
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18432 26206 18552 26234
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17420 25702 17448 25842
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17512 25362 17540 25774
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17408 25288 17460 25294
rect 17788 25276 17816 25842
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 17868 25288 17920 25294
rect 17788 25248 17868 25276
rect 17408 25230 17460 25236
rect 17868 25230 17920 25236
rect 17420 24342 17448 25230
rect 18064 24750 18092 25298
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17408 24336 17460 24342
rect 17408 24278 17460 24284
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 16316 21962 16344 22374
rect 16500 22030 16528 22374
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16040 20330 16068 21286
rect 16316 20942 16344 21898
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16132 19786 16160 20402
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16132 19446 16160 19722
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 15764 18902 15792 19382
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15856 18426 15884 18702
rect 16316 18630 16344 20878
rect 16592 20602 16620 22034
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16684 20398 16712 22918
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 16960 21622 16988 22510
rect 17236 22234 17264 22510
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17512 22166 17540 23666
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17592 23112 17644 23118
rect 17590 23080 17592 23089
rect 17644 23080 17646 23089
rect 17590 23015 17646 23024
rect 17500 22160 17552 22166
rect 17500 22102 17552 22108
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 17040 20426 17092 20432
rect 16672 20392 16724 20398
rect 17040 20368 17092 20374
rect 16672 20334 16724 20340
rect 16684 19786 16712 20334
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19854 16804 20266
rect 17052 20058 17080 20368
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17052 19938 17080 19994
rect 16960 19910 17080 19938
rect 17224 19916 17276 19922
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 19378 16712 19722
rect 16960 19378 16988 19910
rect 17224 19858 17276 19864
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16776 18834 16804 19246
rect 17052 18902 17080 19246
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 17144 18834 17172 19246
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17236 18766 17264 19858
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18902 17356 19110
rect 17696 18902 17724 21898
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17788 19378 17816 19654
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17880 19258 17908 23598
rect 18524 23322 18552 26206
rect 18616 26042 18644 27406
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18616 24886 18644 25094
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18800 23662 18828 41386
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19248 40044 19300 40050
rect 19248 39986 19300 39992
rect 18972 39364 19024 39370
rect 18972 39306 19024 39312
rect 18984 39098 19012 39306
rect 18972 39092 19024 39098
rect 18972 39034 19024 39040
rect 19260 38758 19288 39986
rect 19984 39840 20036 39846
rect 19984 39782 20036 39788
rect 19996 39370 20024 39782
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 20076 38888 20128 38894
rect 20076 38830 20128 38836
rect 20168 38888 20220 38894
rect 20168 38830 20220 38836
rect 19248 38752 19300 38758
rect 19248 38694 19300 38700
rect 19260 38350 19288 38694
rect 20088 38554 20116 38830
rect 20076 38548 20128 38554
rect 20076 38490 20128 38496
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19352 37942 19380 38150
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19340 37936 19392 37942
rect 19340 37878 19392 37884
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19352 37262 19380 37606
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19260 36310 19288 36722
rect 19352 36394 19380 37198
rect 19444 36786 19472 37742
rect 20180 37738 20208 38830
rect 20444 38412 20496 38418
rect 20444 38354 20496 38360
rect 20168 37732 20220 37738
rect 20168 37674 20220 37680
rect 20180 37346 20208 37674
rect 20088 37330 20208 37346
rect 20076 37324 20208 37330
rect 20128 37318 20208 37324
rect 20076 37266 20128 37272
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36922 20024 37062
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19432 36780 19484 36786
rect 19484 36740 19656 36768
rect 19432 36722 19484 36728
rect 19352 36366 19564 36394
rect 19248 36304 19300 36310
rect 19248 36246 19300 36252
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 19260 35494 19288 36110
rect 19352 35698 19380 36110
rect 19444 35698 19472 36366
rect 19536 36242 19564 36366
rect 19628 36310 19656 36740
rect 19616 36304 19668 36310
rect 19616 36246 19668 36252
rect 19984 36304 20036 36310
rect 19984 36246 20036 36252
rect 19524 36236 19576 36242
rect 19524 36178 19576 36184
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19996 35562 20024 36246
rect 19984 35556 20036 35562
rect 19984 35498 20036 35504
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19260 35086 19288 35430
rect 19340 35148 19392 35154
rect 19340 35090 19392 35096
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19156 35012 19208 35018
rect 19156 34954 19208 34960
rect 19168 34406 19196 34954
rect 19352 34746 19380 35090
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19156 34400 19208 34406
rect 19156 34342 19208 34348
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18892 31754 18920 32166
rect 18892 31726 19012 31754
rect 18984 31142 19012 31726
rect 18972 31136 19024 31142
rect 18972 31078 19024 31084
rect 18984 30190 19012 31078
rect 18972 30184 19024 30190
rect 18972 30126 19024 30132
rect 18984 28218 19012 30126
rect 19076 29170 19104 33594
rect 19800 33312 19852 33318
rect 19800 33254 19852 33260
rect 19812 32978 19840 33254
rect 20088 32978 20116 37266
rect 20260 36780 20312 36786
rect 20260 36722 20312 36728
rect 20168 34536 20220 34542
rect 20168 34478 20220 34484
rect 20180 34202 20208 34478
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 19800 32972 19852 32978
rect 19800 32914 19852 32920
rect 20076 32972 20128 32978
rect 20076 32914 20128 32920
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19168 31890 19196 32302
rect 19260 32026 19288 32370
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 20088 32026 20116 32166
rect 19248 32020 19300 32026
rect 19248 31962 19300 31968
rect 20076 32020 20128 32026
rect 20076 31962 20128 31968
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19168 31482 19196 31826
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 19444 31346 19472 31826
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19444 30666 19472 31282
rect 20168 30728 20220 30734
rect 20168 30670 20220 30676
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19352 30326 19380 30534
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19444 30138 19472 30602
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19352 30110 19472 30138
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 19076 28082 19104 29106
rect 19260 28422 19288 29582
rect 19352 29510 19380 30110
rect 20180 29850 20208 30670
rect 20168 29844 20220 29850
rect 20168 29786 20220 29792
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19352 28558 19380 29446
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19076 27878 19104 28018
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 19352 27470 19380 28494
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19536 27674 19564 27950
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 20076 27328 20128 27334
rect 20076 27270 20128 27276
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19260 25702 19288 25842
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19616 25764 19668 25770
rect 19616 25706 19668 25712
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25362 19564 25638
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19628 25226 19656 25706
rect 19996 25498 20024 25774
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19616 25220 19668 25226
rect 19616 25162 19668 25168
rect 19444 24410 19472 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19536 24342 19564 24550
rect 19524 24336 19576 24342
rect 19524 24278 19576 24284
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18524 19922 18552 23258
rect 19536 23186 19564 23462
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 20088 23050 20116 27270
rect 20272 26234 20300 36722
rect 20456 36718 20484 38354
rect 20548 38350 20576 47126
rect 20996 47048 21048 47054
rect 20996 46990 21048 46996
rect 20628 46980 20680 46986
rect 20628 46922 20680 46928
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 20548 37738 20576 38150
rect 20536 37732 20588 37738
rect 20536 37674 20588 37680
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20352 36100 20404 36106
rect 20352 36042 20404 36048
rect 20364 35698 20392 36042
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20444 35624 20496 35630
rect 20444 35566 20496 35572
rect 20456 35290 20484 35566
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20444 35284 20496 35290
rect 20444 35226 20496 35232
rect 20352 35148 20404 35154
rect 20352 35090 20404 35096
rect 20364 33998 20392 35090
rect 20456 34610 20484 35226
rect 20548 35086 20576 35430
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20444 34604 20496 34610
rect 20444 34546 20496 34552
rect 20444 34060 20496 34066
rect 20548 34048 20576 35022
rect 20496 34020 20576 34048
rect 20444 34002 20496 34008
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20352 32836 20404 32842
rect 20352 32778 20404 32784
rect 20364 32434 20392 32778
rect 20548 32434 20576 32846
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20352 30592 20404 30598
rect 20352 30534 20404 30540
rect 20364 30258 20392 30534
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20548 28150 20576 28358
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20272 26206 20576 26234
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18616 22098 18644 22646
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18708 19990 18736 22986
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19168 22642 19196 22918
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19168 22030 19196 22578
rect 19904 22234 19932 22578
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 19892 22228 19944 22234
rect 19892 22170 19944 22176
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19444 20942 19472 21422
rect 19996 21350 20024 21966
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21554 20116 21830
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20534 19380 20742
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18064 19310 18092 19858
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17788 19230 17908 19258
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 16316 18290 16344 18566
rect 17604 18290 17632 18566
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2582 15240 2926
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 800 15516 2314
rect 16132 800 16160 2382
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 1970 16896 2246
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17420 800 17448 16186
rect 17788 15910 17816 19230
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17880 4146 17908 18838
rect 18340 18766 18368 19790
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18290 18092 18566
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18432 18222 18460 18362
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17604 3534 17632 3878
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 2990 17816 3470
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 3058 18276 3334
rect 18340 3194 18368 4082
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18708 3126 18736 19926
rect 19260 19786 19288 20334
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19260 19310 19288 19722
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19352 18902 19380 19382
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19444 16590 19472 20878
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 20088 19854 20116 21490
rect 20180 21486 20208 22374
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 20088 19378 20116 19790
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18358 20024 18566
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19892 18080 19944 18086
rect 20088 18068 20116 18770
rect 19944 18040 20116 18068
rect 19892 18022 19944 18028
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19996 16658 20024 18040
rect 20272 17746 20300 24550
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20364 21418 20392 23666
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 17338 20208 17546
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15706 19380 15982
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19444 15586 19472 16526
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19352 15558 19472 15586
rect 19352 15502 19380 15558
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 15026 19380 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18892 3058 18920 3878
rect 19260 3738 19288 4082
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19352 3194 19380 4558
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19338 3088 19394 3097
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18880 3052 18932 3058
rect 19338 3023 19394 3032
rect 18880 2994 18932 3000
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18708 800 18736 2790
rect 19352 800 19380 3023
rect 19444 2446 19472 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 4264 20024 15982
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19904 4236 20024 4264
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19812 3534 19840 4150
rect 19800 3528 19852 3534
rect 19904 3505 19932 4236
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19800 3470 19852 3476
rect 19890 3496 19946 3505
rect 19890 3431 19946 3440
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 2650 20024 4082
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20088 2446 20116 4966
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20180 3058 20208 3470
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20272 2582 20300 5170
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20364 3738 20392 4558
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20364 3194 20392 3402
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20260 2576 20312 2582
rect 20260 2518 20312 2524
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 870 20208 898
rect 19996 800 20024 870
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20180 762 20208 870
rect 20456 762 20484 3538
rect 20548 2650 20576 26206
rect 20640 4570 20668 46922
rect 21008 46034 21036 46990
rect 21284 46034 21312 49200
rect 21916 47252 21968 47258
rect 21916 47194 21968 47200
rect 20996 46028 21048 46034
rect 20996 45970 21048 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 21928 41414 21956 47194
rect 24584 47048 24636 47054
rect 24584 46990 24636 46996
rect 24596 46578 24624 46990
rect 24584 46572 24636 46578
rect 24584 46514 24636 46520
rect 25148 46510 25176 49200
rect 25412 47048 25464 47054
rect 25412 46990 25464 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25424 46034 25452 46990
rect 25792 46034 25820 49200
rect 25412 46028 25464 46034
rect 25412 45970 25464 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 24584 45960 24636 45966
rect 24584 45902 24636 45908
rect 24596 45626 24624 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 24584 45620 24636 45626
rect 24584 45562 24636 45568
rect 24596 45354 24624 45562
rect 25424 45558 25452 45834
rect 25412 45552 25464 45558
rect 25412 45494 25464 45500
rect 25780 45484 25832 45490
rect 25780 45426 25832 45432
rect 24584 45348 24636 45354
rect 24584 45290 24636 45296
rect 21836 41386 21956 41414
rect 20996 39296 21048 39302
rect 20996 39238 21048 39244
rect 21008 39098 21036 39238
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21008 37874 21036 39034
rect 21836 38962 21864 41386
rect 23480 40112 23532 40118
rect 23480 40054 23532 40060
rect 23492 39642 23520 40054
rect 23848 39976 23900 39982
rect 23848 39918 23900 39924
rect 25136 39976 25188 39982
rect 25136 39918 25188 39924
rect 23480 39636 23532 39642
rect 23480 39578 23532 39584
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 21824 38956 21876 38962
rect 21824 38898 21876 38904
rect 21180 38344 21232 38350
rect 21180 38286 21232 38292
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 21008 36242 21036 37810
rect 20996 36236 21048 36242
rect 20996 36178 21048 36184
rect 21008 35562 21036 36178
rect 21192 36174 21220 38286
rect 21836 37942 21864 38898
rect 22008 38888 22060 38894
rect 22008 38830 22060 38836
rect 22020 38350 22048 38830
rect 22112 38758 22140 39374
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 23296 38752 23348 38758
rect 23296 38694 23348 38700
rect 22008 38344 22060 38350
rect 22008 38286 22060 38292
rect 21824 37936 21876 37942
rect 21824 37878 21876 37884
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 21100 35766 21128 35974
rect 21192 35834 21220 36110
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21088 35760 21140 35766
rect 21088 35702 21140 35708
rect 20996 35556 21048 35562
rect 20996 35498 21048 35504
rect 21192 35290 21220 35770
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 21272 34400 21324 34406
rect 21272 34342 21324 34348
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33658 20760 33798
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 20824 33386 20852 34138
rect 21284 33998 21312 34342
rect 21376 34202 21404 35770
rect 21456 34944 21508 34950
rect 21456 34886 21508 34892
rect 21364 34196 21416 34202
rect 21364 34138 21416 34144
rect 21468 33998 21496 34886
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 20812 33380 20864 33386
rect 20812 33322 20864 33328
rect 20916 33046 20944 33866
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 33114 21036 33458
rect 21088 33448 21140 33454
rect 21088 33390 21140 33396
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 20904 33040 20956 33046
rect 20904 32982 20956 32988
rect 20916 32434 20944 32982
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 21008 31822 21036 32166
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 20732 29646 20760 31758
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 20824 29714 20852 29786
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 16574 20760 29446
rect 20916 29238 20944 29990
rect 21100 29714 21128 33390
rect 21468 32978 21496 33934
rect 21456 32972 21508 32978
rect 21456 32914 21508 32920
rect 21468 32434 21496 32914
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21836 29850 21864 37878
rect 22112 36786 22140 38694
rect 23308 38282 23336 38694
rect 23492 38418 23520 38898
rect 23860 38894 23888 39918
rect 25148 39642 25176 39918
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 25136 39024 25188 39030
rect 25136 38966 25188 38972
rect 23848 38888 23900 38894
rect 23848 38830 23900 38836
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 24768 38888 24820 38894
rect 24768 38830 24820 38836
rect 24136 38554 24164 38830
rect 24124 38548 24176 38554
rect 24124 38490 24176 38496
rect 24780 38418 24808 38830
rect 25148 38554 25176 38966
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38554 25360 38694
rect 25136 38548 25188 38554
rect 25136 38490 25188 38496
rect 25320 38548 25372 38554
rect 25320 38490 25372 38496
rect 23480 38412 23532 38418
rect 23480 38354 23532 38360
rect 24768 38412 24820 38418
rect 24768 38354 24820 38360
rect 22376 38276 22428 38282
rect 22376 38218 22428 38224
rect 23296 38276 23348 38282
rect 23296 38218 23348 38224
rect 22388 38010 22416 38218
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22204 37738 22232 37946
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22192 37732 22244 37738
rect 22192 37674 22244 37680
rect 22572 37466 22600 37810
rect 23492 37670 23520 38354
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 22560 37460 22612 37466
rect 22560 37402 22612 37408
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22204 36106 22232 36518
rect 22468 36236 22520 36242
rect 22468 36178 22520 36184
rect 22192 36100 22244 36106
rect 22192 36042 22244 36048
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22388 35698 22416 35974
rect 22480 35834 22508 36178
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22192 35624 22244 35630
rect 22192 35566 22244 35572
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22020 34610 22048 35226
rect 22204 35154 22232 35566
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 22204 34678 22232 35090
rect 23492 35086 23520 37606
rect 23676 37330 23704 37606
rect 23664 37324 23716 37330
rect 23664 37266 23716 37272
rect 23768 37262 23796 38150
rect 24964 38010 24992 38286
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 25332 37874 25360 38490
rect 25792 37942 25820 45426
rect 26608 40520 26660 40526
rect 26608 40462 26660 40468
rect 26240 40384 26292 40390
rect 26240 40326 26292 40332
rect 26056 39636 26108 39642
rect 26056 39578 26108 39584
rect 25964 38276 26016 38282
rect 25964 38218 26016 38224
rect 25780 37936 25832 37942
rect 25780 37878 25832 37884
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 23756 37256 23808 37262
rect 23756 37198 23808 37204
rect 24676 37256 24728 37262
rect 24676 37198 24728 37204
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 23572 37120 23624 37126
rect 23572 37062 23624 37068
rect 23584 36922 23612 37062
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23768 36854 23796 37198
rect 23756 36848 23808 36854
rect 23756 36790 23808 36796
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 22928 35012 22980 35018
rect 22928 34954 22980 34960
rect 22192 34672 22244 34678
rect 22192 34614 22244 34620
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22560 34468 22612 34474
rect 22560 34410 22612 34416
rect 22572 34082 22600 34410
rect 22848 34202 22876 34478
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 22572 34054 22876 34082
rect 22848 33998 22876 34054
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22756 33658 22784 33934
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22848 32842 22876 33934
rect 22940 33318 22968 34954
rect 23572 34944 23624 34950
rect 23572 34886 23624 34892
rect 23584 34678 23612 34886
rect 23572 34672 23624 34678
rect 23572 34614 23624 34620
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 22836 32836 22888 32842
rect 22836 32778 22888 32784
rect 22940 31890 22968 33254
rect 23020 32836 23072 32842
rect 23020 32778 23072 32784
rect 22928 31884 22980 31890
rect 22928 31826 22980 31832
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22020 30308 22048 31758
rect 22284 31748 22336 31754
rect 22284 31690 22336 31696
rect 22296 31482 22324 31690
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22020 30280 22140 30308
rect 22112 30190 22140 30280
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 21824 29844 21876 29850
rect 21824 29786 21876 29792
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 21088 29572 21140 29578
rect 21088 29514 21140 29520
rect 21100 29238 21128 29514
rect 20904 29232 20956 29238
rect 20904 29174 20956 29180
rect 21088 29232 21140 29238
rect 21088 29174 21140 29180
rect 20916 28558 20944 29174
rect 21100 28626 21128 29174
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 21100 28014 21128 28562
rect 21284 28490 21312 28902
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21192 27538 21220 28358
rect 21284 28150 21312 28426
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 21180 27532 21232 27538
rect 21180 27474 21232 27480
rect 21560 27402 21588 28494
rect 21744 27878 21772 29650
rect 22296 29646 22324 29990
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22008 29504 22060 29510
rect 22008 29446 22060 29452
rect 22020 29170 22048 29446
rect 22112 29306 22140 29582
rect 22100 29300 22152 29306
rect 22100 29242 22152 29248
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22296 29102 22324 29582
rect 22284 29096 22336 29102
rect 22284 29038 22336 29044
rect 22376 29096 22428 29102
rect 22376 29038 22428 29044
rect 22296 28694 22324 29038
rect 22284 28688 22336 28694
rect 22284 28630 22336 28636
rect 22388 28150 22416 29038
rect 22664 28218 22692 30126
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22756 28762 22784 29106
rect 23032 28994 23060 32778
rect 23308 32774 23336 33934
rect 23756 33924 23808 33930
rect 23756 33866 23808 33872
rect 23768 33658 23796 33866
rect 23756 33652 23808 33658
rect 23756 33594 23808 33600
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23584 33318 23612 33526
rect 23860 33522 23888 33594
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23676 32910 23704 33458
rect 23860 33114 23888 33458
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 22940 28966 23060 28994
rect 23308 28994 23336 32710
rect 23676 32570 23704 32846
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23572 31748 23624 31754
rect 23572 31690 23624 31696
rect 23584 30938 23612 31690
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23308 28966 23612 28994
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22744 28756 22796 28762
rect 22744 28698 22796 28704
rect 22848 28558 22876 28902
rect 22940 28558 22968 28966
rect 23112 28688 23164 28694
rect 23112 28630 23164 28636
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21732 27872 21784 27878
rect 21732 27814 21784 27820
rect 21744 27538 21772 27814
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 22020 27470 22048 28018
rect 22008 27464 22060 27470
rect 22008 27406 22060 27412
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21008 25430 21036 25842
rect 20996 25424 21048 25430
rect 20996 25366 21048 25372
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20824 24206 20852 24754
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21622 21036 21898
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21100 21434 21128 27270
rect 21560 25906 21588 27338
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 21192 24410 21220 24686
rect 21284 24410 21312 24754
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 22020 24206 22048 25434
rect 22296 25362 22324 25842
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22388 25226 22416 28086
rect 22664 28014 22692 28154
rect 22940 28150 22968 28358
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22664 26994 22692 27950
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22940 25906 22968 26522
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22928 25900 22980 25906
rect 22928 25842 22980 25848
rect 22572 25430 22600 25842
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 22940 25226 22968 25842
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 22928 25220 22980 25226
rect 22928 25162 22980 25168
rect 22940 24954 22968 25162
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 21744 22658 21772 24142
rect 22572 23866 22600 24822
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21836 22778 21864 23054
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21744 22642 21864 22658
rect 22296 22642 22324 23666
rect 23124 23662 23152 28630
rect 23584 28558 23612 28966
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23308 28218 23336 28494
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23860 27062 23888 27270
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 23216 25158 23244 25842
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23216 24206 23244 25094
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23492 24206 23520 24890
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23216 23730 23244 24142
rect 23308 23798 23336 24142
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 23848 23792 23900 23798
rect 23848 23734 23900 23740
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23112 23656 23164 23662
rect 23112 23598 23164 23604
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 22836 23044 22888 23050
rect 22836 22986 22888 22992
rect 22848 22778 22876 22986
rect 23400 22778 23428 23054
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23584 22642 23612 22918
rect 23860 22642 23888 23734
rect 21744 22636 21876 22642
rect 21744 22630 21824 22636
rect 21824 22578 21876 22584
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 21836 22506 21864 22578
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 22744 22500 22796 22506
rect 22744 22442 22796 22448
rect 21836 21554 21864 22442
rect 22756 21554 22784 22442
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 21100 21406 21220 21434
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21100 21010 21128 21286
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 18834 20852 19654
rect 20916 19174 20944 19790
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20916 18290 20944 19110
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 21008 17202 21036 19858
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21008 16658 21036 17138
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20732 16546 20852 16574
rect 20640 4542 20760 4570
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4146 20668 4422
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20626 4040 20682 4049
rect 20732 4026 20760 4542
rect 20682 3998 20760 4026
rect 20626 3975 20682 3984
rect 20824 3602 20852 16546
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21008 4282 21036 4558
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 21100 4146 21128 4422
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20916 3398 20944 4014
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 21192 2446 21220 21406
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20602 22140 20810
rect 22756 20806 22784 21490
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21836 18426 21864 19246
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 22112 17882 22140 19246
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21744 14482 21772 14758
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21284 2854 21312 4626
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4282 21680 4558
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21928 3398 21956 17546
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17134 22232 17478
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 21916 3392 21968 3398
rect 22020 3369 22048 16458
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 21916 3334 21968 3340
rect 22006 3360 22062 3369
rect 22006 3295 22062 3304
rect 22204 3058 22232 4490
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22296 4146 22324 4422
rect 22388 4214 22416 18634
rect 22756 16114 22784 20742
rect 22848 20466 22876 22578
rect 23756 22024 23808 22030
rect 23860 22012 23888 22578
rect 23808 21984 23888 22012
rect 23756 21966 23808 21972
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23124 21010 23152 21286
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23492 20534 23520 21286
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22848 19854 22876 20402
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22940 20058 22968 20334
rect 23676 20058 23704 20470
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22848 18766 22876 19790
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 23124 18902 23152 19382
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23308 18358 23336 18566
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23400 18222 23428 19178
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23400 17746 23428 18158
rect 23768 17814 23796 21830
rect 23860 21622 23888 21830
rect 23848 21616 23900 21622
rect 23848 21558 23900 21564
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22940 16046 22968 16390
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22480 3534 22508 4422
rect 22572 4282 22600 4558
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22572 3670 22600 4082
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 20640 800 20668 2382
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21928 800 21956 2314
rect 22020 2310 22048 2926
rect 22388 2650 22416 2994
rect 22664 2774 22692 14418
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 22572 2746 22692 2774
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 22572 800 22600 2746
rect 23032 2650 23060 5170
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23124 3534 23152 3878
rect 23216 3670 23244 4558
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23308 3058 23336 4422
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23400 3126 23428 4082
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23492 2774 23520 5170
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23768 3058 23796 5034
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23216 2746 23520 2774
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23216 800 23244 2746
rect 23584 2446 23612 2790
rect 23860 2514 23888 3878
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23952 2106 23980 36722
rect 24688 36378 24716 37198
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 24780 36922 24808 37062
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 25148 36854 25176 37198
rect 24860 36848 24912 36854
rect 24860 36790 24912 36796
rect 25136 36848 25188 36854
rect 25136 36790 25188 36796
rect 24872 36582 24900 36790
rect 25332 36786 25360 37810
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 24872 36174 24900 36518
rect 25056 36310 25084 36722
rect 25424 36378 25452 37742
rect 25596 37188 25648 37194
rect 25596 37130 25648 37136
rect 25608 36718 25636 37130
rect 25976 36786 26004 38218
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 25596 36712 25648 36718
rect 25596 36654 25648 36660
rect 25412 36372 25464 36378
rect 25412 36314 25464 36320
rect 25044 36304 25096 36310
rect 25044 36246 25096 36252
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 25056 36106 25084 36246
rect 25044 36100 25096 36106
rect 25044 36042 25096 36048
rect 24124 35080 24176 35086
rect 24124 35022 24176 35028
rect 24136 34678 24164 35022
rect 24124 34672 24176 34678
rect 24124 34614 24176 34620
rect 25056 34610 25084 36042
rect 25504 34740 25556 34746
rect 25504 34682 25556 34688
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 24216 34468 24268 34474
rect 24216 34410 24268 34416
rect 24228 33658 24256 34410
rect 24308 34400 24360 34406
rect 24308 34342 24360 34348
rect 24320 33930 24348 34342
rect 24780 34202 24808 34546
rect 25228 34536 25280 34542
rect 25228 34478 25280 34484
rect 24952 34400 25004 34406
rect 24952 34342 25004 34348
rect 24768 34196 24820 34202
rect 24768 34138 24820 34144
rect 24308 33924 24360 33930
rect 24308 33866 24360 33872
rect 24216 33652 24268 33658
rect 24216 33594 24268 33600
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 24044 31822 24072 32370
rect 24136 32026 24164 33458
rect 24320 33046 24348 33866
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 24308 33040 24360 33046
rect 24308 32982 24360 32988
rect 24584 32360 24636 32366
rect 24584 32302 24636 32308
rect 24216 32224 24268 32230
rect 24216 32166 24268 32172
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24032 31816 24084 31822
rect 24032 31758 24084 31764
rect 24136 31414 24164 31962
rect 24228 31822 24256 32166
rect 24596 31958 24624 32302
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24124 31408 24176 31414
rect 24124 31350 24176 31356
rect 24596 31346 24624 31894
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24308 30728 24360 30734
rect 24308 30670 24360 30676
rect 24320 29646 24348 30670
rect 24400 30320 24452 30326
rect 24400 30262 24452 30268
rect 24412 29850 24440 30262
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 24320 28558 24348 29582
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24308 28552 24360 28558
rect 24308 28494 24360 28500
rect 24320 26586 24348 28494
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24412 26382 24440 29446
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 28150 24532 28358
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24044 25498 24072 25774
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 24044 23662 24072 25434
rect 24688 24682 24716 33458
rect 24964 32910 24992 34342
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24780 31278 24808 31894
rect 25136 31680 25188 31686
rect 25136 31622 25188 31628
rect 25148 31482 25176 31622
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 24768 31272 24820 31278
rect 24768 31214 24820 31220
rect 25240 30666 25268 34478
rect 25412 33924 25464 33930
rect 25412 33866 25464 33872
rect 25424 33114 25452 33866
rect 25412 33108 25464 33114
rect 25412 33050 25464 33056
rect 25516 32994 25544 34682
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 25424 32966 25544 32994
rect 25228 30660 25280 30666
rect 25228 30602 25280 30608
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24872 30190 24900 30534
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 25332 28506 25360 32914
rect 25424 32910 25452 32966
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25424 32774 25452 32846
rect 25412 32768 25464 32774
rect 25412 32710 25464 32716
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25516 32434 25544 32710
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25608 32230 25636 36654
rect 25976 36582 26004 36722
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25964 32972 26016 32978
rect 25964 32914 26016 32920
rect 25976 32502 26004 32914
rect 25964 32496 26016 32502
rect 25964 32438 26016 32444
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25596 32224 25648 32230
rect 25596 32166 25648 32172
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25424 31346 25452 31826
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25516 31210 25544 32166
rect 25608 31890 25636 32166
rect 25596 31884 25648 31890
rect 25596 31826 25648 31832
rect 25792 31822 25820 32234
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25608 31278 25636 31622
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25504 31204 25556 31210
rect 25504 31146 25556 31152
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25976 30734 26004 31078
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25688 30660 25740 30666
rect 25688 30602 25740 30608
rect 25700 30054 25728 30602
rect 25688 30048 25740 30054
rect 25688 29990 25740 29996
rect 26068 29850 26096 39578
rect 26252 39574 26280 40326
rect 26424 40180 26476 40186
rect 26424 40122 26476 40128
rect 26240 39568 26292 39574
rect 26240 39510 26292 39516
rect 26436 39438 26464 40122
rect 26620 39642 26648 40462
rect 26608 39636 26660 39642
rect 26608 39578 26660 39584
rect 26424 39432 26476 39438
rect 26424 39374 26476 39380
rect 26436 38350 26464 39374
rect 26516 38412 26568 38418
rect 26516 38354 26568 38360
rect 26424 38344 26476 38350
rect 26424 38286 26476 38292
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 26160 36310 26188 36518
rect 26252 36378 26280 36722
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26148 36304 26200 36310
rect 26148 36246 26200 36252
rect 26436 34678 26464 38150
rect 26528 37262 26556 38354
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26528 36922 26556 37198
rect 26516 36916 26568 36922
rect 26516 36858 26568 36864
rect 26528 36802 26556 36858
rect 26528 36774 26648 36802
rect 26620 36718 26648 36774
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26528 36106 26556 36654
rect 26516 36100 26568 36106
rect 26516 36042 26568 36048
rect 26424 34672 26476 34678
rect 26424 34614 26476 34620
rect 26424 34536 26476 34542
rect 26424 34478 26476 34484
rect 26436 33930 26464 34478
rect 26424 33924 26476 33930
rect 26424 33866 26476 33872
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26148 32836 26200 32842
rect 26148 32778 26200 32784
rect 26160 32434 26188 32778
rect 26252 32434 26280 33254
rect 26344 32910 26372 33798
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 26160 30734 26188 32370
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26160 30394 26188 30670
rect 26148 30388 26200 30394
rect 26148 30330 26200 30336
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26528 29782 26556 36042
rect 26516 29776 26568 29782
rect 26516 29718 26568 29724
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 26329 29640 26381 29646
rect 26329 29582 26381 29588
rect 26160 29034 26188 29582
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26148 29028 26200 29034
rect 26148 28970 26200 28976
rect 26252 28966 26280 29446
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 26344 28762 26372 29582
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26436 28626 26464 28970
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26332 28552 26384 28558
rect 25332 28478 25452 28506
rect 26332 28494 26384 28500
rect 25320 28416 25372 28422
rect 25320 28358 25372 28364
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25148 27470 25176 27814
rect 25332 27538 25360 28358
rect 25320 27532 25372 27538
rect 25320 27474 25372 27480
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25332 27130 25360 27338
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25240 26586 25268 26998
rect 25424 26874 25452 28478
rect 25596 28008 25648 28014
rect 25596 27950 25648 27956
rect 25608 27674 25636 27950
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 26344 27606 26372 28494
rect 26516 28416 26568 28422
rect 26516 28358 26568 28364
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 25332 26846 25452 26874
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25056 25294 25084 26318
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 24400 24336 24452 24342
rect 24400 24278 24452 24284
rect 24412 24138 24440 24278
rect 25148 24274 25176 24550
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24032 23656 24084 23662
rect 24032 23598 24084 23604
rect 24044 17882 24072 23598
rect 24216 23248 24268 23254
rect 24216 23190 24268 23196
rect 24228 21962 24256 23190
rect 24412 22438 24440 24074
rect 24676 23520 24728 23526
rect 24676 23462 24728 23468
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24688 23186 24716 23462
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24504 22710 24532 22918
rect 24872 22778 24900 23462
rect 24964 23050 24992 24142
rect 25044 23248 25096 23254
rect 25044 23190 25096 23196
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24504 22094 24532 22646
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24412 22066 24532 22094
rect 24412 21962 24440 22066
rect 24688 22030 24716 22510
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24412 20398 24440 21898
rect 24780 21554 24808 22374
rect 24872 21962 24900 22714
rect 25056 22506 25084 23190
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 25240 22094 25268 24686
rect 25056 22066 25268 22094
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24320 17270 24348 19110
rect 24412 18902 24440 19314
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24412 17542 24440 18634
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 17592 24624 18566
rect 24780 17678 24808 19314
rect 24872 18290 24900 19790
rect 25056 18834 25084 22066
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24676 17604 24728 17610
rect 24596 17564 24676 17592
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24412 16998 24440 17478
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16522 24440 16934
rect 24596 16794 24624 17564
rect 24676 17546 24728 17552
rect 24780 16794 24808 17614
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24400 16516 24452 16522
rect 24400 16458 24452 16464
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24412 3194 24440 4014
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24504 3194 24532 3334
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24596 3058 24624 3878
rect 24688 3534 24716 3946
rect 24780 3602 24808 4966
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24676 3528 24728 3534
rect 24674 3496 24676 3505
rect 24728 3496 24730 3505
rect 24674 3431 24730 3440
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3126 24808 3334
rect 25240 3126 25268 4082
rect 25332 3942 25360 26846
rect 26528 26450 26556 28358
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26516 26444 26568 26450
rect 26516 26386 26568 26392
rect 26620 26382 26648 27610
rect 26712 27606 26740 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 28368 47054 28396 49200
rect 28908 47184 28960 47190
rect 28908 47126 28960 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 26884 45824 26936 45830
rect 26884 45766 26936 45772
rect 26896 40390 26924 45766
rect 28920 41414 28948 47126
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49314 43250 50000
rect 43138 49286 43576 49314
rect 43138 49200 43250 49286
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 29368 46980 29420 46986
rect 29368 46922 29420 46928
rect 28828 41386 28948 41414
rect 26976 40588 27028 40594
rect 26976 40530 27028 40536
rect 26884 40384 26936 40390
rect 26884 40326 26936 40332
rect 26792 36644 26844 36650
rect 26792 36586 26844 36592
rect 26804 36106 26832 36586
rect 26792 36100 26844 36106
rect 26792 36042 26844 36048
rect 26988 33454 27016 40530
rect 27252 38888 27304 38894
rect 27252 38830 27304 38836
rect 27344 38888 27396 38894
rect 27344 38830 27396 38836
rect 27160 38208 27212 38214
rect 27160 38150 27212 38156
rect 27172 37874 27200 38150
rect 27264 38010 27292 38830
rect 27356 38350 27384 38830
rect 27528 38412 27580 38418
rect 27528 38354 27580 38360
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27344 38208 27396 38214
rect 27344 38150 27396 38156
rect 27252 38004 27304 38010
rect 27252 37946 27304 37952
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27356 37466 27384 38150
rect 27540 37806 27568 38354
rect 27528 37800 27580 37806
rect 27528 37742 27580 37748
rect 27344 37460 27396 37466
rect 27344 37402 27396 37408
rect 27344 37324 27396 37330
rect 27344 37266 27396 37272
rect 27356 36786 27384 37266
rect 27344 36780 27396 36786
rect 27344 36722 27396 36728
rect 27068 36032 27120 36038
rect 27068 35974 27120 35980
rect 26976 33448 27028 33454
rect 26976 33390 27028 33396
rect 26988 32026 27016 33390
rect 26976 32020 27028 32026
rect 26976 31962 27028 31968
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26988 31346 27016 31758
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 26988 30938 27016 31282
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 27080 30802 27108 35974
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 27160 34196 27212 34202
rect 27160 34138 27212 34144
rect 27172 33318 27200 34138
rect 27264 33930 27292 34546
rect 27436 34468 27488 34474
rect 27436 34410 27488 34416
rect 27344 34400 27396 34406
rect 27344 34342 27396 34348
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27264 33114 27292 33866
rect 27356 33590 27384 34342
rect 27448 34202 27476 34410
rect 27436 34196 27488 34202
rect 27436 34138 27488 34144
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27344 33584 27396 33590
rect 27344 33526 27396 33532
rect 27448 33522 27476 33866
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27540 33114 27568 37742
rect 27896 37664 27948 37670
rect 27896 37606 27948 37612
rect 27712 34060 27764 34066
rect 27712 34002 27764 34008
rect 27724 33454 27752 34002
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27252 33108 27304 33114
rect 27252 33050 27304 33056
rect 27528 33108 27580 33114
rect 27528 33050 27580 33056
rect 27344 33040 27396 33046
rect 27344 32982 27396 32988
rect 26792 30796 26844 30802
rect 26792 30738 26844 30744
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 26700 27600 26752 27606
rect 26700 27542 26752 27548
rect 26608 26376 26660 26382
rect 26608 26318 26660 26324
rect 26620 25974 26648 26318
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 25412 25968 25464 25974
rect 25412 25910 25464 25916
rect 26608 25968 26660 25974
rect 26608 25910 26660 25916
rect 25424 25498 25452 25910
rect 26620 25770 26648 25910
rect 26608 25764 26660 25770
rect 26608 25706 26660 25712
rect 25412 25492 25464 25498
rect 25412 25434 25464 25440
rect 26712 24818 26740 26250
rect 26804 25498 26832 30738
rect 27356 30598 27384 32982
rect 27528 32836 27580 32842
rect 27528 32778 27580 32784
rect 27540 32450 27568 32778
rect 27448 32434 27568 32450
rect 27436 32428 27568 32434
rect 27488 32422 27568 32428
rect 27436 32370 27488 32376
rect 27448 31822 27476 32370
rect 27908 31958 27936 37606
rect 28172 37120 28224 37126
rect 28172 37062 28224 37068
rect 28080 36100 28132 36106
rect 28080 36042 28132 36048
rect 28092 35630 28120 36042
rect 28080 35624 28132 35630
rect 28080 35566 28132 35572
rect 27988 35012 28040 35018
rect 27988 34954 28040 34960
rect 28000 32910 28028 34954
rect 27988 32904 28040 32910
rect 27988 32846 28040 32852
rect 28000 32609 28028 32846
rect 27986 32600 28042 32609
rect 27986 32535 28042 32544
rect 27896 31952 27948 31958
rect 27896 31894 27948 31900
rect 27436 31816 27488 31822
rect 27436 31758 27488 31764
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27528 30728 27580 30734
rect 27528 30670 27580 30676
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 26976 30388 27028 30394
rect 26976 30330 27028 30336
rect 26884 29776 26936 29782
rect 26884 29718 26936 29724
rect 26896 29238 26924 29718
rect 26884 29232 26936 29238
rect 26884 29174 26936 29180
rect 26988 29170 27016 30330
rect 27356 30326 27384 30534
rect 27540 30394 27568 30670
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27344 30320 27396 30326
rect 27344 30262 27396 30268
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26988 29050 27016 29106
rect 26896 29022 27016 29050
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 26896 24206 26924 29022
rect 27080 28422 27108 29786
rect 27528 29504 27580 29510
rect 27172 29464 27528 29492
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 27080 27334 27108 28018
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 26976 26240 27028 26246
rect 26976 26182 27028 26188
rect 26988 25906 27016 26182
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26896 23798 26924 24142
rect 26884 23792 26936 23798
rect 26884 23734 26936 23740
rect 25688 23588 25740 23594
rect 25688 23530 25740 23536
rect 25412 23316 25464 23322
rect 25596 23316 25648 23322
rect 25464 23276 25596 23304
rect 25412 23258 25464 23264
rect 25596 23258 25648 23264
rect 25700 23254 25728 23530
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 26882 23216 26938 23225
rect 26882 23151 26938 23160
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25700 22642 25728 22918
rect 25778 22672 25834 22681
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25688 22636 25740 22642
rect 25778 22607 25834 22616
rect 25688 22578 25740 22584
rect 25516 22409 25544 22578
rect 25792 22574 25820 22607
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25872 22500 25924 22506
rect 25872 22442 25924 22448
rect 26148 22500 26200 22506
rect 26148 22442 26200 22448
rect 25502 22400 25558 22409
rect 25502 22335 25558 22344
rect 25884 20466 25912 22442
rect 26160 22234 26188 22442
rect 26252 22234 26280 23054
rect 26896 22710 26924 23151
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 26988 22778 27016 22986
rect 26976 22772 27028 22778
rect 26976 22714 27028 22720
rect 26884 22704 26936 22710
rect 27080 22681 27108 27270
rect 27172 26314 27200 29464
rect 27528 29446 27580 29452
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27264 28218 27292 28494
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27264 27538 27292 28154
rect 27356 27946 27384 29106
rect 27632 28642 27660 31282
rect 27540 28614 27660 28642
rect 27540 27962 27568 28614
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27632 28082 27660 28426
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27344 27940 27396 27946
rect 27540 27934 27660 27962
rect 27344 27882 27396 27888
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27160 26308 27212 26314
rect 27160 26250 27212 26256
rect 27252 26308 27304 26314
rect 27252 26250 27304 26256
rect 27264 25906 27292 26250
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27356 25702 27384 27882
rect 27632 27130 27660 27934
rect 27724 27606 27752 31758
rect 28000 31482 28028 32535
rect 27988 31476 28040 31482
rect 27988 31418 28040 31424
rect 28092 31362 28120 35566
rect 28000 31334 28120 31362
rect 27896 30660 27948 30666
rect 27896 30602 27948 30608
rect 27804 30320 27856 30326
rect 27804 30262 27856 30268
rect 27816 29714 27844 30262
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 27816 29170 27844 29650
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27816 28490 27844 29106
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27632 26382 27660 27066
rect 27908 27062 27936 30602
rect 28000 29850 28028 31334
rect 28080 31204 28132 31210
rect 28080 31146 28132 31152
rect 28092 30802 28120 31146
rect 28080 30796 28132 30802
rect 28080 30738 28132 30744
rect 28092 30258 28120 30738
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 27988 29844 28040 29850
rect 27988 29786 28040 29792
rect 28000 29170 28028 29786
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 28000 28082 28028 29106
rect 28080 28620 28132 28626
rect 28080 28562 28132 28568
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 28092 28014 28120 28562
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 27896 27056 27948 27062
rect 27896 26998 27948 27004
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 27908 26314 27936 26998
rect 27988 26444 28040 26450
rect 27988 26386 28040 26392
rect 27896 26308 27948 26314
rect 27896 26250 27948 26256
rect 27436 25900 27488 25906
rect 27436 25842 27488 25848
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 26884 22646 26936 22652
rect 27066 22672 27122 22681
rect 26516 22636 26568 22642
rect 27172 22642 27200 24550
rect 27066 22607 27122 22616
rect 27160 22636 27212 22642
rect 26516 22578 26568 22584
rect 27160 22578 27212 22584
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26436 22030 26464 22102
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 26160 21554 26188 21966
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 26068 21146 26096 21354
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26252 20602 26280 20878
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 25872 20460 25924 20466
rect 25792 20420 25872 20448
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25700 19922 25728 20198
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25792 18766 25820 20420
rect 25872 20402 25924 20408
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25424 17134 25452 18022
rect 25792 17746 25820 18702
rect 26252 18630 26280 20538
rect 26528 20534 26556 22578
rect 27068 22568 27120 22574
rect 27264 22522 27292 25366
rect 27356 22982 27384 25638
rect 27448 25430 27476 25842
rect 27436 25424 27488 25430
rect 27436 25366 27488 25372
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27448 22982 27476 23666
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27816 23186 27844 23462
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27804 23044 27856 23050
rect 27540 23004 27804 23032
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 27068 22510 27120 22516
rect 27080 22234 27108 22510
rect 27172 22494 27292 22522
rect 27068 22228 27120 22234
rect 27068 22170 27120 22176
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26896 20942 26924 21286
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26528 18834 26556 19654
rect 26896 19378 26924 20470
rect 26988 20466 27016 21558
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26988 19718 27016 20402
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 27080 19514 27108 19722
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26896 18714 26924 19314
rect 26896 18686 27016 18714
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26884 18624 26936 18630
rect 26884 18566 26936 18572
rect 26896 18426 26924 18566
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 25792 16522 25820 17682
rect 26252 16658 26280 17682
rect 26344 16794 26372 18022
rect 26988 17678 27016 18686
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26528 17270 26556 17478
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 14074 27108 14282
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27172 12434 27200 22494
rect 27356 22438 27384 22918
rect 27448 22778 27476 22918
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 27344 22432 27396 22438
rect 27344 22374 27396 22380
rect 27264 21146 27292 22374
rect 27448 21962 27476 22714
rect 27540 22234 27568 23004
rect 27804 22986 27856 22992
rect 27710 22672 27766 22681
rect 27710 22607 27766 22616
rect 27724 22574 27752 22607
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27894 22400 27950 22409
rect 27894 22335 27950 22344
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 27436 21956 27488 21962
rect 27436 21898 27488 21904
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27264 20466 27292 21082
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27264 16522 27292 17478
rect 27252 16516 27304 16522
rect 27252 16458 27304 16464
rect 27448 14482 27476 21898
rect 27540 21690 27568 22170
rect 27620 22160 27672 22166
rect 27620 22102 27672 22108
rect 27632 21962 27660 22102
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27908 21894 27936 22335
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27896 21888 27948 21894
rect 27896 21830 27948 21836
rect 27724 21690 27752 21830
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27540 20806 27568 21286
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27540 20602 27568 20742
rect 27816 20602 27844 20810
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27712 17808 27764 17814
rect 27712 17750 27764 17756
rect 27724 16454 27752 17750
rect 27908 17746 27936 21830
rect 28000 18154 28028 26386
rect 28092 26382 28120 27270
rect 28080 26376 28132 26382
rect 28080 26318 28132 26324
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 27988 18148 28040 18154
rect 27988 18090 28040 18096
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27816 17338 27844 17614
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 28000 17202 28028 17614
rect 28092 17610 28120 18226
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27724 16114 27752 16390
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27436 14476 27488 14482
rect 27436 14418 27488 14424
rect 26804 12406 27200 12434
rect 25596 4208 25648 4214
rect 25596 4150 25648 4156
rect 25502 4040 25558 4049
rect 25608 4026 25636 4150
rect 25558 3998 25636 4026
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 25502 3975 25558 3984
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24872 2990 24900 3062
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 24504 800 24532 2314
rect 25148 800 25176 2926
rect 25516 2446 25544 3975
rect 26620 3602 26648 4014
rect 26608 3596 26660 3602
rect 26608 3538 26660 3544
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26712 2582 26740 3470
rect 26700 2576 26752 2582
rect 26700 2518 26752 2524
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26436 800 26464 2382
rect 26804 1970 26832 12406
rect 27344 3528 27396 3534
rect 27342 3496 27344 3505
rect 27396 3496 27398 3505
rect 27342 3431 27398 3440
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26792 1964 26844 1970
rect 26792 1906 26844 1912
rect 27080 800 27108 2994
rect 28000 2514 28028 17138
rect 28184 2650 28212 37062
rect 28632 35012 28684 35018
rect 28632 34954 28684 34960
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 28276 32434 28304 32914
rect 28368 32570 28396 34546
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 28460 32910 28488 33390
rect 28448 32904 28500 32910
rect 28448 32846 28500 32852
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28460 32570 28488 32846
rect 28356 32564 28408 32570
rect 28356 32506 28408 32512
rect 28448 32564 28500 32570
rect 28448 32506 28500 32512
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28276 31890 28304 32370
rect 28264 31884 28316 31890
rect 28264 31826 28316 31832
rect 28368 30734 28396 32506
rect 28552 32230 28580 32846
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28448 30660 28500 30666
rect 28448 30602 28500 30608
rect 28460 30326 28488 30602
rect 28448 30320 28500 30326
rect 28448 30262 28500 30268
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 28368 29850 28396 30058
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 28552 29850 28580 29990
rect 28356 29844 28408 29850
rect 28356 29786 28408 29792
rect 28540 29844 28592 29850
rect 28540 29786 28592 29792
rect 28552 29578 28580 29786
rect 28264 29572 28316 29578
rect 28264 29514 28316 29520
rect 28448 29572 28500 29578
rect 28448 29514 28500 29520
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28276 28218 28304 29514
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28264 28212 28316 28218
rect 28264 28154 28316 28160
rect 28368 28082 28396 28358
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28264 27940 28316 27946
rect 28264 27882 28316 27888
rect 28276 26994 28304 27882
rect 28368 27470 28396 28018
rect 28460 27878 28488 29514
rect 28540 29096 28592 29102
rect 28540 29038 28592 29044
rect 28552 28490 28580 29038
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28552 27946 28580 28426
rect 28540 27940 28592 27946
rect 28540 27882 28592 27888
rect 28448 27872 28500 27878
rect 28448 27814 28500 27820
rect 28460 27470 28488 27814
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 28448 27464 28500 27470
rect 28448 27406 28500 27412
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28276 26382 28304 26930
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28276 23254 28304 23598
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28368 20534 28396 26862
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28460 25974 28488 26250
rect 28448 25968 28500 25974
rect 28448 25910 28500 25916
rect 28460 25362 28488 25910
rect 28448 25356 28500 25362
rect 28448 25298 28500 25304
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 28460 24138 28488 24754
rect 28448 24132 28500 24138
rect 28448 24074 28500 24080
rect 28460 22982 28488 24074
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 28644 22094 28672 34954
rect 28724 33448 28776 33454
rect 28724 33390 28776 33396
rect 28736 31346 28764 33390
rect 28724 31340 28776 31346
rect 28724 31282 28776 31288
rect 28736 29646 28764 31282
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 28736 29170 28764 29582
rect 28724 29164 28776 29170
rect 28724 29106 28776 29112
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 28736 27606 28764 28970
rect 28724 27600 28776 27606
rect 28724 27542 28776 27548
rect 28828 26926 28856 41386
rect 29000 38752 29052 38758
rect 29000 38694 29052 38700
rect 29012 38350 29040 38694
rect 29000 38344 29052 38350
rect 29000 38286 29052 38292
rect 29092 36372 29144 36378
rect 29092 36314 29144 36320
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 29012 35766 29040 36110
rect 29000 35760 29052 35766
rect 29000 35702 29052 35708
rect 29000 35556 29052 35562
rect 29000 35498 29052 35504
rect 29012 35290 29040 35498
rect 29000 35284 29052 35290
rect 29000 35226 29052 35232
rect 28908 34060 28960 34066
rect 28908 34002 28960 34008
rect 28920 33590 28948 34002
rect 29104 33590 29132 36314
rect 29184 35624 29236 35630
rect 29184 35566 29236 35572
rect 29196 35086 29224 35566
rect 29276 35148 29328 35154
rect 29276 35090 29328 35096
rect 29184 35080 29236 35086
rect 29184 35022 29236 35028
rect 29196 34678 29224 35022
rect 29184 34672 29236 34678
rect 29184 34614 29236 34620
rect 29288 34542 29316 35090
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29288 34134 29316 34478
rect 29276 34128 29328 34134
rect 29276 34070 29328 34076
rect 29184 33992 29236 33998
rect 29184 33934 29236 33940
rect 29196 33658 29224 33934
rect 29184 33652 29236 33658
rect 29184 33594 29236 33600
rect 28908 33584 28960 33590
rect 28908 33526 28960 33532
rect 29092 33584 29144 33590
rect 29092 33526 29144 33532
rect 28920 32910 28948 33526
rect 29196 33114 29224 33594
rect 29288 33590 29316 34070
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29184 33108 29236 33114
rect 29184 33050 29236 33056
rect 28908 32904 28960 32910
rect 28908 32846 28960 32852
rect 28998 32600 29054 32609
rect 28908 32564 28960 32570
rect 28998 32535 29000 32544
rect 28908 32506 28960 32512
rect 29052 32535 29054 32544
rect 29000 32506 29052 32512
rect 28920 31686 28948 32506
rect 29196 32366 29224 33050
rect 29184 32360 29236 32366
rect 29184 32302 29236 32308
rect 29184 32224 29236 32230
rect 29184 32166 29236 32172
rect 29092 31816 29144 31822
rect 29092 31758 29144 31764
rect 28908 31680 28960 31686
rect 28908 31622 28960 31628
rect 29000 30660 29052 30666
rect 29000 30602 29052 30608
rect 29012 29306 29040 30602
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28908 28620 28960 28626
rect 28908 28562 28960 28568
rect 28920 27538 28948 28562
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 29104 26926 29132 31758
rect 29196 30802 29224 32166
rect 29184 30796 29236 30802
rect 29184 30738 29236 30744
rect 29196 29170 29224 30738
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29196 28694 29224 29106
rect 29184 28688 29236 28694
rect 29184 28630 29236 28636
rect 29196 27946 29224 28630
rect 29184 27940 29236 27946
rect 29184 27882 29236 27888
rect 28816 26920 28868 26926
rect 28816 26862 28868 26868
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 28724 26240 28776 26246
rect 28724 26182 28776 26188
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28736 25974 28764 26182
rect 28920 26042 28948 26182
rect 29104 26042 29132 26862
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 28724 25968 28776 25974
rect 28724 25910 28776 25916
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28736 24138 28764 24754
rect 29092 24336 29144 24342
rect 29092 24278 29144 24284
rect 28724 24132 28776 24138
rect 28724 24074 28776 24080
rect 28736 23662 28764 24074
rect 28998 23760 29054 23769
rect 28816 23724 28868 23730
rect 28998 23695 29000 23704
rect 28816 23666 28868 23672
rect 29052 23695 29054 23704
rect 29000 23666 29052 23672
rect 28724 23656 28776 23662
rect 28724 23598 28776 23604
rect 28736 23322 28764 23598
rect 28828 23322 28856 23666
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28816 23316 28868 23322
rect 28816 23258 28868 23264
rect 28736 23225 28764 23258
rect 28722 23216 28778 23225
rect 28722 23151 28778 23160
rect 28828 22234 28856 23258
rect 28908 23248 28960 23254
rect 28908 23190 28960 23196
rect 28920 22710 28948 23190
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 29104 22642 29132 24278
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29288 23866 29316 24074
rect 29276 23860 29328 23866
rect 29276 23802 29328 23808
rect 29184 23792 29236 23798
rect 29184 23734 29236 23740
rect 29196 22778 29224 23734
rect 29288 23050 29316 23802
rect 29276 23044 29328 23050
rect 29276 22986 29328 22992
rect 29184 22772 29236 22778
rect 29184 22714 29236 22720
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 28816 22228 28868 22234
rect 28816 22170 28868 22176
rect 28644 22066 28764 22094
rect 28356 20528 28408 20534
rect 28356 20470 28408 20476
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28368 6866 28396 18634
rect 28540 18352 28592 18358
rect 28540 18294 28592 18300
rect 28552 18086 28580 18294
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28552 17202 28580 18022
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28644 17338 28672 17478
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28448 14340 28500 14346
rect 28448 14282 28500 14288
rect 28356 6860 28408 6866
rect 28356 6802 28408 6808
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 28092 2378 28120 2586
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28080 2372 28132 2378
rect 28080 2314 28132 2320
rect 28368 800 28396 2382
rect 28460 1902 28488 14282
rect 28552 4078 28580 17138
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28736 1970 28764 22066
rect 29380 20806 29408 46922
rect 32232 46442 32260 49200
rect 38028 47410 38056 49200
rect 37292 47382 38056 47410
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 36912 47252 36964 47258
rect 36912 47194 36964 47200
rect 35348 47184 35400 47190
rect 35348 47126 35400 47132
rect 34704 47048 34756 47054
rect 34704 46990 34756 46996
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 34428 46504 34480 46510
rect 34428 46446 34480 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 46170 32352 46446
rect 34440 46170 34468 46446
rect 32312 46164 32364 46170
rect 32312 46106 32364 46112
rect 34428 46164 34480 46170
rect 34428 46106 34480 46112
rect 32588 45960 32640 45966
rect 32588 45902 32640 45908
rect 32600 45422 32628 45902
rect 34716 45554 34744 46990
rect 34796 46504 34848 46510
rect 34796 46446 34848 46452
rect 34808 46170 34836 46446
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34796 46164 34848 46170
rect 34796 46106 34848 46112
rect 34716 45526 34836 45554
rect 32588 45416 32640 45422
rect 32588 45358 32640 45364
rect 29920 38956 29972 38962
rect 29920 38898 29972 38904
rect 29828 38820 29880 38826
rect 29828 38762 29880 38768
rect 29840 38418 29868 38762
rect 29932 38554 29960 38898
rect 30012 38888 30064 38894
rect 30012 38830 30064 38836
rect 30104 38888 30156 38894
rect 30104 38830 30156 38836
rect 29920 38548 29972 38554
rect 29920 38490 29972 38496
rect 29828 38412 29880 38418
rect 29828 38354 29880 38360
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 29656 36786 29684 37266
rect 29840 37262 29868 38354
rect 29932 37330 29960 38490
rect 30024 38010 30052 38830
rect 30012 38004 30064 38010
rect 30012 37946 30064 37952
rect 30012 37800 30064 37806
rect 30012 37742 30064 37748
rect 30024 37466 30052 37742
rect 30116 37670 30144 38830
rect 31116 38276 31168 38282
rect 31116 38218 31168 38224
rect 31128 38010 31156 38218
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 30932 37868 30984 37874
rect 30932 37810 30984 37816
rect 30104 37664 30156 37670
rect 30104 37606 30156 37612
rect 30012 37460 30064 37466
rect 30012 37402 30064 37408
rect 29920 37324 29972 37330
rect 29920 37266 29972 37272
rect 29828 37256 29880 37262
rect 29828 37198 29880 37204
rect 29644 36780 29696 36786
rect 29644 36722 29696 36728
rect 29656 36378 29684 36722
rect 29840 36718 29868 37198
rect 29828 36712 29880 36718
rect 29828 36654 29880 36660
rect 29644 36372 29696 36378
rect 29644 36314 29696 36320
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 29748 35018 29776 36110
rect 29840 35154 29868 36654
rect 29932 35766 29960 37266
rect 30116 36922 30144 37606
rect 30104 36916 30156 36922
rect 30104 36858 30156 36864
rect 30380 36848 30432 36854
rect 30380 36790 30432 36796
rect 30104 36712 30156 36718
rect 30104 36654 30156 36660
rect 30196 36712 30248 36718
rect 30196 36654 30248 36660
rect 30116 36378 30144 36654
rect 30104 36372 30156 36378
rect 30104 36314 30156 36320
rect 30208 36242 30236 36654
rect 30196 36236 30248 36242
rect 30196 36178 30248 36184
rect 30208 36122 30236 36178
rect 30208 36094 30328 36122
rect 30196 36032 30248 36038
rect 30196 35974 30248 35980
rect 30208 35766 30236 35974
rect 29920 35760 29972 35766
rect 29920 35702 29972 35708
rect 30196 35760 30248 35766
rect 30196 35702 30248 35708
rect 30300 35698 30328 36094
rect 30392 35834 30420 36790
rect 30840 36576 30892 36582
rect 30840 36518 30892 36524
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 29920 35556 29972 35562
rect 29920 35498 29972 35504
rect 29828 35148 29880 35154
rect 29828 35090 29880 35096
rect 29736 35012 29788 35018
rect 29736 34954 29788 34960
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29748 33998 29776 34546
rect 29932 34542 29960 35498
rect 30012 35080 30064 35086
rect 30012 35022 30064 35028
rect 30024 34746 30052 35022
rect 30104 35012 30156 35018
rect 30104 34954 30156 34960
rect 30012 34740 30064 34746
rect 30012 34682 30064 34688
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29552 33856 29604 33862
rect 29552 33798 29604 33804
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29472 32910 29500 33458
rect 29564 33318 29592 33798
rect 29932 33454 29960 34478
rect 30116 33998 30144 34954
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30288 33992 30340 33998
rect 30288 33934 30340 33940
rect 30024 33658 30052 33934
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 29920 33448 29972 33454
rect 29920 33390 29972 33396
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29656 33046 29684 33254
rect 29644 33040 29696 33046
rect 29644 32982 29696 32988
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29460 32904 29512 32910
rect 29460 32846 29512 32852
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 29460 32496 29512 32502
rect 29460 32438 29512 32444
rect 29472 22094 29500 32438
rect 29564 30734 29592 32710
rect 29748 32434 29776 32914
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29748 32026 29776 32370
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 29920 32360 29972 32366
rect 29920 32302 29972 32308
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 29840 31482 29868 32302
rect 29932 31958 29960 32302
rect 29920 31952 29972 31958
rect 29920 31894 29972 31900
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 29828 31476 29880 31482
rect 29828 31418 29880 31424
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 29644 31272 29696 31278
rect 29644 31214 29696 31220
rect 29656 30938 29684 31214
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29552 30728 29604 30734
rect 29552 30670 29604 30676
rect 29748 29730 29776 31282
rect 30116 30666 30144 31758
rect 30104 30660 30156 30666
rect 30104 30602 30156 30608
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 29656 29702 29776 29730
rect 29656 26024 29684 29702
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29748 28762 29776 29582
rect 29932 29238 29960 29786
rect 30024 29646 30052 30126
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 30208 29492 30236 29582
rect 30024 29464 30236 29492
rect 29920 29232 29972 29238
rect 29920 29174 29972 29180
rect 30024 29102 30052 29464
rect 30012 29096 30064 29102
rect 30012 29038 30064 29044
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 30024 28558 30052 29038
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 29656 25996 29776 26024
rect 29552 24608 29604 24614
rect 29552 24550 29604 24556
rect 29564 23186 29592 24550
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29552 23180 29604 23186
rect 29552 23122 29604 23128
rect 29656 23118 29684 24006
rect 29644 23112 29696 23118
rect 29644 23054 29696 23060
rect 29472 22066 29592 22094
rect 29564 21146 29592 22066
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29656 21554 29684 21966
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 29012 18850 29040 19382
rect 29656 19378 29684 19790
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 28920 18822 29040 18850
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28828 18426 28856 18702
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28816 18284 28868 18290
rect 28816 18226 28868 18232
rect 28828 17202 28856 18226
rect 28920 18222 28948 18822
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 28908 18216 28960 18222
rect 28908 18158 28960 18164
rect 29012 17338 29040 18702
rect 29656 18306 29684 19314
rect 29564 18278 29684 18306
rect 29564 18222 29592 18278
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29644 18148 29696 18154
rect 29644 18090 29696 18096
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29104 17678 29132 18022
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 28828 4146 28856 17138
rect 29012 17134 29040 17274
rect 29104 17202 29132 17614
rect 29184 17604 29236 17610
rect 29184 17546 29236 17552
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29196 17066 29224 17546
rect 29184 17060 29236 17066
rect 29184 17002 29236 17008
rect 29196 16658 29224 17002
rect 29564 16794 29592 17614
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29656 16658 29684 18090
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 28816 4140 28868 4146
rect 28816 4082 28868 4088
rect 29748 2774 29776 25996
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29840 21554 29868 22578
rect 29828 21548 29880 21554
rect 29828 21490 29880 21496
rect 29826 21448 29882 21457
rect 29826 21383 29828 21392
rect 29880 21383 29882 21392
rect 29828 21354 29880 21360
rect 29828 19780 29880 19786
rect 29828 19722 29880 19728
rect 29840 19446 29868 19722
rect 29828 19440 29880 19446
rect 29828 19382 29880 19388
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29840 17338 29868 17614
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29932 17218 29960 25230
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 30024 23769 30052 24142
rect 30010 23760 30066 23769
rect 30010 23695 30066 23704
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 30024 22234 30052 23462
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30116 22778 30144 23054
rect 30104 22772 30156 22778
rect 30104 22714 30156 22720
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 30196 21412 30248 21418
rect 30196 21354 30248 21360
rect 30208 21010 30236 21354
rect 30104 21004 30156 21010
rect 30104 20946 30156 20952
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30012 19848 30064 19854
rect 30012 19790 30064 19796
rect 30024 19514 30052 19790
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30024 18766 30052 19450
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 30116 17338 30144 20946
rect 30208 19990 30236 20946
rect 30196 19984 30248 19990
rect 30196 19926 30248 19932
rect 30196 18148 30248 18154
rect 30196 18090 30248 18096
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 29932 17190 30144 17218
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29932 15706 29960 15982
rect 29920 15700 29972 15706
rect 29920 15642 29972 15648
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 13938 29868 15438
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 30024 3466 30052 17070
rect 30116 5098 30144 17190
rect 30208 15502 30236 18090
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30104 5092 30156 5098
rect 30104 5034 30156 5040
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 30024 3126 30052 3402
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 29564 2746 29776 2774
rect 29564 2038 29592 2746
rect 30300 2650 30328 33934
rect 30392 32910 30420 35770
rect 30484 35630 30512 36110
rect 30472 35624 30524 35630
rect 30472 35566 30524 35572
rect 30484 35086 30512 35566
rect 30852 35494 30880 36518
rect 30944 36174 30972 37810
rect 31116 36848 31168 36854
rect 31116 36790 31168 36796
rect 31128 36378 31156 36790
rect 31116 36372 31168 36378
rect 31116 36314 31168 36320
rect 30932 36168 30984 36174
rect 30932 36110 30984 36116
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30484 33998 30512 35022
rect 30748 34400 30800 34406
rect 30748 34342 30800 34348
rect 30760 34066 30788 34342
rect 30748 34060 30800 34066
rect 30748 34002 30800 34008
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30944 32434 30972 36110
rect 31300 36100 31352 36106
rect 31300 36042 31352 36048
rect 31312 35834 31340 36042
rect 32324 35894 32352 36110
rect 32600 35894 32628 45358
rect 33232 37868 33284 37874
rect 33232 37810 33284 37816
rect 32680 37664 32732 37670
rect 32680 37606 32732 37612
rect 32692 37330 32720 37606
rect 32680 37324 32732 37330
rect 32680 37266 32732 37272
rect 33244 36922 33272 37810
rect 34704 37800 34756 37806
rect 34704 37742 34756 37748
rect 34716 37330 34744 37742
rect 34704 37324 34756 37330
rect 34704 37266 34756 37272
rect 33692 37188 33744 37194
rect 33692 37130 33744 37136
rect 33232 36916 33284 36922
rect 33232 36858 33284 36864
rect 33704 36378 33732 37130
rect 33968 37120 34020 37126
rect 33968 37062 34020 37068
rect 34704 37120 34756 37126
rect 34704 37062 34756 37068
rect 33980 36786 34008 37062
rect 34716 36922 34744 37062
rect 34704 36916 34756 36922
rect 34704 36858 34756 36864
rect 33968 36780 34020 36786
rect 33968 36722 34020 36728
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 32324 35866 32536 35894
rect 32600 35866 32720 35894
rect 31300 35828 31352 35834
rect 31300 35770 31352 35776
rect 31208 35080 31260 35086
rect 31208 35022 31260 35028
rect 31116 34604 31168 34610
rect 31116 34546 31168 34552
rect 31128 33930 31156 34546
rect 31116 33924 31168 33930
rect 31116 33866 31168 33872
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 31036 32978 31064 33526
rect 31128 33114 31156 33866
rect 31116 33108 31168 33114
rect 31116 33050 31168 33056
rect 31024 32972 31076 32978
rect 31024 32914 31076 32920
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 30748 32224 30800 32230
rect 30748 32166 30800 32172
rect 30380 31748 30432 31754
rect 30380 31690 30432 31696
rect 30392 31482 30420 31690
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30760 31346 30788 32166
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30656 31136 30708 31142
rect 30656 31078 30708 31084
rect 30668 29714 30696 31078
rect 30944 29850 30972 32370
rect 31220 31754 31248 35022
rect 32508 34610 32536 35866
rect 32588 35012 32640 35018
rect 32588 34954 32640 34960
rect 32600 34746 32628 34954
rect 32588 34740 32640 34746
rect 32588 34682 32640 34688
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 31300 33856 31352 33862
rect 31300 33798 31352 33804
rect 31312 32978 31340 33798
rect 31588 33386 31616 34546
rect 32508 33522 32536 34546
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 31576 33380 31628 33386
rect 31576 33322 31628 33328
rect 32404 33312 32456 33318
rect 32404 33254 32456 33260
rect 31300 32972 31352 32978
rect 31300 32914 31352 32920
rect 32416 32910 32444 33254
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 31392 32836 31444 32842
rect 31392 32778 31444 32784
rect 31404 32434 31432 32778
rect 31392 32428 31444 32434
rect 31392 32370 31444 32376
rect 31404 31890 31432 32370
rect 31484 32224 31536 32230
rect 31484 32166 31536 32172
rect 32036 32224 32088 32230
rect 32036 32166 32088 32172
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 31220 31726 31340 31754
rect 30932 29844 30984 29850
rect 30932 29786 30984 29792
rect 30656 29708 30708 29714
rect 30656 29650 30708 29656
rect 30944 28558 30972 29786
rect 31024 29232 31076 29238
rect 31024 29174 31076 29180
rect 31036 28762 31064 29174
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 30932 28552 30984 28558
rect 30932 28494 30984 28500
rect 30746 27568 30802 27577
rect 30746 27503 30802 27512
rect 30760 27470 30788 27503
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30944 26994 30972 28494
rect 31206 27024 31262 27033
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 31024 26988 31076 26994
rect 31206 26959 31208 26968
rect 31024 26930 31076 26936
rect 31260 26959 31262 26968
rect 31208 26930 31260 26936
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30932 26784 30984 26790
rect 30932 26726 30984 26732
rect 30392 25974 30420 26726
rect 30944 26314 30972 26726
rect 30932 26308 30984 26314
rect 30932 26250 30984 26256
rect 31036 26246 31064 26930
rect 31024 26240 31076 26246
rect 31024 26182 31076 26188
rect 30380 25968 30432 25974
rect 30380 25910 30432 25916
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30392 23322 30420 24142
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 30668 23186 30696 24006
rect 30656 23180 30708 23186
rect 30656 23122 30708 23128
rect 31208 21140 31260 21146
rect 31208 21082 31260 21088
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30944 19990 30972 20402
rect 30932 19984 30984 19990
rect 30932 19926 30984 19932
rect 31024 19236 31076 19242
rect 31024 19178 31076 19184
rect 31036 18834 31064 19178
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 30564 18760 30616 18766
rect 30564 18702 30616 18708
rect 30576 18358 30604 18702
rect 31024 18692 31076 18698
rect 31024 18634 31076 18640
rect 31036 18426 31064 18634
rect 31024 18420 31076 18426
rect 31024 18362 31076 18368
rect 30564 18352 30616 18358
rect 30564 18294 30616 18300
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30944 4146 30972 18226
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30380 3936 30432 3942
rect 30380 3878 30432 3884
rect 30392 3670 30420 3878
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 31220 2514 31248 21082
rect 31312 2854 31340 31726
rect 31404 31482 31432 31826
rect 31496 31822 31524 32166
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31392 31476 31444 31482
rect 31392 31418 31444 31424
rect 32048 31278 32076 32166
rect 32496 31952 32548 31958
rect 32496 31894 32548 31900
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 31760 31204 31812 31210
rect 31760 31146 31812 31152
rect 31484 30728 31536 30734
rect 31484 30670 31536 30676
rect 31496 29646 31524 30670
rect 31772 30598 31800 31146
rect 32048 30802 32076 31214
rect 32036 30796 32088 30802
rect 32036 30738 32088 30744
rect 32232 30666 32260 31282
rect 32404 31272 32456 31278
rect 32404 31214 32456 31220
rect 32220 30660 32272 30666
rect 32220 30602 32272 30608
rect 31760 30592 31812 30598
rect 31760 30534 31812 30540
rect 31484 29640 31536 29646
rect 31484 29582 31536 29588
rect 31772 28558 31800 30534
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31852 28416 31904 28422
rect 31852 28358 31904 28364
rect 31864 27538 31892 28358
rect 31576 27532 31628 27538
rect 31576 27474 31628 27480
rect 31852 27532 31904 27538
rect 31852 27474 31904 27480
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 31404 26790 31432 27270
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31588 25362 31616 27474
rect 31668 27464 31720 27470
rect 31668 27406 31720 27412
rect 31680 26586 31708 27406
rect 31668 26580 31720 26586
rect 31668 26522 31720 26528
rect 31680 25906 31708 26522
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31956 26042 31984 26250
rect 31944 26036 31996 26042
rect 31944 25978 31996 25984
rect 31668 25900 31720 25906
rect 31668 25842 31720 25848
rect 31576 25356 31628 25362
rect 31576 25298 31628 25304
rect 31680 24614 31708 25842
rect 32128 25220 32180 25226
rect 32128 25162 32180 25168
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 31680 24206 31708 24550
rect 31668 24200 31720 24206
rect 31668 24142 31720 24148
rect 31680 23730 31708 24142
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31668 23724 31720 23730
rect 31668 23666 31720 23672
rect 31772 23118 31800 24006
rect 32140 23322 32168 25162
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 32036 21616 32088 21622
rect 32036 21558 32088 21564
rect 32048 21146 32076 21558
rect 32128 21480 32180 21486
rect 32128 21422 32180 21428
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 32140 20466 32168 21422
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 31208 2508 31260 2514
rect 31208 2450 31260 2456
rect 29644 2440 29696 2446
rect 31404 2394 31432 15982
rect 32232 8838 32260 30602
rect 32416 29306 32444 31214
rect 32508 30122 32536 31894
rect 32496 30116 32548 30122
rect 32496 30058 32548 30064
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 32416 28626 32444 29242
rect 32508 29102 32536 30058
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32404 28620 32456 28626
rect 32404 28562 32456 28568
rect 32416 26450 32444 28562
rect 32588 28484 32640 28490
rect 32588 28426 32640 28432
rect 32600 28218 32628 28426
rect 32588 28212 32640 28218
rect 32588 28154 32640 28160
rect 32494 27024 32550 27033
rect 32494 26959 32496 26968
rect 32548 26959 32550 26968
rect 32496 26930 32548 26936
rect 32404 26444 32456 26450
rect 32404 26386 32456 26392
rect 32416 25906 32444 26386
rect 32508 26246 32536 26930
rect 32692 26586 32720 35866
rect 33980 35154 34008 36722
rect 34612 36712 34664 36718
rect 34612 36654 34664 36660
rect 34624 35290 34652 36654
rect 34612 35284 34664 35290
rect 34612 35226 34664 35232
rect 33968 35148 34020 35154
rect 33968 35090 34020 35096
rect 33508 34944 33560 34950
rect 33508 34886 33560 34892
rect 33520 34474 33548 34886
rect 33508 34468 33560 34474
rect 33508 34410 33560 34416
rect 33980 34406 34008 35090
rect 34060 35012 34112 35018
rect 34060 34954 34112 34960
rect 34072 34610 34100 34954
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 34060 34604 34112 34610
rect 34060 34546 34112 34552
rect 33968 34400 34020 34406
rect 33968 34342 34020 34348
rect 32864 34060 32916 34066
rect 32864 34002 32916 34008
rect 32772 33856 32824 33862
rect 32772 33798 32824 33804
rect 32784 33590 32812 33798
rect 32772 33584 32824 33590
rect 32772 33526 32824 33532
rect 32876 32570 32904 34002
rect 34532 33998 34560 34886
rect 34624 34746 34652 35226
rect 34808 35086 34836 45526
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35256 37324 35308 37330
rect 35256 37266 35308 37272
rect 35164 37120 35216 37126
rect 35164 37062 35216 37068
rect 35176 36922 35204 37062
rect 35268 36938 35296 37266
rect 35360 37262 35388 47126
rect 35440 45960 35492 45966
rect 35440 45902 35492 45908
rect 35348 37256 35400 37262
rect 35348 37198 35400 37204
rect 35164 36916 35216 36922
rect 35268 36910 35388 36938
rect 35164 36858 35216 36864
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 35360 35154 35388 36910
rect 35348 35148 35400 35154
rect 35348 35090 35400 35096
rect 34796 35080 34848 35086
rect 34796 35022 34848 35028
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 34612 34604 34664 34610
rect 34612 34546 34664 34552
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 34624 33998 34652 34546
rect 34808 33998 34836 34546
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 35164 33992 35216 33998
rect 35164 33934 35216 33940
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33060 32910 33088 33458
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 32864 32564 32916 32570
rect 32864 32506 32916 32512
rect 32876 31890 32904 32506
rect 32864 31884 32916 31890
rect 32864 31826 32916 31832
rect 32876 29714 32904 31826
rect 33060 30938 33088 32846
rect 33876 31272 33928 31278
rect 33876 31214 33928 31220
rect 33888 30938 33916 31214
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 34624 30258 34652 33934
rect 35176 33658 35204 33934
rect 35164 33652 35216 33658
rect 35164 33594 35216 33600
rect 34796 33516 34848 33522
rect 34796 33458 34848 33464
rect 34808 33114 34836 33458
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34796 31748 34848 31754
rect 34796 31690 34848 31696
rect 34704 31680 34756 31686
rect 34704 31622 34756 31628
rect 34716 30734 34744 31622
rect 34808 30938 34836 31690
rect 35348 31680 35400 31686
rect 35348 31622 35400 31628
rect 35360 31142 35388 31622
rect 35348 31136 35400 31142
rect 35348 31078 35400 31084
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34796 30932 34848 30938
rect 34796 30874 34848 30880
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 35164 30592 35216 30598
rect 35164 30534 35216 30540
rect 35176 30394 35204 30534
rect 35164 30388 35216 30394
rect 35164 30330 35216 30336
rect 34520 30252 34572 30258
rect 34520 30194 34572 30200
rect 34612 30252 34664 30258
rect 34612 30194 34664 30200
rect 34796 30252 34848 30258
rect 34796 30194 34848 30200
rect 32864 29708 32916 29714
rect 32864 29650 32916 29656
rect 32864 29572 32916 29578
rect 32864 29514 32916 29520
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32784 28082 32812 29446
rect 32876 29306 32904 29514
rect 34060 29504 34112 29510
rect 34060 29446 34112 29452
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 34072 29170 34100 29446
rect 34532 29306 34560 30194
rect 34520 29300 34572 29306
rect 34520 29242 34572 29248
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 34060 29164 34112 29170
rect 34060 29106 34112 29112
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32680 26580 32732 26586
rect 32680 26522 32732 26528
rect 32496 26240 32548 26246
rect 32496 26182 32548 26188
rect 32864 26240 32916 26246
rect 32864 26182 32916 26188
rect 32876 25974 32904 26182
rect 32864 25968 32916 25974
rect 32864 25910 32916 25916
rect 32404 25900 32456 25906
rect 32404 25842 32456 25848
rect 32588 21480 32640 21486
rect 32586 21448 32588 21457
rect 32640 21448 32642 21457
rect 32586 21383 32642 21392
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 32324 18358 32352 19110
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32968 12646 32996 29106
rect 33968 29096 34020 29102
rect 33968 29038 34020 29044
rect 33876 28620 33928 28626
rect 33876 28562 33928 28568
rect 33140 28484 33192 28490
rect 33140 28426 33192 28432
rect 33152 27606 33180 28426
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 33888 27470 33916 28562
rect 33980 27538 34008 29038
rect 34072 28762 34100 29106
rect 34808 28762 34836 30194
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35360 29102 35388 31078
rect 35348 29096 35400 29102
rect 35348 29038 35400 29044
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34060 28756 34112 28762
rect 34060 28698 34112 28704
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 35360 28558 35388 29038
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34704 28484 34756 28490
rect 34704 28426 34756 28432
rect 33968 27532 34020 27538
rect 33968 27474 34020 27480
rect 33876 27464 33928 27470
rect 33876 27406 33928 27412
rect 33888 27062 33916 27406
rect 33980 27130 34008 27474
rect 34716 27402 34744 28426
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 34060 27396 34112 27402
rect 34060 27338 34112 27344
rect 34704 27396 34756 27402
rect 34704 27338 34756 27344
rect 33968 27124 34020 27130
rect 33968 27066 34020 27072
rect 33876 27056 33928 27062
rect 33876 26998 33928 27004
rect 33968 26988 34020 26994
rect 34072 26976 34100 27338
rect 34020 26948 34100 26976
rect 34244 26988 34296 26994
rect 33968 26930 34020 26936
rect 34244 26930 34296 26936
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33336 26382 33364 26726
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33600 26308 33652 26314
rect 33600 26250 33652 26256
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33612 25498 33640 26250
rect 33796 25974 33824 26250
rect 34256 26246 34284 26930
rect 35360 26790 35388 27406
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26382 35388 26726
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34244 26240 34296 26246
rect 34244 26182 34296 26188
rect 34256 26042 34284 26182
rect 34244 26036 34296 26042
rect 34244 25978 34296 25984
rect 33784 25968 33836 25974
rect 33784 25910 33836 25916
rect 35360 25906 35388 26318
rect 35452 25974 35480 45902
rect 36176 45620 36228 45626
rect 36176 45562 36228 45568
rect 35808 35148 35860 35154
rect 35808 35090 35860 35096
rect 35624 34944 35676 34950
rect 35624 34886 35676 34892
rect 35636 34746 35664 34886
rect 35624 34740 35676 34746
rect 35624 34682 35676 34688
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35544 34202 35572 34546
rect 35532 34196 35584 34202
rect 35532 34138 35584 34144
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35728 31346 35756 32846
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 35820 30802 35848 35090
rect 35808 30796 35860 30802
rect 35808 30738 35860 30744
rect 36188 27538 36216 45562
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36832 31482 36860 31622
rect 36820 31476 36872 31482
rect 36820 31418 36872 31424
rect 36176 27532 36228 27538
rect 36176 27474 36228 27480
rect 36188 27334 36216 27474
rect 36176 27328 36228 27334
rect 36176 27270 36228 27276
rect 35532 26988 35584 26994
rect 35532 26930 35584 26936
rect 35440 25968 35492 25974
rect 35440 25910 35492 25916
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 35348 25900 35400 25906
rect 35348 25842 35400 25848
rect 33600 25492 33652 25498
rect 33600 25434 33652 25440
rect 34808 25294 34836 25842
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 33428 24954 33456 25230
rect 33600 25152 33652 25158
rect 33600 25094 33652 25100
rect 33416 24948 33468 24954
rect 33416 24890 33468 24896
rect 33612 24818 33640 25094
rect 33600 24812 33652 24818
rect 33600 24754 33652 24760
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33520 23050 33548 23666
rect 33508 23044 33560 23050
rect 33508 22986 33560 22992
rect 33140 20392 33192 20398
rect 33140 20334 33192 20340
rect 33152 19378 33180 20334
rect 33612 19854 33640 24754
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 34244 24744 34296 24750
rect 34244 24686 34296 24692
rect 33980 23254 34008 24686
rect 34256 24410 34284 24686
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34244 24404 34296 24410
rect 34244 24346 34296 24352
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 35084 23866 35112 24142
rect 35072 23860 35124 23866
rect 35072 23802 35124 23808
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 33968 23248 34020 23254
rect 33968 23190 34020 23196
rect 33980 23118 34008 23190
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 34152 20392 34204 20398
rect 34152 20334 34204 20340
rect 34164 19990 34192 20334
rect 34152 19984 34204 19990
rect 34152 19926 34204 19932
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33140 19236 33192 19242
rect 33140 19178 33192 19184
rect 33048 19168 33100 19174
rect 33048 19110 33100 19116
rect 33060 18834 33088 19110
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 33152 18766 33180 19178
rect 33612 19122 33640 19790
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33968 19712 34020 19718
rect 33968 19654 34020 19660
rect 33888 19446 33916 19654
rect 33876 19440 33928 19446
rect 33876 19382 33928 19388
rect 33980 19310 34008 19654
rect 33968 19304 34020 19310
rect 33968 19246 34020 19252
rect 33612 19094 33732 19122
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33612 17542 33640 18226
rect 33704 18222 33732 19094
rect 33980 18766 34008 19246
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 34164 18222 34192 19926
rect 34612 18692 34664 18698
rect 34612 18634 34664 18640
rect 34624 18358 34652 18634
rect 34612 18352 34664 18358
rect 34612 18294 34664 18300
rect 33692 18216 33744 18222
rect 33692 18158 33744 18164
rect 34152 18216 34204 18222
rect 34152 18158 34204 18164
rect 33600 17536 33652 17542
rect 33600 17478 33652 17484
rect 33612 17202 33640 17478
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33704 16590 33732 18158
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 33796 16794 33824 17070
rect 33784 16788 33836 16794
rect 33784 16730 33836 16736
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 34716 14278 34744 23734
rect 35452 23730 35480 25910
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35544 23050 35572 26930
rect 35900 25696 35952 25702
rect 35900 25638 35952 25644
rect 35912 25362 35940 25638
rect 35900 25356 35952 25362
rect 35900 25298 35952 25304
rect 36924 24206 36952 47194
rect 36912 24200 36964 24206
rect 36912 24142 36964 24148
rect 35808 24132 35860 24138
rect 35808 24074 35860 24080
rect 35820 23866 35848 24074
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35808 23724 35860 23730
rect 35808 23666 35860 23672
rect 35532 23044 35584 23050
rect 35532 22986 35584 22992
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34808 21146 34836 21286
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 35624 20936 35676 20942
rect 35624 20878 35676 20884
rect 34796 20868 34848 20874
rect 34796 20810 34848 20816
rect 34808 19990 34836 20810
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34796 19984 34848 19990
rect 34796 19926 34848 19932
rect 35636 19786 35664 20878
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35728 19922 35756 20334
rect 35716 19916 35768 19922
rect 35716 19858 35768 19864
rect 35624 19780 35676 19786
rect 35624 19722 35676 19728
rect 35532 19372 35584 19378
rect 35532 19314 35584 19320
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 32956 12640 33008 12646
rect 32956 12582 33008 12588
rect 34716 10674 34744 14214
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34704 10668 34756 10674
rect 34704 10610 34756 10616
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 32220 8832 32272 8838
rect 32220 8774 32272 8780
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35452 3602 35480 17070
rect 35544 3738 35572 19314
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 29644 2382 29696 2388
rect 29552 2032 29604 2038
rect 29552 1974 29604 1980
rect 28724 1964 28776 1970
rect 28724 1906 28776 1912
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 29656 800 29684 2382
rect 30944 2366 31432 2394
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29748 1902 29776 2246
rect 29736 1896 29788 1902
rect 29736 1838 29788 1844
rect 30944 800 30972 2366
rect 32232 800 32260 3062
rect 32968 2854 32996 3470
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33152 3126 33180 3334
rect 33796 3194 33824 3470
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35636 2650 35664 19722
rect 35820 17270 35848 23666
rect 37292 21962 37320 47382
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 37372 46980 37424 46986
rect 37372 46922 37424 46928
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 36372 20466 36400 20946
rect 36360 20460 36412 20466
rect 36360 20402 36412 20408
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 37292 19378 37320 20198
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37096 18760 37148 18766
rect 37096 18702 37148 18708
rect 37108 18630 37136 18702
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 37108 18154 37136 18566
rect 37096 18148 37148 18154
rect 37096 18090 37148 18096
rect 35808 17264 35860 17270
rect 35808 17206 35860 17212
rect 37384 5370 37412 46922
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 47122 39344 49200
rect 39304 47116 39356 47122
rect 39304 47058 39356 47064
rect 39304 46980 39356 46986
rect 39304 46922 39356 46928
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38304 46170 38332 46446
rect 38660 46368 38712 46374
rect 38660 46310 38712 46316
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38672 24818 38700 46310
rect 39212 40928 39264 40934
rect 39212 40870 39264 40876
rect 38660 24812 38712 24818
rect 38660 24754 38712 24760
rect 39224 23730 39252 40870
rect 39316 30734 39344 46922
rect 39960 46374 39988 49200
rect 41248 47462 41276 49200
rect 40040 47456 40092 47462
rect 40040 47398 40092 47404
rect 41236 47456 41288 47462
rect 41236 47398 41288 47404
rect 39948 46368 40000 46374
rect 39948 46310 40000 46316
rect 40052 35894 40080 47398
rect 41892 47240 41920 49200
rect 41892 47212 42012 47240
rect 41880 47048 41932 47054
rect 41880 46990 41932 46996
rect 41236 46368 41288 46374
rect 41236 46310 41288 46316
rect 41248 46034 41276 46310
rect 41236 46028 41288 46034
rect 41236 45970 41288 45976
rect 41420 45892 41472 45898
rect 41420 45834 41472 45840
rect 41432 45558 41460 45834
rect 41420 45552 41472 45558
rect 41420 45494 41472 45500
rect 41892 45490 41920 46990
rect 41984 46034 42012 47212
rect 42536 46442 42564 49200
rect 43076 46980 43128 46986
rect 43076 46922 43128 46928
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41972 46028 42024 46034
rect 41972 45970 42024 45976
rect 42628 45626 42656 46446
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 41052 45484 41104 45490
rect 41052 45426 41104 45432
rect 41880 45484 41932 45490
rect 41880 45426 41932 45432
rect 41064 44266 41092 45426
rect 42892 45416 42944 45422
rect 42892 45358 42944 45364
rect 42904 45082 42932 45358
rect 42892 45076 42944 45082
rect 42892 45018 42944 45024
rect 41052 44260 41104 44266
rect 41052 44202 41104 44208
rect 40052 35866 40264 35894
rect 39304 30728 39356 30734
rect 39304 30670 39356 30676
rect 40132 27532 40184 27538
rect 40132 27474 40184 27480
rect 40040 27396 40092 27402
rect 40040 27338 40092 27344
rect 40052 27130 40080 27338
rect 40040 27124 40092 27130
rect 40040 27066 40092 27072
rect 39856 26988 39908 26994
rect 39856 26930 39908 26936
rect 39868 26586 39896 26930
rect 39856 26580 39908 26586
rect 39856 26522 39908 26528
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 40040 23724 40092 23730
rect 40144 23712 40172 27474
rect 40236 24342 40264 35866
rect 40224 24336 40276 24342
rect 40224 24278 40276 24284
rect 41064 23798 41092 44202
rect 41696 32020 41748 32026
rect 41696 31962 41748 31968
rect 41052 23792 41104 23798
rect 41052 23734 41104 23740
rect 40092 23684 40172 23712
rect 40040 23666 40092 23672
rect 38384 23656 38436 23662
rect 38384 23598 38436 23604
rect 38292 19712 38344 19718
rect 38292 19654 38344 19660
rect 38304 19514 38332 19654
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 37464 19304 37516 19310
rect 37464 19246 37516 19252
rect 37476 18902 37504 19246
rect 37464 18896 37516 18902
rect 37464 18838 37516 18844
rect 38396 6914 38424 23598
rect 40040 23520 40092 23526
rect 40040 23462 40092 23468
rect 40052 23186 40080 23462
rect 40144 23186 40172 23684
rect 40224 23656 40276 23662
rect 40224 23598 40276 23604
rect 40040 23180 40092 23186
rect 40040 23122 40092 23128
rect 40132 23180 40184 23186
rect 40132 23122 40184 23128
rect 40236 22778 40264 23598
rect 41420 23520 41472 23526
rect 41420 23462 41472 23468
rect 41432 23118 41460 23462
rect 41420 23112 41472 23118
rect 41420 23054 41472 23060
rect 41604 22976 41656 22982
rect 41604 22918 41656 22924
rect 40224 22772 40276 22778
rect 40224 22714 40276 22720
rect 40224 22636 40276 22642
rect 40224 22578 40276 22584
rect 40038 22536 40094 22545
rect 40038 22471 40094 22480
rect 40052 22438 40080 22471
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 40052 22030 40080 22374
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40236 21962 40264 22578
rect 41616 22506 41644 22918
rect 41604 22500 41656 22506
rect 41604 22442 41656 22448
rect 41708 22098 41736 31962
rect 43088 31686 43116 46922
rect 43548 45554 43576 49286
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49314 46470 50000
rect 46124 49286 46470 49314
rect 43824 47054 43852 49200
rect 44468 47190 44496 49200
rect 44456 47184 44508 47190
rect 44456 47126 44508 47132
rect 43812 47048 43864 47054
rect 43812 46990 43864 46996
rect 44456 47048 44508 47054
rect 44456 46990 44508 46996
rect 43548 45526 44128 45554
rect 44100 45422 44128 45526
rect 44088 45416 44140 45422
rect 44088 45358 44140 45364
rect 44468 45082 44496 46990
rect 45112 46102 45140 49200
rect 45560 47932 45612 47938
rect 45560 47874 45612 47880
rect 45572 47410 45600 47874
rect 45480 47382 45600 47410
rect 45480 47002 45508 47382
rect 45376 46980 45428 46986
rect 45480 46974 45600 47002
rect 45376 46922 45428 46928
rect 45192 46504 45244 46510
rect 45192 46446 45244 46452
rect 45204 46170 45232 46446
rect 45192 46164 45244 46170
rect 45192 46106 45244 46112
rect 45100 46096 45152 46102
rect 45100 46038 45152 46044
rect 44916 45416 44968 45422
rect 44916 45358 44968 45364
rect 45192 45416 45244 45422
rect 45192 45358 45244 45364
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 44928 44402 44956 45358
rect 45204 45082 45232 45358
rect 45388 45082 45416 46922
rect 45572 45626 45600 46974
rect 45652 46096 45704 46102
rect 45652 46038 45704 46044
rect 45560 45620 45612 45626
rect 45560 45562 45612 45568
rect 45664 45554 45692 46038
rect 45756 45966 45784 49200
rect 46124 47938 46152 49286
rect 46358 49200 46470 49286
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 46112 47932 46164 47938
rect 46112 47874 46164 47880
rect 46754 47696 46810 47705
rect 46754 47631 46810 47640
rect 46768 46510 46796 47631
rect 46848 47252 46900 47258
rect 46848 47194 46900 47200
rect 46860 47025 46888 47194
rect 46846 47016 46902 47025
rect 46846 46951 46902 46960
rect 46756 46504 46808 46510
rect 46756 46446 46808 46452
rect 46664 46436 46716 46442
rect 46664 46378 46716 46384
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 46296 45892 46348 45898
rect 46296 45834 46348 45840
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 45664 45526 45784 45554
rect 45756 45422 45784 45526
rect 45744 45416 45796 45422
rect 45744 45358 45796 45364
rect 45192 45076 45244 45082
rect 45192 45018 45244 45024
rect 45376 45076 45428 45082
rect 45376 45018 45428 45024
rect 45560 44872 45612 44878
rect 45560 44814 45612 44820
rect 45744 44872 45796 44878
rect 45744 44814 45796 44820
rect 44916 44396 44968 44402
rect 44916 44338 44968 44344
rect 45572 38962 45600 44814
rect 45560 38956 45612 38962
rect 45560 38898 45612 38904
rect 45572 35894 45600 38898
rect 45572 35866 45692 35894
rect 43076 31680 43128 31686
rect 43076 31622 43128 31628
rect 45558 26616 45614 26625
rect 45558 26551 45614 26560
rect 45100 26240 45152 26246
rect 45100 26182 45152 26188
rect 45112 25974 45140 26182
rect 45100 25968 45152 25974
rect 45100 25910 45152 25916
rect 45100 25832 45152 25838
rect 45100 25774 45152 25780
rect 42892 24948 42944 24954
rect 42892 24890 42944 24896
rect 41880 23656 41932 23662
rect 41880 23598 41932 23604
rect 41892 22438 41920 23598
rect 42904 23594 42932 24890
rect 43076 24404 43128 24410
rect 43076 24346 43128 24352
rect 43444 24404 43496 24410
rect 43444 24346 43496 24352
rect 43088 24206 43116 24346
rect 43076 24200 43128 24206
rect 43076 24142 43128 24148
rect 43260 24200 43312 24206
rect 43260 24142 43312 24148
rect 43076 23792 43128 23798
rect 43076 23734 43128 23740
rect 42892 23588 42944 23594
rect 42892 23530 42944 23536
rect 43088 22778 43116 23734
rect 43168 23724 43220 23730
rect 43168 23666 43220 23672
rect 43076 22772 43128 22778
rect 43076 22714 43128 22720
rect 41880 22432 41932 22438
rect 41880 22374 41932 22380
rect 41696 22092 41748 22098
rect 41892 22094 41920 22374
rect 41696 22034 41748 22040
rect 41800 22066 41920 22094
rect 42536 22066 42840 22094
rect 40224 21956 40276 21962
rect 40224 21898 40276 21904
rect 40500 21956 40552 21962
rect 40500 21898 40552 21904
rect 40236 21350 40264 21898
rect 40224 21344 40276 21350
rect 40224 21286 40276 21292
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 39132 8294 39160 19314
rect 39120 8288 39172 8294
rect 39120 8230 39172 8236
rect 38304 6886 38424 6914
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37372 5364 37424 5370
rect 37372 5306 37424 5312
rect 37292 4978 37320 5306
rect 37384 5166 37412 5306
rect 37556 5296 37608 5302
rect 37556 5238 37608 5244
rect 37372 5160 37424 5166
rect 37372 5102 37424 5108
rect 37372 5024 37424 5030
rect 37292 4972 37372 4978
rect 37292 4966 37424 4972
rect 37292 4950 37412 4966
rect 37568 4282 37596 5238
rect 38304 5166 38332 6886
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 40040 5568 40092 5574
rect 40040 5510 40092 5516
rect 40052 5234 40080 5510
rect 40040 5228 40092 5234
rect 40040 5170 40092 5176
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 37556 4276 37608 4282
rect 37556 4218 37608 4224
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 37292 2922 37320 3538
rect 37752 3194 37780 4082
rect 38304 3602 38332 5102
rect 40144 4758 40172 5646
rect 40224 5160 40276 5166
rect 40224 5102 40276 5108
rect 40236 4826 40264 5102
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 40132 4752 40184 4758
rect 40132 4694 40184 4700
rect 40408 4616 40460 4622
rect 40408 4558 40460 4564
rect 40420 4282 40448 4558
rect 40408 4276 40460 4282
rect 40408 4218 40460 4224
rect 40512 4146 40540 21898
rect 41708 21554 41736 22034
rect 41696 21548 41748 21554
rect 41696 21490 41748 21496
rect 41708 20466 41736 21490
rect 41800 21434 41828 22066
rect 42536 22030 42564 22066
rect 42524 22024 42576 22030
rect 42524 21966 42576 21972
rect 42248 21956 42300 21962
rect 42248 21898 42300 21904
rect 42432 21956 42484 21962
rect 42432 21898 42484 21904
rect 41800 21406 41920 21434
rect 41696 20460 41748 20466
rect 41696 20402 41748 20408
rect 41892 18222 41920 21406
rect 42260 21350 42288 21898
rect 42340 21888 42392 21894
rect 42340 21830 42392 21836
rect 42248 21344 42300 21350
rect 42248 21286 42300 21292
rect 42352 20942 42380 21830
rect 42444 21690 42472 21898
rect 42432 21684 42484 21690
rect 42432 21626 42484 21632
rect 42536 21554 42564 21966
rect 42524 21548 42576 21554
rect 42524 21490 42576 21496
rect 42708 21548 42760 21554
rect 42708 21490 42760 21496
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 42720 20874 42748 21490
rect 42708 20868 42760 20874
rect 42708 20810 42760 20816
rect 42720 20330 42748 20810
rect 42812 20466 42840 22066
rect 43180 21690 43208 23666
rect 43272 23118 43300 24142
rect 43456 23118 43484 24346
rect 43904 24200 43956 24206
rect 43904 24142 43956 24148
rect 43916 23866 43944 24142
rect 43996 24064 44048 24070
rect 43996 24006 44048 24012
rect 43904 23860 43956 23866
rect 43904 23802 43956 23808
rect 43916 23254 43944 23802
rect 44008 23730 44036 24006
rect 43996 23724 44048 23730
rect 43996 23666 44048 23672
rect 43904 23248 43956 23254
rect 43904 23190 43956 23196
rect 43260 23112 43312 23118
rect 43260 23054 43312 23060
rect 43444 23112 43496 23118
rect 43444 23054 43496 23060
rect 44456 23112 44508 23118
rect 44456 23054 44508 23060
rect 43272 22574 43300 23054
rect 43456 22642 43484 23054
rect 44468 22778 44496 23054
rect 44456 22772 44508 22778
rect 44456 22714 44508 22720
rect 45112 22642 45140 25774
rect 45572 25226 45600 26551
rect 45560 25220 45612 25226
rect 45560 25162 45612 25168
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45572 23866 45600 24142
rect 45664 23882 45692 35866
rect 45756 24041 45784 44814
rect 46308 44402 46336 45834
rect 46492 44538 46520 45834
rect 46676 44538 46704 46378
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 47768 47184 47820 47190
rect 47768 47126 47820 47132
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47308 46368 47360 46374
rect 47308 46310 47360 46316
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46848 45348 46900 45354
rect 46848 45290 46900 45296
rect 46480 44532 46532 44538
rect 46480 44474 46532 44480
rect 46664 44532 46716 44538
rect 46664 44474 46716 44480
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46480 44192 46532 44198
rect 46480 44134 46532 44140
rect 46492 43858 46520 44134
rect 46480 43852 46532 43858
rect 46480 43794 46532 43800
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46860 41138 46888 45290
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46848 41132 46900 41138
rect 46848 41074 46900 41080
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 46388 38752 46440 38758
rect 46388 38694 46440 38700
rect 46572 38752 46624 38758
rect 46572 38694 46624 38700
rect 46400 38418 46428 38694
rect 46388 38412 46440 38418
rect 46388 38354 46440 38360
rect 46112 38344 46164 38350
rect 46112 38286 46164 38292
rect 45836 31816 45888 31822
rect 45836 31758 45888 31764
rect 45742 24032 45798 24041
rect 45742 23967 45798 23976
rect 45560 23860 45612 23866
rect 45664 23854 45784 23882
rect 45560 23802 45612 23808
rect 45652 23792 45704 23798
rect 45652 23734 45704 23740
rect 45560 23520 45612 23526
rect 45560 23462 45612 23468
rect 45284 23044 45336 23050
rect 45284 22986 45336 22992
rect 43444 22636 43496 22642
rect 43444 22578 43496 22584
rect 45100 22636 45152 22642
rect 45100 22578 45152 22584
rect 43260 22568 43312 22574
rect 43260 22510 43312 22516
rect 43720 22568 43772 22574
rect 43720 22510 43772 22516
rect 44180 22568 44232 22574
rect 44180 22510 44232 22516
rect 43168 21684 43220 21690
rect 43168 21626 43220 21632
rect 43260 21548 43312 21554
rect 43260 21490 43312 21496
rect 43272 20942 43300 21490
rect 43260 20936 43312 20942
rect 43260 20878 43312 20884
rect 43628 20936 43680 20942
rect 43628 20878 43680 20884
rect 42800 20460 42852 20466
rect 42800 20402 42852 20408
rect 43076 20460 43128 20466
rect 43076 20402 43128 20408
rect 42708 20324 42760 20330
rect 42708 20266 42760 20272
rect 42984 20324 43036 20330
rect 42984 20266 43036 20272
rect 42996 19854 43024 20266
rect 42984 19848 43036 19854
rect 42984 19790 43036 19796
rect 41880 18216 41932 18222
rect 41880 18158 41932 18164
rect 41892 5166 41920 18158
rect 42340 5296 42392 5302
rect 42340 5238 42392 5244
rect 41880 5160 41932 5166
rect 41880 5102 41932 5108
rect 40776 4616 40828 4622
rect 40776 4558 40828 4564
rect 40788 4214 40816 4558
rect 40776 4208 40828 4214
rect 40776 4150 40828 4156
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 40224 4072 40276 4078
rect 40276 4020 40356 4026
rect 40224 4014 40356 4020
rect 39408 3670 39436 4014
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 38292 3596 38344 3602
rect 38292 3538 38344 3544
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 38660 3460 38712 3466
rect 38660 3402 38712 3408
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 38672 3058 38700 3402
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 37280 2916 37332 2922
rect 37280 2858 37332 2864
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 37384 2446 37412 2790
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 35452 800 35480 2382
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 800 36124 2314
rect 38028 800 38056 2382
rect 38672 2310 38700 2994
rect 39132 2650 39160 3470
rect 39408 2990 39436 3606
rect 39592 3534 39620 4014
rect 40236 3998 40356 4014
rect 40328 3942 40356 3998
rect 40316 3936 40368 3942
rect 40316 3878 40368 3884
rect 40512 3738 40540 4082
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40500 3732 40552 3738
rect 40500 3674 40552 3680
rect 39580 3528 39632 3534
rect 39580 3470 39632 3476
rect 39764 3460 39816 3466
rect 39764 3402 39816 3408
rect 39776 3194 39804 3402
rect 39948 3392 40000 3398
rect 39948 3334 40000 3340
rect 39764 3188 39816 3194
rect 39764 3130 39816 3136
rect 39960 3058 39988 3334
rect 40788 3058 40816 4014
rect 41892 3602 41920 5102
rect 42352 4826 42380 5238
rect 42340 4820 42392 4826
rect 42340 4762 42392 4768
rect 42892 4616 42944 4622
rect 42892 4558 42944 4564
rect 41696 3596 41748 3602
rect 41696 3538 41748 3544
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 40972 3194 41000 3470
rect 40960 3188 41012 3194
rect 40960 3130 41012 3136
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 41708 2990 41736 3538
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42430 3360 42486 3369
rect 42430 3295 42486 3304
rect 39396 2984 39448 2990
rect 39396 2926 39448 2932
rect 41696 2984 41748 2990
rect 41696 2926 41748 2932
rect 41708 2650 41736 2926
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 41696 2644 41748 2650
rect 41696 2586 41748 2592
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 39396 2372 39448 2378
rect 39396 2314 39448 2320
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39408 1170 39436 2314
rect 39316 1142 39436 1170
rect 39316 800 39344 1142
rect 39960 800 39988 2382
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 42444 1714 42472 3295
rect 42720 3126 42748 3470
rect 42708 3120 42760 3126
rect 42708 3062 42760 3068
rect 42812 3058 42840 3538
rect 42800 3052 42852 3058
rect 42800 2994 42852 3000
rect 42904 2650 42932 4558
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42996 3126 43024 3334
rect 42984 3120 43036 3126
rect 42984 3062 43036 3068
rect 42524 2644 42576 2650
rect 42524 2586 42576 2592
rect 42892 2644 42944 2650
rect 42892 2586 42944 2592
rect 42536 1902 42564 2586
rect 43088 2582 43116 20402
rect 43168 20392 43220 20398
rect 43168 20334 43220 20340
rect 43180 19854 43208 20334
rect 43640 20058 43668 20878
rect 43628 20052 43680 20058
rect 43628 19994 43680 20000
rect 43168 19848 43220 19854
rect 43168 19790 43220 19796
rect 43628 19168 43680 19174
rect 43628 19110 43680 19116
rect 43640 18834 43668 19110
rect 43628 18828 43680 18834
rect 43628 18770 43680 18776
rect 43732 5166 43760 22510
rect 44192 21962 44220 22510
rect 44548 22024 44600 22030
rect 44548 21966 44600 21972
rect 44180 21956 44232 21962
rect 44180 21898 44232 21904
rect 44272 21956 44324 21962
rect 44272 21898 44324 21904
rect 43904 20800 43956 20806
rect 43904 20742 43956 20748
rect 43916 20398 43944 20742
rect 43904 20392 43956 20398
rect 43904 20334 43956 20340
rect 43812 20324 43864 20330
rect 43812 20266 43864 20272
rect 43824 19854 43852 20266
rect 43812 19848 43864 19854
rect 43812 19790 43864 19796
rect 43824 18766 43852 19790
rect 43916 19446 43944 20334
rect 44180 20256 44232 20262
rect 44180 20198 44232 20204
rect 43904 19440 43956 19446
rect 43904 19382 43956 19388
rect 44088 19304 44140 19310
rect 44088 19246 44140 19252
rect 43812 18760 43864 18766
rect 43812 18702 43864 18708
rect 44100 18698 44128 19246
rect 44192 18766 44220 20198
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 43720 5160 43772 5166
rect 43720 5102 43772 5108
rect 43732 4214 43760 5102
rect 43260 4208 43312 4214
rect 43260 4150 43312 4156
rect 43720 4208 43772 4214
rect 43720 4150 43772 4156
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 43076 2576 43128 2582
rect 43076 2518 43128 2524
rect 42524 1896 42576 1902
rect 42524 1838 42576 1844
rect 42444 1686 42564 1714
rect 42536 800 42564 1686
rect 43180 800 43208 2926
rect 43272 2514 43300 4150
rect 43720 4072 43772 4078
rect 43548 4020 43720 4026
rect 43548 4014 43772 4020
rect 43548 3998 43760 4014
rect 43548 3942 43576 3998
rect 43536 3936 43588 3942
rect 43536 3878 43588 3884
rect 44284 3670 44312 21898
rect 44560 21554 44588 21966
rect 44548 21548 44600 21554
rect 44548 21490 44600 21496
rect 45008 21480 45060 21486
rect 45008 21422 45060 21428
rect 45020 19854 45048 21422
rect 44548 19848 44600 19854
rect 44548 19790 44600 19796
rect 45008 19848 45060 19854
rect 45008 19790 45060 19796
rect 44560 19378 44588 19790
rect 44548 19372 44600 19378
rect 44548 19314 44600 19320
rect 44456 18420 44508 18426
rect 44456 18362 44508 18368
rect 44468 17678 44496 18362
rect 44560 17882 44588 19314
rect 45020 18630 45048 19790
rect 45112 19310 45140 22578
rect 45296 22030 45324 22986
rect 45572 22710 45600 23462
rect 45664 23186 45692 23734
rect 45652 23180 45704 23186
rect 45652 23122 45704 23128
rect 45560 22704 45612 22710
rect 45560 22646 45612 22652
rect 45560 22092 45612 22098
rect 45560 22034 45612 22040
rect 45284 22024 45336 22030
rect 45284 21966 45336 21972
rect 45376 21548 45428 21554
rect 45376 21490 45428 21496
rect 45388 20942 45416 21490
rect 45376 20936 45428 20942
rect 45376 20878 45428 20884
rect 45572 20534 45600 22034
rect 45756 21622 45784 23854
rect 45744 21616 45796 21622
rect 45744 21558 45796 21564
rect 45756 20874 45784 21558
rect 45744 20868 45796 20874
rect 45744 20810 45796 20816
rect 45560 20528 45612 20534
rect 45560 20470 45612 20476
rect 45652 19848 45704 19854
rect 45652 19790 45704 19796
rect 45100 19304 45152 19310
rect 45100 19246 45152 19252
rect 45192 18760 45244 18766
rect 45192 18702 45244 18708
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 45008 18624 45060 18630
rect 45008 18566 45060 18572
rect 44732 18284 44784 18290
rect 44732 18226 44784 18232
rect 44548 17876 44600 17882
rect 44548 17818 44600 17824
rect 44744 17814 44772 18226
rect 45204 18154 45232 18702
rect 45284 18624 45336 18630
rect 45284 18566 45336 18572
rect 45296 18290 45324 18566
rect 45284 18284 45336 18290
rect 45284 18226 45336 18232
rect 45192 18148 45244 18154
rect 45192 18090 45244 18096
rect 44732 17808 44784 17814
rect 44732 17750 44784 17756
rect 45204 17678 45232 18090
rect 45388 17746 45416 18702
rect 45664 18222 45692 19790
rect 45652 18216 45704 18222
rect 45652 18158 45704 18164
rect 45376 17740 45428 17746
rect 45376 17682 45428 17688
rect 44456 17672 44508 17678
rect 44456 17614 44508 17620
rect 45192 17672 45244 17678
rect 45192 17614 45244 17620
rect 45664 16726 45692 18158
rect 45652 16720 45704 16726
rect 45652 16662 45704 16668
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 45192 16516 45244 16522
rect 45192 16458 45244 16464
rect 45204 16250 45232 16458
rect 45192 16244 45244 16250
rect 45192 16186 45244 16192
rect 45480 16182 45508 16594
rect 45468 16176 45520 16182
rect 45468 16118 45520 16124
rect 45756 16114 45784 20810
rect 45744 16108 45796 16114
rect 45744 16050 45796 16056
rect 45560 16040 45612 16046
rect 45560 15982 45612 15988
rect 45572 15745 45600 15982
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45652 9580 45704 9586
rect 45652 9522 45704 9528
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 45664 3534 45692 9522
rect 45848 9450 45876 31758
rect 46018 31376 46074 31385
rect 46018 31311 46074 31320
rect 45928 24744 45980 24750
rect 45928 24686 45980 24692
rect 45940 21962 45968 24686
rect 46032 24274 46060 31311
rect 46020 24268 46072 24274
rect 46020 24210 46072 24216
rect 46018 24032 46074 24041
rect 46018 23967 46074 23976
rect 46032 21962 46060 23967
rect 46124 23798 46152 38286
rect 46296 37868 46348 37874
rect 46296 37810 46348 37816
rect 46308 26234 46336 37810
rect 46480 37664 46532 37670
rect 46480 37606 46532 37612
rect 46492 37330 46520 37606
rect 46480 37324 46532 37330
rect 46480 37266 46532 37272
rect 46480 32428 46532 32434
rect 46480 32370 46532 32376
rect 46216 26206 46336 26234
rect 46112 23792 46164 23798
rect 46112 23734 46164 23740
rect 46112 23656 46164 23662
rect 46112 23598 46164 23604
rect 45928 21956 45980 21962
rect 45928 21898 45980 21904
rect 46020 21956 46072 21962
rect 46020 21898 46072 21904
rect 45928 19508 45980 19514
rect 45928 19450 45980 19456
rect 45940 19242 45968 19450
rect 45928 19236 45980 19242
rect 45928 19178 45980 19184
rect 46032 18970 46060 21898
rect 46124 21865 46152 23598
rect 46110 21856 46166 21865
rect 46110 21791 46166 21800
rect 46216 21486 46244 26206
rect 46296 24812 46348 24818
rect 46296 24754 46348 24760
rect 46388 24812 46440 24818
rect 46388 24754 46440 24760
rect 46308 23905 46336 24754
rect 46294 23896 46350 23905
rect 46294 23831 46350 23840
rect 46400 23225 46428 24754
rect 46492 24750 46520 32370
rect 46480 24744 46532 24750
rect 46480 24686 46532 24692
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46386 23216 46442 23225
rect 46386 23151 46442 23160
rect 46584 22982 46612 38694
rect 46756 33516 46808 33522
rect 46756 33458 46808 33464
rect 46768 33425 46796 33458
rect 46754 33416 46810 33425
rect 46754 33351 46810 33360
rect 46756 31884 46808 31890
rect 46756 31826 46808 31832
rect 46768 29050 46796 31826
rect 46860 30138 46888 41074
rect 47032 40520 47084 40526
rect 47032 40462 47084 40468
rect 47044 39574 47072 40462
rect 47032 39568 47084 39574
rect 47032 39510 47084 39516
rect 47124 35488 47176 35494
rect 47124 35430 47176 35436
rect 47032 35080 47084 35086
rect 47032 35022 47084 35028
rect 46940 32836 46992 32842
rect 46940 32778 46992 32784
rect 46952 32570 46980 32778
rect 46940 32564 46992 32570
rect 46940 32506 46992 32512
rect 46860 30110 46980 30138
rect 46846 30016 46902 30025
rect 46846 29951 46902 29960
rect 46860 29850 46888 29951
rect 46848 29844 46900 29850
rect 46848 29786 46900 29792
rect 46952 29730 46980 30110
rect 46676 29022 46796 29050
rect 46860 29702 46980 29730
rect 46572 22976 46624 22982
rect 46572 22918 46624 22924
rect 46204 21480 46256 21486
rect 46204 21422 46256 21428
rect 46112 19780 46164 19786
rect 46112 19722 46164 19728
rect 46124 19446 46152 19722
rect 46112 19440 46164 19446
rect 46112 19382 46164 19388
rect 46020 18964 46072 18970
rect 46020 18906 46072 18912
rect 45926 18456 45982 18465
rect 45926 18391 45982 18400
rect 45940 18358 45968 18391
rect 45928 18352 45980 18358
rect 45928 18294 45980 18300
rect 45928 18216 45980 18222
rect 45928 18158 45980 18164
rect 45940 17610 45968 18158
rect 45928 17604 45980 17610
rect 45928 17546 45980 17552
rect 45836 9444 45888 9450
rect 45836 9386 45888 9392
rect 45744 8288 45796 8294
rect 45742 8256 45744 8265
rect 45796 8256 45798 8265
rect 45742 8191 45798 8200
rect 45940 7954 45968 17546
rect 46112 8492 46164 8498
rect 46112 8434 46164 8440
rect 45928 7948 45980 7954
rect 45928 7890 45980 7896
rect 45940 7274 45968 7890
rect 46124 7478 46152 8434
rect 46112 7472 46164 7478
rect 46112 7414 46164 7420
rect 46020 7336 46072 7342
rect 46020 7278 46072 7284
rect 45928 7268 45980 7274
rect 45928 7210 45980 7216
rect 46032 4146 46060 7278
rect 46124 4758 46152 7414
rect 46112 4752 46164 4758
rect 46112 4694 46164 4700
rect 46020 4140 46072 4146
rect 46020 4082 46072 4088
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 45204 3058 45232 3470
rect 46216 3466 46244 21422
rect 46480 20868 46532 20874
rect 46480 20810 46532 20816
rect 46492 20058 46520 20810
rect 46480 20052 46532 20058
rect 46480 19994 46532 20000
rect 46676 19990 46704 29022
rect 46860 26234 46888 29702
rect 46940 28552 46992 28558
rect 46940 28494 46992 28500
rect 46952 27606 46980 28494
rect 47044 28218 47072 35022
rect 47136 34066 47164 35430
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 47032 28212 47084 28218
rect 47032 28154 47084 28160
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 46768 26206 46888 26234
rect 46768 23322 46796 26206
rect 46846 25936 46902 25945
rect 46846 25871 46902 25880
rect 46860 25838 46888 25871
rect 46848 25832 46900 25838
rect 46848 25774 46900 25780
rect 46940 25220 46992 25226
rect 46940 25162 46992 25168
rect 46952 24818 46980 25162
rect 46848 24812 46900 24818
rect 46848 24754 46900 24760
rect 46940 24812 46992 24818
rect 46940 24754 46992 24760
rect 46756 23316 46808 23322
rect 46756 23258 46808 23264
rect 46860 22624 46888 24754
rect 46940 23180 46992 23186
rect 46940 23122 46992 23128
rect 46768 22596 46888 22624
rect 46768 21350 46796 22596
rect 46952 22574 46980 23122
rect 46940 22568 46992 22574
rect 46846 22536 46902 22545
rect 46940 22510 46992 22516
rect 46846 22471 46848 22480
rect 46900 22471 46902 22480
rect 46848 22442 46900 22448
rect 46952 22438 46980 22510
rect 46940 22432 46992 22438
rect 46940 22374 46992 22380
rect 46756 21344 46808 21350
rect 46756 21286 46808 21292
rect 46664 19984 46716 19990
rect 46664 19926 46716 19932
rect 46388 19372 46440 19378
rect 46388 19314 46440 19320
rect 46400 19174 46428 19314
rect 46388 19168 46440 19174
rect 46388 19110 46440 19116
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 16794 46336 17614
rect 46768 17218 46796 21286
rect 46952 20482 46980 22374
rect 47320 22094 47348 46310
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47492 44396 47544 44402
rect 47492 44338 47544 44344
rect 47400 44328 47452 44334
rect 47400 44270 47452 44276
rect 47412 43314 47440 44270
rect 47400 43308 47452 43314
rect 47400 43250 47452 43256
rect 47412 32434 47440 43250
rect 47504 35894 47532 44338
rect 47584 44260 47636 44266
rect 47584 44202 47636 44208
rect 47596 40050 47624 44202
rect 47688 43450 47716 44746
rect 47676 43444 47728 43450
rect 47676 43386 47728 43392
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47584 40044 47636 40050
rect 47584 39986 47636 39992
rect 47780 38706 47808 47126
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47964 46345 47992 46514
rect 47950 46336 48006 46345
rect 47950 46271 48006 46280
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48044 45280 48096 45286
rect 48044 45222 48096 45228
rect 47860 44736 47912 44742
rect 47860 44678 47912 44684
rect 47872 42226 47900 44678
rect 47860 42220 47912 42226
rect 47860 42162 47912 42168
rect 47872 40746 47900 42162
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47872 40718 47992 40746
rect 47860 38956 47912 38962
rect 47860 38898 47912 38904
rect 47872 38865 47900 38898
rect 47858 38856 47914 38865
rect 47858 38791 47914 38800
rect 47780 38678 47900 38706
rect 47768 37664 47820 37670
rect 47768 37606 47820 37612
rect 47780 37194 47808 37606
rect 47768 37188 47820 37194
rect 47768 37130 47820 37136
rect 47504 35866 47716 35894
rect 47584 34060 47636 34066
rect 47584 34002 47636 34008
rect 47492 33516 47544 33522
rect 47492 33458 47544 33464
rect 47400 32428 47452 32434
rect 47400 32370 47452 32376
rect 47504 31958 47532 33458
rect 47596 32026 47624 34002
rect 47584 32020 47636 32026
rect 47584 31962 47636 31968
rect 47492 31952 47544 31958
rect 47492 31894 47544 31900
rect 47596 31890 47624 31962
rect 47584 31884 47636 31890
rect 47584 31826 47636 31832
rect 47400 29504 47452 29510
rect 47400 29446 47452 29452
rect 47412 24138 47440 29446
rect 47688 28082 47716 35866
rect 47872 35086 47900 38678
rect 47860 35080 47912 35086
rect 47860 35022 47912 35028
rect 47860 34944 47912 34950
rect 47860 34886 47912 34892
rect 47768 34604 47820 34610
rect 47768 34546 47820 34552
rect 47780 33658 47808 34546
rect 47768 33652 47820 33658
rect 47768 33594 47820 33600
rect 47872 33318 47900 34886
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47964 32586 47992 40718
rect 48056 40610 48084 45222
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48134 41576 48190 41585
rect 48134 41511 48136 41520
rect 48188 41511 48190 41520
rect 48136 41482 48188 41488
rect 48056 40582 48268 40610
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48042 39536 48098 39545
rect 48148 39506 48176 40151
rect 48042 39471 48098 39480
rect 48136 39500 48188 39506
rect 48056 38418 48084 39471
rect 48136 39442 48188 39448
rect 48044 38412 48096 38418
rect 48044 38354 48096 38360
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48148 37330 48176 38111
rect 48136 37324 48188 37330
rect 48136 37266 48188 37272
rect 48136 35692 48188 35698
rect 48136 35634 48188 35640
rect 48044 35080 48096 35086
rect 48044 35022 48096 35028
rect 48056 34105 48084 35022
rect 48148 34785 48176 35634
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48042 34096 48098 34105
rect 48042 34031 48098 34040
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 47872 32558 47992 32586
rect 47676 28076 47728 28082
rect 47676 28018 47728 28024
rect 47688 27962 47716 28018
rect 47596 27934 47716 27962
rect 47596 27334 47624 27934
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27538 47716 27814
rect 47676 27532 47728 27538
rect 47676 27474 47728 27480
rect 47584 27328 47636 27334
rect 47584 27270 47636 27276
rect 47676 26376 47728 26382
rect 47676 26318 47728 26324
rect 47688 25362 47716 26318
rect 47872 26234 47900 32558
rect 47952 32428 48004 32434
rect 47952 32370 48004 32376
rect 47964 32065 47992 32370
rect 47950 32056 48006 32065
rect 47950 31991 48006 32000
rect 48136 29640 48188 29646
rect 48136 29582 48188 29588
rect 48148 29345 48176 29582
rect 48134 29336 48190 29345
rect 48134 29271 48190 29280
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 47872 26206 47992 26234
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47676 25356 47728 25362
rect 47676 25298 47728 25304
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47400 24132 47452 24138
rect 47400 24074 47452 24080
rect 47412 23526 47440 24074
rect 47400 23520 47452 23526
rect 47400 23462 47452 23468
rect 47136 22066 47348 22094
rect 47032 22024 47084 22030
rect 47032 21966 47084 21972
rect 47044 20602 47072 21966
rect 47032 20596 47084 20602
rect 47032 20538 47084 20544
rect 46952 20454 47072 20482
rect 47044 20398 47072 20454
rect 47032 20392 47084 20398
rect 47032 20334 47084 20340
rect 47044 19922 47072 20334
rect 47032 19916 47084 19922
rect 47032 19858 47084 19864
rect 47136 19514 47164 22066
rect 47412 21978 47440 23462
rect 47504 23050 47532 24754
rect 47584 24676 47636 24682
rect 47584 24618 47636 24624
rect 47492 23044 47544 23050
rect 47492 22986 47544 22992
rect 47228 21950 47440 21978
rect 47228 21622 47256 21950
rect 47504 21842 47532 22986
rect 47596 22642 47624 24618
rect 47780 24342 47808 25638
rect 47964 24818 47992 26206
rect 48134 25256 48190 25265
rect 48134 25191 48136 25200
rect 48188 25191 48190 25200
rect 48136 25162 48188 25168
rect 47952 24812 48004 24818
rect 47952 24754 48004 24760
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 47768 24336 47820 24342
rect 47768 24278 47820 24284
rect 48148 24274 48176 24511
rect 48240 24410 48268 40582
rect 48228 24404 48280 24410
rect 48228 24346 48280 24352
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 47676 24064 47728 24070
rect 47676 24006 47728 24012
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47320 21814 47532 21842
rect 47216 21616 47268 21622
rect 47216 21558 47268 21564
rect 47216 20800 47268 20806
rect 47216 20742 47268 20748
rect 47124 19508 47176 19514
rect 47124 19450 47176 19456
rect 46768 17190 46980 17218
rect 46664 17128 46716 17134
rect 46848 17128 46900 17134
rect 46664 17070 46716 17076
rect 46846 17096 46848 17105
rect 46900 17096 46902 17105
rect 46296 16788 46348 16794
rect 46296 16730 46348 16736
rect 46676 16522 46704 17070
rect 46756 17060 46808 17066
rect 46846 17031 46902 17040
rect 46756 17002 46808 17008
rect 46664 16516 46716 16522
rect 46664 16458 46716 16464
rect 46768 16114 46796 17002
rect 46952 16658 46980 17190
rect 46940 16652 46992 16658
rect 46940 16594 46992 16600
rect 46664 16108 46716 16114
rect 46664 16050 46716 16056
rect 46756 16108 46808 16114
rect 46756 16050 46808 16056
rect 46676 13938 46704 16050
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 46480 13728 46532 13734
rect 46480 13670 46532 13676
rect 46492 13394 46520 13670
rect 46480 13388 46532 13394
rect 46480 13330 46532 13336
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 46308 12850 46336 13262
rect 46296 12844 46348 12850
rect 46296 12786 46348 12792
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46940 9988 46992 9994
rect 46940 9930 46992 9936
rect 46952 9654 46980 9930
rect 46940 9648 46992 9654
rect 46940 9590 46992 9596
rect 46388 8288 46440 8294
rect 46388 8230 46440 8236
rect 46400 7886 46428 8230
rect 46388 7880 46440 7886
rect 46388 7822 46440 7828
rect 46940 7812 46992 7818
rect 46940 7754 46992 7760
rect 46952 7546 46980 7754
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 47228 6798 47256 20742
rect 47320 20210 47348 21814
rect 47596 21706 47624 22578
rect 47688 22438 47716 24006
rect 47952 23724 48004 23730
rect 47952 23666 48004 23672
rect 47860 22568 47912 22574
rect 47860 22510 47912 22516
rect 47676 22432 47728 22438
rect 47676 22374 47728 22380
rect 47504 21690 47624 21706
rect 47492 21684 47624 21690
rect 47544 21678 47624 21684
rect 47492 21626 47544 21632
rect 47504 20466 47532 21626
rect 47688 20534 47716 22374
rect 47872 21554 47900 22510
rect 47964 22094 47992 23666
rect 47964 22066 48084 22094
rect 48056 21554 48084 22066
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 48044 21548 48096 21554
rect 48044 21490 48096 21496
rect 47872 20806 47900 21490
rect 47860 20800 47912 20806
rect 47860 20742 47912 20748
rect 47676 20528 47728 20534
rect 47676 20470 47728 20476
rect 47492 20460 47544 20466
rect 47492 20402 47544 20408
rect 47952 20392 48004 20398
rect 47952 20334 48004 20340
rect 47320 20182 47532 20210
rect 47400 19168 47452 19174
rect 47400 19110 47452 19116
rect 47308 16584 47360 16590
rect 47308 16526 47360 16532
rect 47320 9586 47348 16526
rect 47308 9580 47360 9586
rect 47308 9522 47360 9528
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 47216 6792 47268 6798
rect 47216 6734 47268 6740
rect 46756 5228 46808 5234
rect 46756 5170 46808 5176
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 46308 3602 46336 3878
rect 46492 3602 46520 4422
rect 46664 4208 46716 4214
rect 46664 4150 46716 4156
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46676 3505 46704 4150
rect 46662 3496 46718 3505
rect 46204 3460 46256 3466
rect 46662 3431 46718 3440
rect 46204 3402 46256 3408
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45100 2916 45152 2922
rect 45100 2858 45152 2864
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 45112 800 45140 2858
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45480 1970 45508 2246
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 46400 800 46428 2314
rect 20180 734 20484 762
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 5170
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 46860 4185 46888 4558
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 47412 2514 47440 19110
rect 47504 18290 47532 20182
rect 47676 19372 47728 19378
rect 47676 19314 47728 19320
rect 47688 19174 47716 19314
rect 47768 19236 47820 19242
rect 47768 19178 47820 19184
rect 47676 19168 47728 19174
rect 47676 19110 47728 19116
rect 47780 18902 47808 19178
rect 47768 18896 47820 18902
rect 47768 18838 47820 18844
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47492 18284 47544 18290
rect 47492 18226 47544 18232
rect 47504 4690 47532 18226
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47688 17338 47716 17546
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 47676 11076 47728 11082
rect 47676 11018 47728 11024
rect 47688 10810 47716 11018
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 47492 4684 47544 4690
rect 47492 4626 47544 4632
rect 47780 3194 47808 18838
rect 47964 12434 47992 20334
rect 48056 19310 48084 21490
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 19304 48096 19310
rect 48044 19246 48096 19252
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 16425 48176 17546
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 47964 12406 48084 12434
rect 47858 9616 47914 9625
rect 47858 9551 47860 9560
rect 47912 9551 47914 9560
rect 47860 9522 47912 9528
rect 47860 8968 47912 8974
rect 47858 8936 47860 8945
rect 47912 8936 47914 8945
rect 47858 8871 47914 8880
rect 48056 6458 48084 12406
rect 48148 12345 48176 13194
rect 48134 12336 48190 12345
rect 48134 12271 48190 12280
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 48044 6452 48096 6458
rect 48044 6394 48096 6400
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 47964 6225 47992 6258
rect 47950 6216 48006 6225
rect 47950 6151 48006 6160
rect 47860 4208 47912 4214
rect 47860 4150 47912 4156
rect 47768 3188 47820 3194
rect 47768 3130 47820 3136
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47400 2508 47452 2514
rect 47400 2450 47452 2456
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47044 800 47072 2382
rect 47688 800 47716 2926
rect 47872 1465 47900 4150
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48320 3052 48372 3058
rect 48320 2994 48372 3000
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 47858 1456 47914 1465
rect 47858 1391 47914 1400
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48056 785 48084 2382
rect 48332 800 48360 2994
rect 48976 800 49004 3402
rect 48042 776 48098 785
rect 48042 711 48098 720
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 1398 42880 1454 42936
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1582 35400 1638 35456
rect 1582 32680 1638 32736
rect 1858 32000 1914 32056
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 1398 17720 1454 17776
rect 1858 16360 1914 16416
rect 1858 12280 1914 12336
rect 3422 46960 3478 47016
rect 2778 46280 2834 46336
rect 2318 27512 2374 27568
rect 2778 36760 2834 36816
rect 2410 22480 2466 22536
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3514 44920 3570 44976
rect 3698 43560 3754 43616
rect 3882 39480 3938 39536
rect 3882 31320 3938 31376
rect 3974 28620 4030 28656
rect 3974 28600 3976 28620
rect 3976 28600 4028 28620
rect 4028 28600 4030 28620
rect 3974 19760 4030 19816
rect 2226 19080 2282 19136
rect 3974 18400 4030 18456
rect 2778 15000 2834 15056
rect 3146 10240 3202 10296
rect 3514 17040 3570 17096
rect 3974 13676 3976 13696
rect 3976 13676 4028 13696
rect 4028 13676 4030 13696
rect 3974 13640 4030 13676
rect 3330 7520 3386 7576
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3422 3440 3478 3496
rect 3514 1400 3570 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 17590 23060 17592 23080
rect 17592 23060 17644 23080
rect 17644 23060 17646 23080
rect 17590 23024 17646 23060
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19338 3032 19394 3088
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 3440 19946 3496
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 2870 720 2926 776
rect 20626 3984 20682 4040
rect 22006 3304 22062 3360
rect 24674 3476 24676 3496
rect 24676 3476 24728 3496
rect 24728 3476 24730 3496
rect 24674 3440 24730 3476
rect 27986 32544 28042 32600
rect 26882 23160 26938 23216
rect 25778 22616 25834 22672
rect 25502 22344 25558 22400
rect 27066 22616 27122 22672
rect 27710 22616 27766 22672
rect 27894 22344 27950 22400
rect 25502 3984 25558 4040
rect 27342 3476 27344 3496
rect 27344 3476 27396 3496
rect 27396 3476 27398 3496
rect 27342 3440 27398 3476
rect 28998 32564 29054 32600
rect 28998 32544 29000 32564
rect 29000 32544 29052 32564
rect 29052 32544 29054 32564
rect 28998 23724 29054 23760
rect 28998 23704 29000 23724
rect 29000 23704 29052 23724
rect 29052 23704 29054 23724
rect 28722 23160 28778 23216
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 29826 21412 29882 21448
rect 29826 21392 29828 21412
rect 29828 21392 29880 21412
rect 29880 21392 29882 21412
rect 30010 23704 30066 23760
rect 30746 27512 30802 27568
rect 31206 26988 31262 27024
rect 31206 26968 31208 26988
rect 31208 26968 31260 26988
rect 31260 26968 31262 26988
rect 32494 26988 32550 27024
rect 32494 26968 32496 26988
rect 32496 26968 32548 26988
rect 32548 26968 32550 26988
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 32586 21428 32588 21448
rect 32588 21428 32640 21448
rect 32640 21428 32642 21448
rect 32586 21392 32642 21428
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40038 22480 40094 22536
rect 46754 47640 46810 47696
rect 46846 46960 46902 47016
rect 45558 26560 45614 26616
rect 45742 23976 45798 24032
rect 42430 3304 42486 3360
rect 45558 15680 45614 15736
rect 46018 31320 46074 31376
rect 46018 23976 46074 24032
rect 46110 21800 46166 21856
rect 46294 23840 46350 23896
rect 46386 23160 46442 23216
rect 46754 33360 46810 33416
rect 46846 29960 46902 30016
rect 45926 18400 45982 18456
rect 45742 8236 45744 8256
rect 45744 8236 45796 8256
rect 45796 8236 45798 8256
rect 45742 8200 45798 8236
rect 46846 25880 46902 25936
rect 46846 22500 46902 22536
rect 46846 22480 46848 22500
rect 46848 22480 46900 22500
rect 46900 22480 46902 22500
rect 47950 46280 48006 46336
rect 48134 45600 48190 45656
rect 47950 40840 48006 40896
rect 47858 38800 47914 38856
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41540 48190 41576
rect 48134 41520 48136 41540
rect 48136 41520 48188 41540
rect 48188 41520 48190 41540
rect 48134 40160 48190 40216
rect 48042 39480 48098 39536
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48042 34040 48098 34096
rect 48134 32680 48190 32736
rect 47950 32000 48006 32056
rect 48134 29280 48190 29336
rect 48134 27920 48190 27976
rect 48134 25220 48190 25256
rect 48134 25200 48136 25220
rect 48136 25200 48188 25220
rect 48188 25200 48190 25220
rect 48134 24520 48190 24576
rect 46846 17076 46848 17096
rect 46848 17076 46900 17096
rect 46900 17076 46902 17096
rect 46846 17040 46902 17076
rect 47306 7520 47362 7576
rect 46662 3440 46718 3496
rect 46846 4120 46902 4176
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 48134 16360 48190 16416
rect 47858 9580 47914 9616
rect 47858 9560 47860 9580
rect 47860 9560 47912 9580
rect 47912 9560 47914 9580
rect 47858 8916 47860 8936
rect 47860 8916 47912 8936
rect 47912 8916 47914 8936
rect 47858 8880 47914 8916
rect 48134 12280 48190 12336
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 47950 6160 48006 6216
rect 47858 1400 47914 1456
rect 46754 40 46810 96
rect 48042 720 48098 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 46749 47698 46815 47701
rect 49200 47698 50000 47788
rect 46749 47696 50000 47698
rect 46749 47640 46754 47696
rect 46810 47640 50000 47696
rect 46749 47638 50000 47640
rect 46749 47635 46815 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 46841 47018 46907 47021
rect 49200 47018 50000 47108
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3509 44978 3575 44981
rect 0 44976 3575 44978
rect 0 44920 3514 44976
rect 3570 44920 3575 44976
rect 0 44918 3575 44920
rect 0 44828 800 44918
rect 3509 44915 3575 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3693 43618 3759 43621
rect 0 43616 3759 43618
rect 0 43560 3698 43616
rect 3754 43560 3759 43616
rect 0 43558 3759 43560
rect 0 43468 800 43558
rect 3693 43555 3759 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3877 39538 3943 39541
rect 0 39536 3943 39538
rect 0 39480 3882 39536
rect 3938 39480 3943 39536
rect 0 39478 3943 39480
rect 0 39388 800 39478
rect 3877 39475 3943 39478
rect 48037 39538 48103 39541
rect 49200 39538 50000 39628
rect 48037 39536 50000 39538
rect 48037 39480 48042 39536
rect 48098 39480 50000 39536
rect 48037 39478 50000 39480
rect 48037 39475 48103 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47853 38858 47919 38861
rect 49200 38858 50000 38948
rect 47853 38856 50000 38858
rect 47853 38800 47858 38856
rect 47914 38800 50000 38856
rect 47853 38798 50000 38800
rect 47853 38795 47919 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48037 34098 48103 34101
rect 49200 34098 50000 34188
rect 48037 34096 50000 34098
rect 48037 34040 48042 34096
rect 48098 34040 50000 34096
rect 48037 34038 50000 34040
rect 48037 34035 48103 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 46749 33418 46815 33421
rect 49200 33418 50000 33508
rect 46749 33416 50000 33418
rect 46749 33360 46754 33416
rect 46810 33360 50000 33416
rect 46749 33358 50000 33360
rect 46749 33355 46815 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 27981 32602 28047 32605
rect 28993 32602 29059 32605
rect 27981 32600 29059 32602
rect 27981 32544 27986 32600
rect 28042 32544 28998 32600
rect 29054 32544 29059 32600
rect 49200 32588 50000 32678
rect 27981 32542 29059 32544
rect 27981 32539 28047 32542
rect 28993 32539 29059 32542
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 47945 32058 48011 32061
rect 49200 32058 50000 32148
rect 47945 32056 50000 32058
rect 47945 32000 47950 32056
rect 48006 32000 50000 32056
rect 47945 31998 50000 32000
rect 47945 31995 48011 31998
rect 49200 31908 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3877 31378 3943 31381
rect 0 31376 3943 31378
rect 0 31320 3882 31376
rect 3938 31320 3943 31376
rect 0 31318 3943 31320
rect 0 31228 800 31318
rect 3877 31315 3943 31318
rect 46013 31378 46079 31381
rect 49200 31378 50000 31468
rect 46013 31376 50000 31378
rect 46013 31320 46018 31376
rect 46074 31320 50000 31376
rect 46013 31318 50000 31320
rect 46013 31315 46079 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 46841 30018 46907 30021
rect 49200 30018 50000 30108
rect 46841 30016 50000 30018
rect 46841 29960 46846 30016
rect 46902 29960 50000 30016
rect 46841 29958 50000 29960
rect 46841 29955 46907 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 48129 29338 48195 29341
rect 49200 29338 50000 29428
rect 48129 29336 50000 29338
rect 48129 29280 48134 29336
rect 48190 29280 50000 29336
rect 48129 29278 50000 29280
rect 48129 29275 48195 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3969 28658 4035 28661
rect 0 28656 4035 28658
rect 0 28600 3974 28656
rect 4030 28600 4035 28656
rect 0 28598 4035 28600
rect 0 28508 800 28598
rect 3969 28595 4035 28598
rect 45686 28596 45692 28660
rect 45756 28658 45762 28660
rect 49200 28658 50000 28748
rect 45756 28598 50000 28658
rect 45756 28596 45762 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 2313 27570 2379 27573
rect 30741 27570 30807 27573
rect 2313 27568 30807 27570
rect 2313 27512 2318 27568
rect 2374 27512 30746 27568
rect 30802 27512 30807 27568
rect 2313 27510 30807 27512
rect 2313 27507 2379 27510
rect 30741 27507 30807 27510
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 31201 27026 31267 27029
rect 32489 27026 32555 27029
rect 31201 27024 32555 27026
rect 31201 26968 31206 27024
rect 31262 26968 32494 27024
rect 32550 26968 32555 27024
rect 31201 26966 32555 26968
rect 31201 26963 31267 26966
rect 32489 26963 32555 26966
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 45553 26618 45619 26621
rect 49200 26618 50000 26708
rect 45553 26616 50000 26618
rect 45553 26560 45558 26616
rect 45614 26560 50000 26616
rect 45553 26558 50000 26560
rect 45553 26555 45619 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46841 25938 46907 25941
rect 49200 25938 50000 26028
rect 46841 25936 50000 25938
rect 46841 25880 46846 25936
rect 46902 25880 50000 25936
rect 46841 25878 50000 25880
rect 46841 25875 46907 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25108 800 25198
rect 1853 25195 1919 25198
rect 48129 25258 48195 25261
rect 49200 25258 50000 25348
rect 48129 25256 50000 25258
rect 48129 25200 48134 25256
rect 48190 25200 50000 25256
rect 48129 25198 50000 25200
rect 48129 25195 48195 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 45737 24034 45803 24037
rect 46013 24034 46079 24037
rect 45737 24032 46079 24034
rect 0 23748 800 23988
rect 45737 23976 45742 24032
rect 45798 23976 46018 24032
rect 46074 23976 46079 24032
rect 45737 23974 46079 23976
rect 45737 23971 45803 23974
rect 46013 23971 46079 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46289 23898 46355 23901
rect 49200 23898 50000 23988
rect 46289 23896 50000 23898
rect 46289 23840 46294 23896
rect 46350 23840 50000 23896
rect 46289 23838 50000 23840
rect 46289 23835 46355 23838
rect 28993 23762 29059 23765
rect 30005 23762 30071 23765
rect 28993 23760 30071 23762
rect 28993 23704 28998 23760
rect 29054 23704 30010 23760
rect 30066 23704 30071 23760
rect 49200 23748 50000 23838
rect 28993 23702 30071 23704
rect 28993 23699 29059 23702
rect 30005 23699 30071 23702
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 26877 23218 26943 23221
rect 28717 23218 28783 23221
rect 26877 23216 28783 23218
rect 26877 23160 26882 23216
rect 26938 23160 28722 23216
rect 28778 23160 28783 23216
rect 26877 23158 28783 23160
rect 26877 23155 26943 23158
rect 28717 23155 28783 23158
rect 46381 23218 46447 23221
rect 49200 23218 50000 23308
rect 46381 23216 50000 23218
rect 46381 23160 46386 23216
rect 46442 23160 50000 23216
rect 46381 23158 50000 23160
rect 46381 23155 46447 23158
rect 17585 23082 17651 23085
rect 45318 23082 45324 23084
rect 17585 23080 45324 23082
rect 17585 23024 17590 23080
rect 17646 23024 45324 23080
rect 17585 23022 45324 23024
rect 17585 23019 17651 23022
rect 45318 23020 45324 23022
rect 45388 23020 45394 23084
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 25773 22674 25839 22677
rect 27061 22674 27127 22677
rect 27705 22674 27771 22677
rect 25773 22672 27771 22674
rect 0 22388 800 22628
rect 25773 22616 25778 22672
rect 25834 22616 27066 22672
rect 27122 22616 27710 22672
rect 27766 22616 27771 22672
rect 25773 22614 27771 22616
rect 25773 22611 25839 22614
rect 27061 22611 27127 22614
rect 27705 22611 27771 22614
rect 2405 22538 2471 22541
rect 40033 22538 40099 22541
rect 2405 22536 40099 22538
rect 2405 22480 2410 22536
rect 2466 22480 40038 22536
rect 40094 22480 40099 22536
rect 2405 22478 40099 22480
rect 2405 22475 2471 22478
rect 40033 22475 40099 22478
rect 46841 22538 46907 22541
rect 49200 22538 50000 22628
rect 46841 22536 50000 22538
rect 46841 22480 46846 22536
rect 46902 22480 50000 22536
rect 46841 22478 50000 22480
rect 46841 22475 46907 22478
rect 25497 22402 25563 22405
rect 27889 22402 27955 22405
rect 25497 22400 27955 22402
rect 25497 22344 25502 22400
rect 25558 22344 27894 22400
rect 27950 22344 27955 22400
rect 49200 22388 50000 22478
rect 25497 22342 27955 22344
rect 25497 22339 25563 22342
rect 27889 22339 27955 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 46105 21858 46171 21861
rect 49200 21858 50000 21948
rect 46105 21856 50000 21858
rect 46105 21800 46110 21856
rect 46166 21800 50000 21856
rect 46105 21798 50000 21800
rect 46105 21795 46171 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 29821 21450 29887 21453
rect 32581 21450 32647 21453
rect 29821 21448 32647 21450
rect 29821 21392 29826 21448
rect 29882 21392 32586 21448
rect 32642 21392 32647 21448
rect 29821 21390 32647 21392
rect 29821 21387 29887 21390
rect 32581 21387 32647 21390
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18308 800 18398
rect 3969 18395 4035 18398
rect 45921 18458 45987 18461
rect 49200 18458 50000 18548
rect 45921 18456 50000 18458
rect 45921 18400 45926 18456
rect 45982 18400 50000 18456
rect 45921 18398 50000 18400
rect 45921 18395 45987 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 16948 800 17038
rect 3509 17035 3575 17038
rect 46841 17098 46907 17101
rect 49200 17098 50000 17188
rect 46841 17096 50000 17098
rect 46841 17040 46846 17096
rect 46902 17040 50000 17096
rect 46841 17038 50000 17040
rect 46841 17035 46907 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1853 12338 1919 12341
rect 0 12336 1919 12338
rect 0 12280 1858 12336
rect 1914 12280 1919 12336
rect 0 12278 1919 12280
rect 0 12188 800 12278
rect 1853 12275 1919 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3141 10298 3207 10301
rect 0 10296 3207 10298
rect 0 10240 3146 10296
rect 3202 10240 3207 10296
rect 0 10238 3207 10240
rect 0 10148 800 10238
rect 3141 10235 3207 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 47853 9618 47919 9621
rect 49200 9618 50000 9708
rect 47853 9616 50000 9618
rect 47853 9560 47858 9616
rect 47914 9560 50000 9616
rect 47853 9558 50000 9560
rect 47853 9555 47919 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47853 8938 47919 8941
rect 49200 8938 50000 9028
rect 47853 8936 50000 8938
rect 47853 8880 47858 8936
rect 47914 8880 50000 8936
rect 47853 8878 50000 8880
rect 47853 8875 47919 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45737 8258 45803 8261
rect 49200 8258 50000 8348
rect 45737 8256 50000 8258
rect 45737 8200 45742 8256
rect 45798 8200 50000 8256
rect 45737 8198 50000 8200
rect 45737 8195 45803 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3325 7578 3391 7581
rect 0 7576 3391 7578
rect 0 7520 3330 7576
rect 3386 7520 3391 7576
rect 0 7518 3391 7520
rect 0 7428 800 7518
rect 3325 7515 3391 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 47945 6218 48011 6221
rect 49200 6218 50000 6308
rect 47945 6216 50000 6218
rect 47945 6160 47950 6216
rect 48006 6160 50000 6216
rect 47945 6158 50000 6160
rect 47945 6155 48011 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 20621 4042 20687 4045
rect 25497 4042 25563 4045
rect 20621 4040 25563 4042
rect 20621 3984 20626 4040
rect 20682 3984 25502 4040
rect 25558 3984 25563 4040
rect 49200 4028 50000 4118
rect 20621 3982 25563 3984
rect 20621 3979 20687 3982
rect 25497 3979 25563 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 19885 3498 19951 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 19382 3496 19951 3498
rect 19382 3440 19890 3496
rect 19946 3440 19951 3496
rect 19382 3438 19951 3440
rect 19382 3093 19442 3438
rect 19885 3435 19951 3438
rect 24669 3498 24735 3501
rect 27337 3498 27403 3501
rect 24669 3496 27403 3498
rect 24669 3440 24674 3496
rect 24730 3440 27342 3496
rect 27398 3440 27403 3496
rect 24669 3438 27403 3440
rect 24669 3435 24735 3438
rect 27337 3435 27403 3438
rect 46657 3498 46723 3501
rect 49200 3498 50000 3588
rect 46657 3496 50000 3498
rect 46657 3440 46662 3496
rect 46718 3440 50000 3496
rect 46657 3438 50000 3440
rect 46657 3435 46723 3438
rect 22001 3362 22067 3365
rect 42425 3362 42491 3365
rect 22001 3360 42491 3362
rect 22001 3304 22006 3360
rect 22062 3304 42430 3360
rect 42486 3304 42491 3360
rect 49200 3348 50000 3438
rect 22001 3302 42491 3304
rect 22001 3299 22067 3302
rect 42425 3299 42491 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 19333 3088 19442 3093
rect 19333 3032 19338 3088
rect 19394 3032 19442 3088
rect 19333 3030 19442 3032
rect 19333 3027 19399 3030
rect 0 2668 800 2908
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1308 800 1398
rect 3509 1395 3575 1398
rect 47853 1458 47919 1461
rect 49200 1458 50000 1548
rect 47853 1456 50000 1458
rect 47853 1400 47858 1456
rect 47914 1400 50000 1456
rect 47853 1398 50000 1400
rect 47853 1395 47919 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 48037 778 48103 781
rect 49200 778 50000 868
rect 48037 776 50000 778
rect 48037 720 48042 776
rect 48098 720 50000 776
rect 48037 718 50000 720
rect 48037 715 48103 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 45692 28596 45756 28660
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 45324 23020 45388 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 45691 28660 45757 28661
rect 45691 28596 45692 28660
rect 45756 28596 45757 28660
rect 45691 28595 45757 28596
rect 45694 28250 45754 28595
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 45326 28190 45754 28250
rect 45326 23085 45386 28190
rect 45323 23084 45389 23085
rect 45323 23020 45324 23084
rect 45388 23020 45389 23084
rect 45323 23019 45389 23020
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 24748 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 35420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 20056 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 29440 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 43792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 38640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 30912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_207
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1644511149
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_314
timestamp 1644511149
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1644511149
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_412
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_71
timestamp 1644511149
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_203
timestamp 1644511149
transform 1 0 19780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_210
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_216
timestamp 1644511149
transform 1 0 20976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_242
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_287
timestamp 1644511149
transform 1 0 27508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_299
timestamp 1644511149
transform 1 0 28612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_311
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_323
timestamp 1644511149
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1644511149
transform 1 0 35972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_399
timestamp 1644511149
transform 1 0 37812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_411
timestamp 1644511149
transform 1 0 38916 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_423
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_474
timestamp 1644511149
transform 1 0 44712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1644511149
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1644511149
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp 1644511149
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1644511149
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1644511149
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_278
timestamp 1644511149
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1644511149
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_409
timestamp 1644511149
transform 1 0 38732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_417
timestamp 1644511149
transform 1 0 39468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1644511149
transform 1 0 40572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1644511149
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_461
timestamp 1644511149
transform 1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_468
timestamp 1644511149
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_21
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1644511149
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_63
timestamp 1644511149
transform 1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_79
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_87
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_140
timestamp 1644511149
transform 1 0 13984 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1644511149
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_255
timestamp 1644511149
transform 1 0 24564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_313
timestamp 1644511149
transform 1 0 29900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1644511149
transform 1 0 30360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_396
timestamp 1644511149
transform 1 0 37536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_408
timestamp 1644511149
transform 1 0 38640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_433
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp 1644511149
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_464
timestamp 1644511149
transform 1 0 43792 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_476
timestamp 1644511149
transform 1 0 44896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_484
timestamp 1644511149
transform 1 0 45632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_490
timestamp 1644511149
transform 1 0 46184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_201
timestamp 1644511149
transform 1 0 19596 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1644511149
transform 1 0 20608 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_226
timestamp 1644511149
transform 1 0 21896 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1644511149
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_416
timestamp 1644511149
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_428
timestamp 1644511149
transform 1 0 40480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_435
timestamp 1644511149
transform 1 0 41124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_442
timestamp 1644511149
transform 1 0 41768 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_451
timestamp 1644511149
transform 1 0 42596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_463
timestamp 1644511149
transform 1 0 43700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1644511149
transform 1 0 46920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_204
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1644511149
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_236
timestamp 1644511149
transform 1 0 22816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_240
timestamp 1644511149
transform 1 0 23184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_244
timestamp 1644511149
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_256
timestamp 1644511149
transform 1 0 24656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_268
timestamp 1644511149
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_406
timestamp 1644511149
transform 1 0 38456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_410
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_422
timestamp 1644511149
transform 1 0 39928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_444
timestamp 1644511149
transform 1 0 41952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_462
timestamp 1644511149
transform 1 0 43608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_466
timestamp 1644511149
transform 1 0 43976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_478
timestamp 1644511149
transform 1 0 45080 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_490
timestamp 1644511149
transform 1 0 46184 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1644511149
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_428
timestamp 1644511149
transform 1 0 40480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_440
timestamp 1644511149
transform 1 0 41584 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_452
timestamp 1644511149
transform 1 0 42688 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_464
timestamp 1644511149
transform 1 0 43792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_500
timestamp 1644511149
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_493
timestamp 1644511149
transform 1 0 46460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_510
timestamp 1644511149
transform 1 0 48024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_487
timestamp 1644511149
transform 1 0 45908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_495
timestamp 1644511149
transform 1 0 46644 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1644511149
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_512
timestamp 1644511149
transform 1 0 48208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1644511149
transform 1 0 9016 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1644511149
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_284
timestamp 1644511149
transform 1 0 27232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_296
timestamp 1644511149
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_320
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_498
timestamp 1644511149
transform 1 0 46920 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_218
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1644511149
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1644511149
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_200
timestamp 1644511149
transform 1 0 19504 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_212
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_224
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_236
timestamp 1644511149
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1644511149
transform 1 0 30084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1644511149
transform 1 0 31188 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1644511149
transform 1 0 32292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1644511149
transform 1 0 33396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1644511149
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_477
timestamp 1644511149
transform 1 0 44988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_481
timestamp 1644511149
transform 1 0 45356 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_493
timestamp 1644511149
transform 1 0 46460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1644511149
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_235
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1644511149
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1644511149
transform 1 0 24840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_291
timestamp 1644511149
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1644511149
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1644511149
transform 1 0 29808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_348
timestamp 1644511149
transform 1 0 33120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_498
timestamp 1644511149
transform 1 0 46920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_505
timestamp 1644511149
transform 1 0 47564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_209
timestamp 1644511149
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_246
timestamp 1644511149
transform 1 0 23736 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1644511149
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_374
timestamp 1644511149
transform 1 0 35512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_386
timestamp 1644511149
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1644511149
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1644511149
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_322
timestamp 1644511149
transform 1 0 30728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_334
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_485
timestamp 1644511149
transform 1 0 45724 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_143
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_155
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1644511149
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_204
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_229
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_268
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1644511149
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_296
timestamp 1644511149
transform 1 0 28336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_306
timestamp 1644511149
transform 1 0 29256 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_315
timestamp 1644511149
transform 1 0 30084 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_323
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1644511149
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1644511149
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_383
timestamp 1644511149
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_465
timestamp 1644511149
transform 1 0 43884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_469
timestamp 1644511149
transform 1 0 44252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_486
timestamp 1644511149
transform 1 0 45816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_495
timestamp 1644511149
transform 1 0 46644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_166
timestamp 1644511149
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_179
timestamp 1644511149
transform 1 0 17572 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_200
timestamp 1644511149
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_211
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_258
timestamp 1644511149
transform 1 0 24840 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_266
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1644511149
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_318
timestamp 1644511149
transform 1 0 30360 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_341
timestamp 1644511149
transform 1 0 32476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1644511149
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_394
timestamp 1644511149
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_406
timestamp 1644511149
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1644511149
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_465
timestamp 1644511149
transform 1 0 43884 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_482
timestamp 1644511149
transform 1 0 45448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_490
timestamp 1644511149
transform 1 0 46184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_132
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_140
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_158
timestamp 1644511149
transform 1 0 15640 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_201
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_245
timestamp 1644511149
transform 1 0 23644 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_284
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_296
timestamp 1644511149
transform 1 0 28336 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_308
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_314
timestamp 1644511149
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_350
timestamp 1644511149
transform 1 0 33304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_375
timestamp 1644511149
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1644511149
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_414
timestamp 1644511149
transform 1 0 39192 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_426
timestamp 1644511149
transform 1 0 40296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_438
timestamp 1644511149
transform 1 0 41400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1644511149
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_457
timestamp 1644511149
transform 1 0 43148 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_463
timestamp 1644511149
transform 1 0 43700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_480
timestamp 1644511149
transform 1 0 45264 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1644511149
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_116
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_124
timestamp 1644511149
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_160
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1644511149
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_216
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_260
timestamp 1644511149
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_284
timestamp 1644511149
transform 1 0 27232 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_316
timestamp 1644511149
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_325
timestamp 1644511149
transform 1 0 31004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_337
timestamp 1644511149
transform 1 0 32108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_349
timestamp 1644511149
transform 1 0 33212 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1644511149
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_382
timestamp 1644511149
transform 1 0 36248 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_394
timestamp 1644511149
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_406
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1644511149
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_453
timestamp 1644511149
transform 1 0 42780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_458
timestamp 1644511149
transform 1 0 43240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_468
timestamp 1644511149
transform 1 0 44160 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_483
timestamp 1644511149
transform 1 0 45540 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_508
timestamp 1644511149
transform 1 0 47840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_116
timestamp 1644511149
transform 1 0 11776 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_127
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_212
timestamp 1644511149
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_236
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_260
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1644511149
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_285
timestamp 1644511149
transform 1 0 27324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_292
timestamp 1644511149
transform 1 0 27968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_304
timestamp 1644511149
transform 1 0 29072 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_316
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1644511149
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_377
timestamp 1644511149
transform 1 0 35788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1644511149
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_455
timestamp 1644511149
transform 1 0 42964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_467
timestamp 1644511149
transform 1 0 44068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_474
timestamp 1644511149
transform 1 0 44712 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_478
timestamp 1644511149
transform 1 0 45080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_510
timestamp 1644511149
transform 1 0 48024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_96
timestamp 1644511149
transform 1 0 9936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1644511149
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_123
timestamp 1644511149
transform 1 0 12420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1644511149
transform 1 0 13156 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_148
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_156
timestamp 1644511149
transform 1 0 15456 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_173
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1644511149
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1644511149
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_322
timestamp 1644511149
transform 1 0 30728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1644511149
transform 1 0 31648 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1644511149
transform 1 0 33396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_371
timestamp 1644511149
transform 1 0 35236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_375
timestamp 1644511149
transform 1 0 35604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_387
timestamp 1644511149
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_399
timestamp 1644511149
transform 1 0 37812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_411
timestamp 1644511149
transform 1 0 38916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_442
timestamp 1644511149
transform 1 0 41768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_449
timestamp 1644511149
transform 1 0 42412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_466
timestamp 1644511149
transform 1 0 43976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1644511149
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_91
timestamp 1644511149
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_98
timestamp 1644511149
transform 1 0 10120 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1644511149
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_180
timestamp 1644511149
transform 1 0 17664 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_192
timestamp 1644511149
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_228
timestamp 1644511149
transform 1 0 22080 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_232
timestamp 1644511149
transform 1 0 22448 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1644511149
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_271
timestamp 1644511149
transform 1 0 26036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_302
timestamp 1644511149
transform 1 0 28888 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_314
timestamp 1644511149
transform 1 0 29992 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_322
timestamp 1644511149
transform 1 0 30728 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_358
timestamp 1644511149
transform 1 0 34040 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_370
timestamp 1644511149
transform 1 0 35144 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_382
timestamp 1644511149
transform 1 0 36248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1644511149
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1644511149
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_459
timestamp 1644511149
transform 1 0 43332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_463
timestamp 1644511149
transform 1 0 43700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_468
timestamp 1644511149
transform 1 0 44160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_478
timestamp 1644511149
transform 1 0 45080 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_494
timestamp 1644511149
transform 1 0 46552 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1644511149
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1644511149
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_113
timestamp 1644511149
transform 1 0 11500 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1644511149
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1644511149
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_158
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_172
timestamp 1644511149
transform 1 0 16928 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_185
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_244
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_257
timestamp 1644511149
transform 1 0 24748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_269
timestamp 1644511149
transform 1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_276
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1644511149
transform 1 0 30084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1644511149
transform 1 0 31188 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1644511149
transform 1 0 33396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_427
timestamp 1644511149
transform 1 0 40388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_439
timestamp 1644511149
transform 1 0 41492 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_447
timestamp 1644511149
transform 1 0 42228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_455
timestamp 1644511149
transform 1 0 42964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_493
timestamp 1644511149
transform 1 0 46460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_507
timestamp 1644511149
transform 1 0 47748 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_515
timestamp 1644511149
transform 1 0 48484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_89
timestamp 1644511149
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_95
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1644511149
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_141
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_159
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1644511149
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_208
timestamp 1644511149
transform 1 0 20240 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_214
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1644511149
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_229
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_250
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1644511149
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_290
timestamp 1644511149
transform 1 0 27784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_302
timestamp 1644511149
transform 1 0 28888 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_307
timestamp 1644511149
transform 1 0 29348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_421
timestamp 1644511149
transform 1 0 39836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_428
timestamp 1644511149
transform 1 0 40480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_435
timestamp 1644511149
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_458
timestamp 1644511149
transform 1 0 43240 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_464
timestamp 1644511149
transform 1 0 43792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1644511149
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1644511149
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_110
timestamp 1644511149
transform 1 0 11224 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1644511149
transform 1 0 12696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_149
timestamp 1644511149
transform 1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_268
timestamp 1644511149
transform 1 0 25760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_272
timestamp 1644511149
transform 1 0 26128 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_294
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1644511149
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_314
timestamp 1644511149
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_338
timestamp 1644511149
transform 1 0 32200 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_346
timestamp 1644511149
transform 1 0 32936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_369
timestamp 1644511149
transform 1 0 35052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_393
timestamp 1644511149
transform 1 0 37260 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_405
timestamp 1644511149
transform 1 0 38364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1644511149
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_434
timestamp 1644511149
transform 1 0 41032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_444
timestamp 1644511149
transform 1 0 41952 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_454
timestamp 1644511149
transform 1 0 42872 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_461
timestamp 1644511149
transform 1 0 43516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1644511149
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_481
timestamp 1644511149
transform 1 0 45356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_506
timestamp 1644511149
transform 1 0 47656 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_514
timestamp 1644511149
transform 1 0 48392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1644511149
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 1644511149
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_151
timestamp 1644511149
transform 1 0 14996 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_176
timestamp 1644511149
transform 1 0 17296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_186
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_198
timestamp 1644511149
transform 1 0 19320 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_203
timestamp 1644511149
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_241
timestamp 1644511149
transform 1 0 23276 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_263
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1644511149
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_291
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_295
timestamp 1644511149
transform 1 0 28244 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_306
timestamp 1644511149
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_310
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_340
timestamp 1644511149
transform 1 0 32384 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_372
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1644511149
transform 1 0 35972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_411
timestamp 1644511149
transform 1 0 38916 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1644511149
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1644511149
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_453
timestamp 1644511149
transform 1 0 42780 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_479
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_486
timestamp 1644511149
transform 1 0 45816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_511
timestamp 1644511149
transform 1 0 48116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_515
timestamp 1644511149
transform 1 0 48484 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1644511149
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_106
timestamp 1644511149
transform 1 0 10856 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1644511149
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_122
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1644511149
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_162
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_187
timestamp 1644511149
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_220
timestamp 1644511149
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1644511149
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_313
timestamp 1644511149
transform 1 0 29900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_320
timestamp 1644511149
transform 1 0 30544 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_335
timestamp 1644511149
transform 1 0 31924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_347
timestamp 1644511149
transform 1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_351
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_355
timestamp 1644511149
transform 1 0 33764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_390
timestamp 1644511149
transform 1 0 36984 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_402
timestamp 1644511149
transform 1 0 38088 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1644511149
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_453
timestamp 1644511149
transform 1 0 42780 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_461
timestamp 1644511149
transform 1 0 43516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_468
timestamp 1644511149
transform 1 0 44160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_483
timestamp 1644511149
transform 1 0 45540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1644511149
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_144
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_154
timestamp 1644511149
transform 1 0 15272 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1644511149
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_209
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_302
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_326
timestamp 1644511149
transform 1 0 31096 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1644511149
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_356
timestamp 1644511149
transform 1 0 33856 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1644511149
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_489
timestamp 1644511149
transform 1 0 46092 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_493
timestamp 1644511149
transform 1 0 46460 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1644511149
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_118
timestamp 1644511149
transform 1 0 11960 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_126
timestamp 1644511149
transform 1 0 12696 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_145
timestamp 1644511149
transform 1 0 14444 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_182
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_188
timestamp 1644511149
transform 1 0 18400 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_218
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_222
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1644511149
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1644511149
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_275
timestamp 1644511149
transform 1 0 26404 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_326
timestamp 1644511149
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_338
timestamp 1644511149
transform 1 0 32200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1644511149
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1644511149
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_372
timestamp 1644511149
transform 1 0 35328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_397
timestamp 1644511149
transform 1 0 37628 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_409
timestamp 1644511149
transform 1 0 38732 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1644511149
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_73
timestamp 1644511149
transform 1 0 7820 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_95
timestamp 1644511149
transform 1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1644511149
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_116
timestamp 1644511149
transform 1 0 11776 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_128
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_140
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_146
timestamp 1644511149
transform 1 0 14536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_151
timestamp 1644511149
transform 1 0 14996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_184
timestamp 1644511149
transform 1 0 18032 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_192
timestamp 1644511149
transform 1 0 18768 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_209
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1644511149
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_244
timestamp 1644511149
transform 1 0 23552 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_289
timestamp 1644511149
transform 1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_318
timestamp 1644511149
transform 1 0 30360 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_326
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_369
timestamp 1644511149
transform 1 0 35052 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_377
timestamp 1644511149
transform 1 0 35788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_384
timestamp 1644511149
transform 1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_477
timestamp 1644511149
transform 1 0 44988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_499
timestamp 1644511149
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1644511149
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_92
timestamp 1644511149
transform 1 0 9568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_101
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_116
timestamp 1644511149
transform 1 0 11776 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_128
timestamp 1644511149
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_132
timestamp 1644511149
transform 1 0 13248 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_162
timestamp 1644511149
transform 1 0 16008 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_257
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_264
timestamp 1644511149
transform 1 0 25392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_272
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_282
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_352
timestamp 1644511149
transform 1 0 33488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1644511149
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_371
timestamp 1644511149
transform 1 0 35236 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_378
timestamp 1644511149
transform 1 0 35880 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_390
timestamp 1644511149
transform 1 0 36984 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_402
timestamp 1644511149
transform 1 0 38088 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_414
timestamp 1644511149
transform 1 0 39192 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_480
timestamp 1644511149
transform 1 0 45264 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_492
timestamp 1644511149
transform 1 0 46368 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_515
timestamp 1644511149
transform 1 0 48484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1644511149
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_94
timestamp 1644511149
transform 1 0 9752 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_123
timestamp 1644511149
transform 1 0 12420 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_190
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_202
timestamp 1644511149
transform 1 0 19688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1644511149
transform 1 0 23460 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_313
timestamp 1644511149
transform 1 0 29900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_320
timestamp 1644511149
transform 1 0 30544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1644511149
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_340
timestamp 1644511149
transform 1 0 32384 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_348
timestamp 1644511149
transform 1 0 33120 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_353
timestamp 1644511149
transform 1 0 33580 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_374
timestamp 1644511149
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1644511149
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_424
timestamp 1644511149
transform 1 0 40112 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_436
timestamp 1644511149
transform 1 0 41216 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_176
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_182
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1644511149
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_223
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_231
timestamp 1644511149
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_256
timestamp 1644511149
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_267
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_276
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1644511149
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_349
timestamp 1644511149
transform 1 0 33212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_358
timestamp 1644511149
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_371
timestamp 1644511149
transform 1 0 35236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1644511149
transform 1 0 36432 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1644511149
transform 1 0 37536 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1644511149
transform 1 0 38640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_442
timestamp 1644511149
transform 1 0 41768 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_454
timestamp 1644511149
transform 1 0 42872 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_466
timestamp 1644511149
transform 1 0 43976 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1644511149
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_75
timestamp 1644511149
transform 1 0 8004 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_80
timestamp 1644511149
transform 1 0 8464 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_88
timestamp 1644511149
transform 1 0 9200 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1644511149
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_99
timestamp 1644511149
transform 1 0 10212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1644511149
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_130
timestamp 1644511149
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_178
timestamp 1644511149
transform 1 0 17480 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_189
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_254
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_259
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_291
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_302
timestamp 1644511149
transform 1 0 28888 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_314
timestamp 1644511149
transform 1 0 29992 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_326
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1644511149
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_341
timestamp 1644511149
transform 1 0 32476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_345
timestamp 1644511149
transform 1 0 32844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_357
timestamp 1644511149
transform 1 0 33948 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_369
timestamp 1644511149
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1644511149
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_110
timestamp 1644511149
transform 1 0 11224 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_126
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1644511149
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_149
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1644511149
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_205
timestamp 1644511149
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_212
timestamp 1644511149
transform 1 0 20608 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_225
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_256
timestamp 1644511149
transform 1 0 24656 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_285
timestamp 1644511149
transform 1 0 27324 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_296
timestamp 1644511149
transform 1 0 28336 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_300
timestamp 1644511149
transform 1 0 28704 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_316
timestamp 1644511149
transform 1 0 30176 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_322
timestamp 1644511149
transform 1 0 30728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_326
timestamp 1644511149
transform 1 0 31096 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_336
timestamp 1644511149
transform 1 0 32016 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1644511149
transform 1 0 35328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1644511149
transform 1 0 36432 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_396
timestamp 1644511149
transform 1 0 37536 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_408
timestamp 1644511149
transform 1 0 38640 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_507
timestamp 1644511149
transform 1 0 47748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_515
timestamp 1644511149
transform 1 0 48484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_87
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_91
timestamp 1644511149
transform 1 0 9476 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_103
timestamp 1644511149
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_122
timestamp 1644511149
transform 1 0 12328 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_133
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_141
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_184
timestamp 1644511149
transform 1 0 18032 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_192
timestamp 1644511149
transform 1 0 18768 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_199
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_211
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_231
timestamp 1644511149
transform 1 0 22356 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_251
timestamp 1644511149
transform 1 0 24196 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_263
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1644511149
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_298
timestamp 1644511149
transform 1 0 28520 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_307
timestamp 1644511149
transform 1 0 29348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_352
timestamp 1644511149
transform 1 0 33488 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_363
timestamp 1644511149
transform 1 0 34500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_371
timestamp 1644511149
transform 1 0 35236 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_383
timestamp 1644511149
transform 1 0 36340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_110
timestamp 1644511149
transform 1 0 11224 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_116
timestamp 1644511149
transform 1 0 11776 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1644511149
transform 1 0 12604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1644511149
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_145
timestamp 1644511149
transform 1 0 14444 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_173
timestamp 1644511149
transform 1 0 17020 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1644511149
transform 1 0 17664 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_201
timestamp 1644511149
transform 1 0 19596 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_208
timestamp 1644511149
transform 1 0 20240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1644511149
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_230
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_237
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_256
timestamp 1644511149
transform 1 0 24656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_268
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_278
timestamp 1644511149
transform 1 0 26680 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_287
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_326
timestamp 1644511149
transform 1 0 31096 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_338
timestamp 1644511149
transform 1 0 32200 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_342
timestamp 1644511149
transform 1 0 32568 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_352
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_89
timestamp 1644511149
transform 1 0 9292 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_95
timestamp 1644511149
transform 1 0 9844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1644511149
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1644511149
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_119
timestamp 1644511149
transform 1 0 12052 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_140
timestamp 1644511149
transform 1 0 13984 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_146
timestamp 1644511149
transform 1 0 14536 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_154
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1644511149
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1644511149
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_233
timestamp 1644511149
transform 1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_262
timestamp 1644511149
transform 1 0 25208 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1644511149
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_289
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_303
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_308
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_320
timestamp 1644511149
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_366
timestamp 1644511149
transform 1 0 34776 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_378
timestamp 1644511149
transform 1 0 35880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 1644511149
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_125
timestamp 1644511149
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1644511149
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_147
timestamp 1644511149
transform 1 0 14628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_152
timestamp 1644511149
transform 1 0 15088 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_164
timestamp 1644511149
transform 1 0 16192 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_186
timestamp 1644511149
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_204
timestamp 1644511149
transform 1 0 19872 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_211
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_223
timestamp 1644511149
transform 1 0 21620 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_235
timestamp 1644511149
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_241
timestamp 1644511149
transform 1 0 23276 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_276
timestamp 1644511149
transform 1 0 26496 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_280
timestamp 1644511149
transform 1 0 26864 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_287
timestamp 1644511149
transform 1 0 27508 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1644511149
transform 1 0 29808 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_324
timestamp 1644511149
transform 1 0 30912 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_334
timestamp 1644511149
transform 1 0 31832 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_359
timestamp 1644511149
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_374
timestamp 1644511149
transform 1 0 35512 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_386
timestamp 1644511149
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_398
timestamp 1644511149
transform 1 0 37720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_410
timestamp 1644511149
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 1644511149
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_26
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_130
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_142
timestamp 1644511149
transform 1 0 14168 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1644511149
transform 1 0 14996 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1644511149
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_175
timestamp 1644511149
transform 1 0 17204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1644511149
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_203
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_215
timestamp 1644511149
transform 1 0 20884 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_233
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_290
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_298
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_303
timestamp 1644511149
transform 1 0 28980 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_316
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_323
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1644511149
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_342
timestamp 1644511149
transform 1 0 32568 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_350
timestamp 1644511149
transform 1 0 33304 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_372
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_50
timestamp 1644511149
transform 1 0 5704 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_62
timestamp 1644511149
transform 1 0 6808 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_74
timestamp 1644511149
transform 1 0 7912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1644511149
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_200
timestamp 1644511149
transform 1 0 19504 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_208
timestamp 1644511149
transform 1 0 20240 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_215
timestamp 1644511149
transform 1 0 20884 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_223
timestamp 1644511149
transform 1 0 21620 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1644511149
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1644511149
transform 1 0 25944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_288
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_296
timestamp 1644511149
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_335
timestamp 1644511149
transform 1 0 31924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_355
timestamp 1644511149
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_374
timestamp 1644511149
transform 1 0 35512 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_386
timestamp 1644511149
transform 1 0 36616 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_410
timestamp 1644511149
transform 1 0 38824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1644511149
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_508
timestamp 1644511149
transform 1 0 47840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_212
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1644511149
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_255
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_285
timestamp 1644511149
transform 1 0 27324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_290
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_303
timestamp 1644511149
transform 1 0 28980 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_316
timestamp 1644511149
transform 1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_324
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1644511149
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_341
timestamp 1644511149
transform 1 0 32476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_353
timestamp 1644511149
transform 1 0 33580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_365
timestamp 1644511149
transform 1 0 34684 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_377
timestamp 1644511149
transform 1 0 35788 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1644511149
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_512
timestamp 1644511149
transform 1 0 48208 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_14
timestamp 1644511149
transform 1 0 2392 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1644511149
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_207
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_218
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_227
timestamp 1644511149
transform 1 0 21988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_257
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_267
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_290
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_296
timestamp 1644511149
transform 1 0 28336 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1644511149
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_313
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_368
timestamp 1644511149
transform 1 0 34960 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_380
timestamp 1644511149
transform 1 0 36064 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_392
timestamp 1644511149
transform 1 0 37168 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_404
timestamp 1644511149
transform 1 0 38272 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_416
timestamp 1644511149
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_483
timestamp 1644511149
transform 1 0 45540 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_487
timestamp 1644511149
transform 1 0 45908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_215
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_239
timestamp 1644511149
transform 1 0 23092 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_289
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_297
timestamp 1644511149
transform 1 0 28428 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_304
timestamp 1644511149
transform 1 0 29072 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_327
timestamp 1644511149
transform 1 0 31188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_342
timestamp 1644511149
transform 1 0 32568 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_350
timestamp 1644511149
transform 1 0 33304 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_371
timestamp 1644511149
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1644511149
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_493
timestamp 1644511149
transform 1 0 46460 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1644511149
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_511
timestamp 1644511149
transform 1 0 48116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_515
timestamp 1644511149
transform 1 0 48484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_205
timestamp 1644511149
transform 1 0 19964 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_215
timestamp 1644511149
transform 1 0 20884 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_222
timestamp 1644511149
transform 1 0 21528 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_234
timestamp 1644511149
transform 1 0 22632 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_244
timestamp 1644511149
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1644511149
transform 1 0 26956 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_292
timestamp 1644511149
transform 1 0 27968 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_322
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_334
timestamp 1644511149
transform 1 0 31832 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_342
timestamp 1644511149
transform 1 0 32568 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_347
timestamp 1644511149
transform 1 0 33028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_368
timestamp 1644511149
transform 1 0 34960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_380
timestamp 1644511149
transform 1 0 36064 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_392
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_404
timestamp 1644511149
transform 1 0 38272 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1644511149
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_198
timestamp 1644511149
transform 1 0 19320 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_206
timestamp 1644511149
transform 1 0 20056 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1644511149
transform 1 0 22172 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_253
timestamp 1644511149
transform 1 0 24380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_263
timestamp 1644511149
transform 1 0 25300 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1644511149
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_286
timestamp 1644511149
transform 1 0 27416 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_294
timestamp 1644511149
transform 1 0 28152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1644511149
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_318
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1644511149
transform 1 0 31004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_344
timestamp 1644511149
transform 1 0 32752 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_352
timestamp 1644511149
transform 1 0 33488 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_370
timestamp 1644511149
transform 1 0 35144 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_377
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1644511149
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_173
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_186
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1644511149
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_208
timestamp 1644511149
transform 1 0 20240 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_218
timestamp 1644511149
transform 1 0 21160 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_230
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_243
timestamp 1644511149
transform 1 0 23460 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_247
timestamp 1644511149
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_313
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_323
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_327
timestamp 1644511149
transform 1 0 31188 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_348
timestamp 1644511149
transform 1 0 33120 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1644511149
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_374
timestamp 1644511149
transform 1 0 35512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_386
timestamp 1644511149
transform 1 0 36616 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_398
timestamp 1644511149
transform 1 0 37720 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_410
timestamp 1644511149
transform 1 0 38824 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_418
timestamp 1644511149
transform 1 0 39560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_186
timestamp 1644511149
transform 1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_197
timestamp 1644511149
transform 1 0 19228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_203
timestamp 1644511149
transform 1 0 19780 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_212
timestamp 1644511149
transform 1 0 20608 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_234
timestamp 1644511149
transform 1 0 22632 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_246
timestamp 1644511149
transform 1 0 23736 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_258
timestamp 1644511149
transform 1 0 24840 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_270
timestamp 1644511149
transform 1 0 25944 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1644511149
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_320
timestamp 1644511149
transform 1 0 30544 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_512
timestamp 1644511149
transform 1 0 48208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_207
timestamp 1644511149
transform 1 0 20148 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_214
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_238
timestamp 1644511149
transform 1 0 23000 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1644511149
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_259
timestamp 1644511149
transform 1 0 24932 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_267
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_275
timestamp 1644511149
transform 1 0 26404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_284
timestamp 1644511149
transform 1 0 27232 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_296
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_318
timestamp 1644511149
transform 1 0 30360 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1644511149
transform 1 0 31188 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_351
timestamp 1644511149
transform 1 0 33396 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1644511149
transform 1 0 33764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_200
timestamp 1644511149
transform 1 0 19504 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 1644511149
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1644511149
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_231
timestamp 1644511149
transform 1 0 22356 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_252
timestamp 1644511149
transform 1 0 24288 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_256
timestamp 1644511149
transform 1 0 24656 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_262
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_287
timestamp 1644511149
transform 1 0 27508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_299
timestamp 1644511149
transform 1 0 28612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_308
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1644511149
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_345
timestamp 1644511149
transform 1 0 32844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_357
timestamp 1644511149
transform 1 0 33948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_368
timestamp 1644511149
transform 1 0 34960 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_380
timestamp 1644511149
transform 1 0 36064 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_185
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_206
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1644511149
transform 1 0 21160 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_238
timestamp 1644511149
transform 1 0 23000 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_259
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_271
timestamp 1644511149
transform 1 0 26036 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1644511149
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_316
timestamp 1644511149
transform 1 0 30176 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_328
timestamp 1644511149
transform 1 0 31280 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_374
timestamp 1644511149
transform 1 0 35512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_386
timestamp 1644511149
transform 1 0 36616 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1644511149
transform 1 0 37720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_410
timestamp 1644511149
transform 1 0 38824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_418
timestamp 1644511149
transform 1 0 39560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_177
timestamp 1644511149
transform 1 0 17388 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_199
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_212
timestamp 1644511149
transform 1 0 20608 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_234
timestamp 1644511149
transform 1 0 22632 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_242
timestamp 1644511149
transform 1 0 23368 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_254
timestamp 1644511149
transform 1 0 24472 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_258
timestamp 1644511149
transform 1 0 24840 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_268
timestamp 1644511149
transform 1 0 25760 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_284
timestamp 1644511149
transform 1 0 27232 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_296
timestamp 1644511149
transform 1 0 28336 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_310
timestamp 1644511149
transform 1 0 29624 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_321
timestamp 1644511149
transform 1 0 30636 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_328
timestamp 1644511149
transform 1 0 31280 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_345
timestamp 1644511149
transform 1 0 32844 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_493
timestamp 1644511149
transform 1 0 46460 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_498
timestamp 1644511149
transform 1 0 46920 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_200
timestamp 1644511149
transform 1 0 19504 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_206
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_216
timestamp 1644511149
transform 1 0 20976 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_224
timestamp 1644511149
transform 1 0 21712 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_256
timestamp 1644511149
transform 1 0 24656 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_263
timestamp 1644511149
transform 1 0 25300 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_269
timestamp 1644511149
transform 1 0 25852 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_276
timestamp 1644511149
transform 1 0 26496 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_329
timestamp 1644511149
transform 1 0 31372 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_341
timestamp 1644511149
transform 1 0 32476 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_353
timestamp 1644511149
transform 1 0 33580 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_361
timestamp 1644511149
transform 1 0 34316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_511
timestamp 1644511149
transform 1 0 48116 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_515
timestamp 1644511149
transform 1 0 48484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_197
timestamp 1644511149
transform 1 0 19228 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_210
timestamp 1644511149
transform 1 0 20424 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_222
timestamp 1644511149
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_230
timestamp 1644511149
transform 1 0 22264 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_238
timestamp 1644511149
transform 1 0 23000 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_243
timestamp 1644511149
transform 1 0 23460 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_267
timestamp 1644511149
transform 1 0 25668 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_302
timestamp 1644511149
transform 1 0 28888 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_308
timestamp 1644511149
transform 1 0 29440 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_318
timestamp 1644511149
transform 1 0 30360 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_330
timestamp 1644511149
transform 1 0 31464 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_492
timestamp 1644511149
transform 1 0 46368 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_217
timestamp 1644511149
transform 1 0 21068 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_229
timestamp 1644511149
transform 1 0 22172 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_235
timestamp 1644511149
transform 1 0 22724 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_264
timestamp 1644511149
transform 1 0 25392 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_270
timestamp 1644511149
transform 1 0 25944 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_278
timestamp 1644511149
transform 1 0 26680 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_290
timestamp 1644511149
transform 1 0 27784 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1644511149
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_201
timestamp 1644511149
transform 1 0 19596 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_207
timestamp 1644511149
transform 1 0 20148 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_219
timestamp 1644511149
transform 1 0 21252 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_270
timestamp 1644511149
transform 1 0 25944 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1644511149
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_282
timestamp 1644511149
transform 1 0 27048 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_294
timestamp 1644511149
transform 1 0 28152 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1644511149
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_500
timestamp 1644511149
transform 1 0 47104 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1644511149
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_477
timestamp 1644511149
transform 1 0 44988 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_483
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_487
timestamp 1644511149
transform 1 0 45908 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_494
timestamp 1644511149
transform 1 0 46552 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1644511149
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_456
timestamp 1644511149
transform 1 0 43056 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_468
timestamp 1644511149
transform 1 0 44160 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_14
timestamp 1644511149
transform 1 0 2392 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_26
timestamp 1644511149
transform 1 0 3496 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_38
timestamp 1644511149
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1644511149
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_433
timestamp 1644511149
transform 1 0 40940 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_437
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_444
timestamp 1644511149
transform 1 0 41952 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_498
timestamp 1644511149
transform 1 0 46920 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_117
timestamp 1644511149
transform 1 0 11868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_188
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_200
timestamp 1644511149
transform 1 0 19504 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_212
timestamp 1644511149
transform 1 0 20608 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_338
timestamp 1644511149
transform 1 0 32200 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_350
timestamp 1644511149
transform 1 0 33304 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_354
timestamp 1644511149
transform 1 0 33672 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1644511149
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_368
timestamp 1644511149
transform 1 0 34960 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_380
timestamp 1644511149
transform 1 0 36064 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_392
timestamp 1644511149
transform 1 0 37168 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_400
timestamp 1644511149
transform 1 0 37904 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_461
timestamp 1644511149
transform 1 0 43516 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_465
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_32
timestamp 1644511149
transform 1 0 4048 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_44
timestamp 1644511149
transform 1 0 5152 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_218
timestamp 1644511149
transform 1 0 21160 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_383
timestamp 1644511149
transform 1 0 36340 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_63
timestamp 1644511149
transform 1 0 6900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1644511149
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_207
timestamp 1644511149
transform 1 0 20148 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_213
timestamp 1644511149
transform 1 0 20700 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_217
timestamp 1644511149
transform 1 0 21068 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1644511149
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_240
timestamp 1644511149
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1644511149
transform 1 0 24840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_317
timestamp 1644511149
transform 1 0 30268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_431
timestamp 1644511149
transform 1 0 40756 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_439
timestamp 1644511149
transform 1 0 41492 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_453
timestamp 1644511149
transform 1 0 42780 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_458
timestamp 1644511149
transform 1 0 43240 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0627_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0628_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0629_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0632_
timestamp 1644511149
transform 1 0 27232 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0633_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0634_
timestamp 1644511149
transform 1 0 26036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0635_
timestamp 1644511149
transform 1 0 25944 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0636_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0637_
timestamp 1644511149
transform 1 0 27140 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0639_
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0640_
timestamp 1644511149
transform 1 0 20240 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0641_
timestamp 1644511149
transform 1 0 20884 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0643_
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1644511149
transform 1 0 33488 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0647_
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0648_
timestamp 1644511149
transform 1 0 12696 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0650_
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0651_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0652_
timestamp 1644511149
transform 1 0 25300 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0653_
timestamp 1644511149
transform 1 0 16744 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0654_
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_2  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0656_
timestamp 1644511149
transform 1 0 16744 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1644511149
transform 1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0660_
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1644511149
transform 1 0 19872 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0666_
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0670_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1644511149
transform 1 0 14260 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0673_
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0675_
timestamp 1644511149
transform 1 0 12328 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0676_
timestamp 1644511149
transform 1 0 11960 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1644511149
transform 1 0 12420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0678_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0679_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0681_
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1644511149
transform 1 0 10580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0684_
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0686_
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 1644511149
transform 1 0 11316 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1644511149
transform 1 0 12972 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1644511149
transform 1 0 8648 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1644511149
transform 1 0 11500 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0699_
timestamp 1644511149
transform 1 0 9936 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0700_
timestamp 1644511149
transform 1 0 9292 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1644511149
transform 1 0 10212 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0703_
timestamp 1644511149
transform 1 0 19044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0705_
timestamp 1644511149
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0706_
timestamp 1644511149
transform 1 0 10028 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 13432 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0709_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0710_
timestamp 1644511149
transform 1 0 11684 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp 1644511149
transform 1 0 12972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1644511149
transform 1 0 11868 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 1644511149
transform 1 0 12328 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0715_
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0717_
timestamp 1644511149
transform 1 0 14628 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0719_
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0720_
timestamp 1644511149
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0721_
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0722_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0723_
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1644511149
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0727_
timestamp 1644511149
transform 1 0 15824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0729_
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1644511149
transform 1 0 19044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 1644511149
transform 1 0 21620 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0732_
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1644511149
transform 1 0 20884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0735_
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0736_
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0737_
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0738_
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1644511149
transform 1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0742_
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0743_
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0744_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0746_
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0747_
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0749_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0750_
timestamp 1644511149
transform 1 0 23552 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1644511149
transform 1 0 22908 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0752_
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0753_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0754_
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0755_
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0756_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1644511149
transform 1 0 26404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0758_
timestamp 1644511149
transform 1 0 24472 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0759_
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1644511149
transform 1 0 27048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0761_
timestamp 1644511149
transform 1 0 25392 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0763_
timestamp 1644511149
transform 1 0 28336 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_1  _0764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0768_
timestamp 1644511149
transform 1 0 25852 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0770_
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0771_
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0772_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0774_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0775_
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1644511149
transform 1 0 31648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0779_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0782_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0784_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0787_
timestamp 1644511149
transform 1 0 20148 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0789_
timestamp 1644511149
transform 1 0 20976 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0790_
timestamp 1644511149
transform 1 0 22632 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0791_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0792_
timestamp 1644511149
transform 1 0 21620 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0795_
timestamp 1644511149
transform 1 0 32292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0796_
timestamp 1644511149
transform 1 0 28796 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0797_
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0798_
timestamp 1644511149
transform 1 0 32200 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0799_
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0800_
timestamp 1644511149
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0801_
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0803_
timestamp 1644511149
transform 1 0 20056 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0804_
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _0805_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0806_
timestamp 1644511149
transform 1 0 28612 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0807_
timestamp 1644511149
transform 1 0 20424 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1644511149
transform 1 0 20516 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0811_
timestamp 1644511149
transform 1 0 27416 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1644511149
transform 1 0 19320 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0814_
timestamp 1644511149
transform 1 0 27140 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0815_
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1644511149
transform 1 0 21252 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0817_
timestamp 1644511149
transform 1 0 19320 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0818_
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0819_
timestamp 1644511149
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0820_
timestamp 1644511149
transform 1 0 28612 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0821_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0822_
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0823_
timestamp 1644511149
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1644511149
transform 1 0 20148 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1644511149
transform 1 0 18952 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0827_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1644511149
transform 1 0 19228 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1644511149
transform 1 0 19872 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0831_
timestamp 1644511149
transform 1 0 18216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0832_
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 1644511149
transform 1 0 18584 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0834_
timestamp 1644511149
transform 1 0 16652 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0835_
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0836_
timestamp 1644511149
transform 1 0 27324 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _0837_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0838_
timestamp 1644511149
transform 1 0 25944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0839_
timestamp 1644511149
transform 1 0 26036 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1644511149
transform 1 0 26220 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 1644511149
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0842_
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0843_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0844_
timestamp 1644511149
transform 1 0 26772 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0845_
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1644511149
transform 1 0 24932 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1644511149
transform 1 0 26864 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0852_
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0853_
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1644511149
transform 1 0 23460 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1644511149
transform 1 0 22356 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1644511149
transform 1 0 24472 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1644511149
transform 1 0 30728 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0861_
timestamp 1644511149
transform 1 0 28428 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0862_
timestamp 1644511149
transform 1 0 24656 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0865_
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0867_
timestamp 1644511149
transform 1 0 22724 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1644511149
transform 1 0 25484 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0869_
timestamp 1644511149
transform 1 0 24748 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0871_
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1644511149
transform 1 0 22632 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0873_
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0874_
timestamp 1644511149
transform 1 0 29072 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1644511149
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0876_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0877_
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0880_
timestamp 1644511149
transform 1 0 28980 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0881_
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _0882_
timestamp 1644511149
transform 1 0 27416 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0884_
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0885_
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0888_
timestamp 1644511149
transform 1 0 26404 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0890_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0891_
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0892_
timestamp 1644511149
transform 1 0 27048 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0893_
timestamp 1644511149
transform 1 0 22816 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0895_
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0896_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0897_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1644511149
transform 1 0 28888 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0899_
timestamp 1644511149
transform 1 0 28336 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0900_
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0901_
timestamp 1644511149
transform 1 0 28612 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0902_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0903_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0905_
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1644511149
transform 1 0 29348 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1644511149
transform 1 0 30544 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0908_
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0909_
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0910_
timestamp 1644511149
transform 1 0 30912 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0911_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0912_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0913_
timestamp 1644511149
transform 1 0 29808 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 1644511149
transform 1 0 29532 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0916_
timestamp 1644511149
transform 1 0 28612 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0918_
timestamp 1644511149
transform 1 0 29900 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1644511149
transform 1 0 34684 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0920_
timestamp 1644511149
transform 1 0 33488 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0921_
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0922_
timestamp 1644511149
transform 1 0 29992 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0923_
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 1644511149
transform 1 0 33120 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 1644511149
transform 1 0 32936 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1644511149
transform 1 0 35512 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 1644511149
transform 1 0 33396 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform 1 0 32752 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0933_
timestamp 1644511149
transform 1 0 34868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1644511149
transform 1 0 34500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0938_
timestamp 1644511149
transform 1 0 33856 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1644511149
transform 1 0 32660 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1644511149
transform 1 0 32660 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1644511149
transform 1 0 32568 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 1644511149
transform 1 0 33948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1644511149
transform 1 0 33212 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0945_
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0948_
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1644511149
transform 1 0 35144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0950_
timestamp 1644511149
transform 1 0 34776 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 33672 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 30912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 39836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 11960 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 31924 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0968_
timestamp 1644511149
transform 1 0 35236 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 35696 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 46276 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 25024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0981_
timestamp 1644511149
transform 1 0 18032 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0987_
timestamp 1644511149
transform 1 0 14904 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 12788 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 14076 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0993_
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 15364 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 41032 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43700 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 45632 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1012_
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1018_
timestamp 1644511149
transform 1 0 45356 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1020_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 45080 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 46092 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 46644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1024_
timestamp 1644511149
transform 1 0 45448 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 46644 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 43240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1030_
timestamp 1644511149
transform 1 0 44528 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 45264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 37076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1036_
timestamp 1644511149
transform 1 0 41400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1037_
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 8372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1043_
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1049_
timestamp 1644511149
transform 1 0 42320 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1644511149
transform 1 0 46644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 42780 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1055_
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1061_
timestamp 1644511149
transform 1 0 17296 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform 1 0 47288 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1644511149
transform 1 0 36156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1068_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1069_
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1071_
timestamp 1644511149
transform 1 0 32752 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33028 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46000 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1075_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1076_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1644511149
transform 1 0 45540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1078_
timestamp 1644511149
transform 1 0 45632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1080_
timestamp 1644511149
transform 1 0 46828 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _1081_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1083_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1084_
timestamp 1644511149
transform 1 0 39928 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1644511149
transform 1 0 40848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1087_
timestamp 1644511149
transform 1 0 40480 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1089_
timestamp 1644511149
transform 1 0 39928 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1092_
timestamp 1644511149
transform 1 0 43056 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 1644511149
transform 1 0 43240 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1094_
timestamp 1644511149
transform 1 0 43884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1096_
timestamp 1644511149
transform 1 0 42964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1097_
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1098_
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1099_
timestamp 1644511149
transform 1 0 28612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1100_
timestamp 1644511149
transform 1 0 28704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1101_
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1644511149
transform 1 0 46184 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1105_
timestamp 1644511149
transform 1 0 44436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1106_
timestamp 1644511149
transform 1 0 43608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1107_
timestamp 1644511149
transform 1 0 42688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1108_
timestamp 1644511149
transform 1 0 42780 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43148 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1644511149
transform 1 0 42504 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1644511149
transform 1 0 42136 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1113_
timestamp 1644511149
transform 1 0 43608 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1644511149
transform 1 0 43976 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1115_
timestamp 1644511149
transform 1 0 44068 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1116_
timestamp 1644511149
transform 1 0 45172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1118_
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1120_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1121_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp 1644511149
transform 1 0 29624 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1125_
timestamp 1644511149
transform 1 0 29716 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1644511149
transform 1 0 29716 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1127_
timestamp 1644511149
transform 1 0 30544 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1129_
timestamp 1644511149
transform 1 0 42964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1130_
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1131_
timestamp 1644511149
transform 1 0 39008 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1132_
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _1133_
timestamp 1644511149
transform 1 0 31096 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1134_
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1135_
timestamp 1644511149
transform 1 0 25668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1137_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1139_
timestamp 1644511149
transform 1 0 46092 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1140_
timestamp 1644511149
transform 1 0 46184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1141_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1142_
timestamp 1644511149
transform 1 0 36156 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1143_
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1144_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1145_
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1146_
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1147_
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1149_
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1644511149
transform 1 0 33856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1644511149
transform 1 0 32936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1153_
timestamp 1644511149
transform 1 0 31464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1644511149
transform 1 0 35696 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1644511149
transform 1 0 33488 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1644511149
transform 1 0 32476 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1644511149
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1644511149
transform 1 0 30728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1644511149
transform 1 0 31004 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1644511149
transform 1 0 31004 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1644511149
transform 1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1165_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1644511149
transform 1 0 23368 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1171_
timestamp 1644511149
transform 1 0 23000 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1644511149
transform 1 0 23552 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1644511149
transform 1 0 23184 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1644511149
transform 1 0 25024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1644511149
transform 1 0 21896 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1644511149
transform 1 0 22816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1644511149
transform 1 0 19872 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1644511149
transform 1 0 22080 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1183_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1644511149
transform 1 0 19504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1188_
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1189_
timestamp 1644511149
transform 1 0 29716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1190_
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1191_
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1192_
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1193_
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1195_
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1196_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1197_
timestamp 1644511149
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1198_
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1200_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1201_
timestamp 1644511149
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1202_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1644511149
transform 1 0 20056 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1204_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1205_
timestamp 1644511149
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1206_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1207_
timestamp 1644511149
transform 1 0 14720 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1208_
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1209_
timestamp 1644511149
transform 1 0 12696 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1644511149
transform 1 0 9200 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1212_
timestamp 1644511149
transform 1 0 8096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1213_
timestamp 1644511149
transform 1 0 8004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1214_
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1215_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1216_
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1218_
timestamp 1644511149
transform 1 0 10672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1219_
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1220_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1222_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1223_
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1644511149
transform 1 0 19320 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1644511149
transform 1 0 32476 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1644511149
transform 1 0 32384 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1644511149
transform 1 0 33488 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 1644511149
transform 1 0 33396 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1644511149
transform 1 0 32384 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1232_
timestamp 1644511149
transform 1 0 31280 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1233_
timestamp 1644511149
transform 1 0 31004 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1235_
timestamp 1644511149
transform 1 0 29808 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1644511149
transform 1 0 30084 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1644511149
transform 1 0 28520 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 1644511149
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1644511149
transform 1 0 21988 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1644511149
transform 1 0 22540 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1644511149
transform 1 0 25116 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1247_
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1248_
timestamp 1644511149
transform 1 0 23828 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1249_
timestamp 1644511149
transform 1 0 24104 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 1644511149
transform 1 0 17480 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 1644511149
transform 1 0 17572 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1252_
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1644511149
transform 1 0 21160 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 1644511149
transform 1 0 17848 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1257_
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1258_
timestamp 1644511149
transform 1 0 30360 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1259_
timestamp 1644511149
transform 1 0 29716 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1260_
timestamp 1644511149
transform 1 0 26220 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1261_
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1644511149
transform 1 0 25392 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1263_
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 1644511149
transform 1 0 24104 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1267_
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1269_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1270_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1271_
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 1644511149
transform 1 0 14996 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1274_
timestamp 1644511149
transform 1 0 15088 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1275_
timestamp 1644511149
transform 1 0 12144 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1276_
timestamp 1644511149
transform 1 0 11684 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1277_
timestamp 1644511149
transform 1 0 9384 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1278_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1279_
timestamp 1644511149
transform 1 0 7912 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1280_
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 1644511149
transform 1 0 9016 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1282_
timestamp 1644511149
transform 1 0 9844 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1283_
timestamp 1644511149
transform 1 0 11592 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1284_
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1644511149
transform 1 0 14260 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1286_
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1290_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1291__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1292__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1293__83
timestamp 1644511149
transform 1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1294__84
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1295__85
timestamp 1644511149
transform 1 0 47472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1296__86
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1297__87
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1298__88
timestamp 1644511149
transform 1 0 24564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1299__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1300__90
timestamp 1644511149
transform 1 0 25208 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1301__91
timestamp 1644511149
transform 1 0 47932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1302__92
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1303__93
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1304__94
timestamp 1644511149
transform 1 0 33396 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1305__95
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1306__96
timestamp 1644511149
transform 1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1307__97
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1308__98
timestamp 1644511149
transform 1 0 43608 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1309__99
timestamp 1644511149
transform 1 0 41492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1310__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1311__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1312__102
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1313__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1314__104
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1315__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1316__106
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1317__107
timestamp 1644511149
transform 1 0 46828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1318__108
timestamp 1644511149
transform 1 0 45908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1319__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1320__110
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1321__111
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1322__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1323__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1324__114
timestamp 1644511149
transform 1 0 43424 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1325__115
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1326__116
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1327__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1328__118
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1329__119
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1330__120
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1331__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1332__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1333__123
timestamp 1644511149
transform 1 0 45632 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1334__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1335__125
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1336__126
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1337__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1338__128
timestamp 1644511149
transform 1 0 47472 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1339__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1340__130
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1341__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1342__132
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1343__133
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1344__134
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1345__135
timestamp 1644511149
transform 1 0 44712 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 30544 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 33580 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 45080 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 33672 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 46184 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 32936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 34408 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1378_
timestamp 1644511149
transform 1 0 35696 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1379_
timestamp 1644511149
transform 1 0 35052 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1380_
timestamp 1644511149
transform 1 0 26680 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1381_
timestamp 1644511149
transform 1 0 20608 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1382_
timestamp 1644511149
transform 1 0 26496 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1383_
timestamp 1644511149
transform 1 0 29716 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1384_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1385_
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1386_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1387_
timestamp 1644511149
transform 1 0 22724 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1388_
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1389_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1390_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1391_
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1392_
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1393_
timestamp 1644511149
transform 1 0 14812 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1394_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1395_
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1396_
timestamp 1644511149
transform 1 0 9568 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1397_
timestamp 1644511149
transform 1 0 11684 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1398_
timestamp 1644511149
transform 1 0 9016 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1399_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1400_
timestamp 1644511149
transform 1 0 14260 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1401_
timestamp 1644511149
transform 1 0 9292 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1402_
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1403_
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1404_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1405_
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1406_
timestamp 1644511149
transform 1 0 15732 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1407_
timestamp 1644511149
transform 1 0 20148 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1408_
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1409_
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1410_
timestamp 1644511149
transform 1 0 9292 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1411_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1412_
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1413_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1414_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1415_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1416_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1417_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1418_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1419_
timestamp 1644511149
transform 1 0 41216 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1420_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1421_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1422_
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1423_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1424_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1425_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1426_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1427_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1428_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1429_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1430_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1431_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1432_
timestamp 1644511149
transform 1 0 19228 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1433_
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1434_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1435_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1436_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1437_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1438_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1439_
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1440_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1441_
timestamp 1644511149
transform 1 0 44988 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26128 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 28980 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 29900 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 47288 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 47932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 46184 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 46736 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1644511149
transform 1 0 47840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 42872 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1644511149
transform 1 0 46184 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1644511149
transform 1 0 43608 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1644511149
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 43884 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 43976 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 39376 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 40020 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 40848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 41492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 40204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 19872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2024 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 46828 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 34592 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29900 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35052 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46644 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 42596 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 37536 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 32292 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 45724 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 40020 0 -1 23936
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
