magic
tech sky130A
magscale 1 2
timestamp 1654172904
<< viali >>
rect 19441 47141 19475 47175
rect 29929 47141 29963 47175
rect 47961 47141 47995 47175
rect 14105 47073 14139 47107
rect 16957 47073 16991 47107
rect 30757 47073 30791 47107
rect 43177 47073 43211 47107
rect 47041 47073 47075 47107
rect 2145 47005 2179 47039
rect 2973 47005 3007 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6837 47005 6871 47039
rect 7757 47005 7791 47039
rect 9413 47005 9447 47039
rect 11621 47005 11655 47039
rect 12357 47005 12391 47039
rect 13093 47005 13127 47039
rect 14381 47005 14415 47039
rect 16681 47005 16715 47039
rect 19257 47005 19291 47039
rect 20269 47005 20303 47039
rect 20913 47005 20947 47039
rect 22017 47005 22051 47039
rect 24777 47005 24811 47039
rect 25513 47005 25547 47039
rect 28641 47005 28675 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38393 47005 38427 47039
rect 41889 47005 41923 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 2513 46937 2547 46971
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 7941 46937 7975 46971
rect 9597 46937 9631 46971
rect 11805 46937 11839 46971
rect 12541 46937 12575 46971
rect 13461 46937 13495 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 3157 46869 3191 46903
rect 6929 46869 6963 46903
rect 21833 46869 21867 46903
rect 28457 46869 28491 46903
rect 1869 46597 1903 46631
rect 28457 46597 28491 46631
rect 30113 46597 30147 46631
rect 19441 46529 19475 46563
rect 24593 46529 24627 46563
rect 28273 46529 28307 46563
rect 38117 46529 38151 46563
rect 41705 46529 41739 46563
rect 42441 46529 42475 46563
rect 47869 46529 47903 46563
rect 3433 46461 3467 46495
rect 3617 46461 3651 46495
rect 4169 46461 4203 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 11989 46461 12023 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19625 46461 19659 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41797 46461 41831 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 2145 46325 2179 46359
rect 2881 46325 2915 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 3893 46121 3927 46155
rect 4629 46121 4663 46155
rect 11253 46121 11287 46155
rect 14289 46121 14323 46155
rect 20177 46121 20211 46155
rect 24685 46121 24719 46155
rect 38301 46121 38335 46155
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41337 45985 41371 46019
rect 41981 45985 42015 46019
rect 47041 45985 47075 46019
rect 2881 45917 2915 45951
rect 3801 45917 3835 45951
rect 11161 45917 11195 45951
rect 20085 45917 20119 45951
rect 24593 45917 24627 45951
rect 38209 45917 38243 45951
rect 43913 45917 43947 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 20913 45849 20947 45883
rect 25421 45849 25455 45883
rect 41521 45849 41555 45883
rect 46489 45849 46523 45883
rect 2973 45781 3007 45815
rect 44097 45781 44131 45815
rect 45753 45781 45787 45815
rect 13829 45577 13863 45611
rect 20913 45577 20947 45611
rect 25421 45577 25455 45611
rect 32229 45577 32263 45611
rect 41521 45577 41555 45611
rect 2237 45509 2271 45543
rect 42901 45509 42935 45543
rect 43913 45509 43947 45543
rect 46949 45509 46983 45543
rect 47961 45509 47995 45543
rect 13737 45441 13771 45475
rect 20821 45441 20855 45475
rect 25329 45441 25363 45475
rect 32137 45441 32171 45475
rect 41429 45441 41463 45475
rect 42809 45441 42843 45475
rect 46857 45441 46891 45475
rect 2053 45373 2087 45407
rect 3065 45373 3099 45407
rect 44557 45373 44591 45407
rect 44741 45373 44775 45407
rect 45661 45373 45695 45407
rect 44005 45237 44039 45271
rect 48053 45237 48087 45271
rect 42901 45033 42935 45067
rect 44465 45033 44499 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 46949 44489 46983 44523
rect 45109 44353 45143 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 47685 44149 47719 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1869 43265 1903 43299
rect 25881 43265 25915 43299
rect 47041 43265 47075 43299
rect 47777 43265 47811 43299
rect 1961 43061 1995 43095
rect 25973 43061 26007 43095
rect 25973 42721 26007 42755
rect 27629 42721 27663 42755
rect 25789 42653 25823 42687
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 25237 42313 25271 42347
rect 47685 42313 47719 42347
rect 25145 42177 25179 42211
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 2237 41225 2271 41259
rect 46857 41225 46891 41259
rect 2145 41089 2179 41123
rect 46765 41089 46799 41123
rect 47961 41089 47995 41123
rect 48145 40953 48179 40987
rect 47685 40681 47719 40715
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 47777 39797 47811 39831
rect 46305 39457 46339 39491
rect 48145 39457 48179 39491
rect 46489 39321 46523 39355
rect 46949 39049 46983 39083
rect 46857 38913 46891 38947
rect 47777 38913 47811 38947
rect 47869 38709 47903 38743
rect 46305 38301 46339 38335
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 47685 37961 47719 37995
rect 19625 37825 19659 37859
rect 47593 37825 47627 37859
rect 24409 37757 24443 37791
rect 24685 37757 24719 37791
rect 19441 37621 19475 37655
rect 26157 37621 26191 37655
rect 25053 37417 25087 37451
rect 47685 37417 47719 37451
rect 19533 37281 19567 37315
rect 26341 37281 26375 37315
rect 27261 37281 27295 37315
rect 19257 37213 19291 37247
rect 22753 37213 22787 37247
rect 23581 37213 23615 37247
rect 25237 37213 25271 37247
rect 26985 37213 27019 37247
rect 21005 37077 21039 37111
rect 22937 37077 22971 37111
rect 23673 37077 23707 37111
rect 26617 37077 26651 37111
rect 27077 37077 27111 37111
rect 19441 36873 19475 36907
rect 20361 36873 20395 36907
rect 21189 36873 21223 36907
rect 20269 36805 20303 36839
rect 19073 36737 19107 36771
rect 21097 36737 21131 36771
rect 25329 36737 25363 36771
rect 19165 36669 19199 36703
rect 20545 36669 20579 36703
rect 22661 36669 22695 36703
rect 22937 36669 22971 36703
rect 25421 36669 25455 36703
rect 25697 36669 25731 36703
rect 19901 36533 19935 36567
rect 24409 36533 24443 36567
rect 19717 36329 19751 36363
rect 22753 36329 22787 36363
rect 24501 36329 24535 36363
rect 23121 36261 23155 36295
rect 2789 36193 2823 36227
rect 20177 36193 20211 36227
rect 20361 36193 20395 36227
rect 1409 36125 1443 36159
rect 20085 36125 20119 36159
rect 22937 36125 22971 36159
rect 23213 36125 23247 36159
rect 24409 36125 24443 36159
rect 1593 36057 1627 36091
rect 2053 35649 2087 35683
rect 22477 35649 22511 35683
rect 23765 35649 23799 35683
rect 27169 35649 27203 35683
rect 28273 35581 28307 35615
rect 28549 35581 28583 35615
rect 23949 35513 23983 35547
rect 22569 35445 22603 35479
rect 27261 35445 27295 35479
rect 30021 35445 30055 35479
rect 2237 35241 2271 35275
rect 19717 35241 19751 35275
rect 24961 35241 24995 35275
rect 29653 35241 29687 35275
rect 18705 35173 18739 35207
rect 16957 35105 16991 35139
rect 19625 35105 19659 35139
rect 21557 35105 21591 35139
rect 25145 35105 25179 35139
rect 26157 35105 26191 35139
rect 26433 35105 26467 35139
rect 1593 35037 1627 35071
rect 2145 35037 2179 35071
rect 14749 35037 14783 35071
rect 19533 35037 19567 35071
rect 20913 35037 20947 35071
rect 25237 35037 25271 35071
rect 29561 35037 29595 35071
rect 31125 35037 31159 35071
rect 47317 35037 47351 35071
rect 47593 35037 47627 35071
rect 15025 34969 15059 35003
rect 17233 34969 17267 35003
rect 21833 34969 21867 35003
rect 24961 34969 24995 35003
rect 1409 34901 1443 34935
rect 16497 34901 16531 34935
rect 19901 34901 19935 34935
rect 21005 34901 21039 34935
rect 23305 34901 23339 34935
rect 25421 34901 25455 34935
rect 27905 34901 27939 34935
rect 31217 34901 31251 34935
rect 17141 34697 17175 34731
rect 18521 34697 18555 34731
rect 22569 34697 22603 34731
rect 29009 34697 29043 34731
rect 27077 34629 27111 34663
rect 15853 34561 15887 34595
rect 17049 34561 17083 34595
rect 17785 34561 17819 34595
rect 17969 34561 18003 34595
rect 18337 34561 18371 34595
rect 18981 34561 19015 34595
rect 19165 34561 19199 34595
rect 19533 34561 19567 34595
rect 19717 34561 19751 34595
rect 20361 34561 20395 34595
rect 20545 34561 20579 34595
rect 20637 34561 20671 34595
rect 21833 34561 21867 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 22385 34561 22419 34595
rect 24225 34561 24259 34595
rect 26985 34561 27019 34595
rect 28273 34561 28307 34595
rect 28457 34561 28491 34595
rect 28641 34561 28675 34595
rect 28825 34561 28859 34595
rect 29837 34561 29871 34595
rect 48145 34561 48179 34595
rect 18061 34493 18095 34527
rect 18153 34493 18187 34527
rect 19257 34493 19291 34527
rect 19349 34493 19383 34527
rect 22109 34493 22143 34527
rect 24501 34493 24535 34527
rect 28549 34493 28583 34527
rect 30113 34493 30147 34527
rect 25973 34425 26007 34459
rect 16037 34357 16071 34391
rect 20177 34357 20211 34391
rect 31585 34357 31619 34391
rect 47961 34357 47995 34391
rect 16405 34153 16439 34187
rect 25237 34153 25271 34187
rect 28733 34153 28767 34187
rect 29009 34153 29043 34187
rect 30297 34153 30331 34187
rect 31125 34153 31159 34187
rect 27813 34085 27847 34119
rect 20177 34017 20211 34051
rect 24961 34017 24995 34051
rect 28733 34017 28767 34051
rect 29831 34017 29865 34051
rect 31217 34017 31251 34051
rect 46305 34017 46339 34051
rect 16313 33949 16347 33983
rect 25053 33949 25087 33983
rect 25697 33949 25731 33983
rect 27629 33949 27663 33983
rect 28457 33949 28491 33983
rect 29561 33927 29595 33961
rect 29745 33947 29779 33981
rect 29929 33949 29963 33983
rect 30113 33949 30147 33983
rect 30941 33949 30975 33983
rect 31769 33949 31803 33983
rect 20453 33881 20487 33915
rect 25881 33881 25915 33915
rect 30757 33881 30791 33915
rect 46489 33881 46523 33915
rect 48145 33881 48179 33915
rect 21925 33813 21959 33847
rect 24593 33813 24627 33847
rect 26065 33813 26099 33847
rect 30665 33813 30699 33847
rect 31861 33813 31895 33847
rect 18061 33609 18095 33643
rect 19533 33609 19567 33643
rect 20545 33609 20579 33643
rect 22385 33609 22419 33643
rect 23765 33609 23799 33643
rect 23949 33609 23983 33643
rect 27261 33609 27295 33643
rect 28733 33609 28767 33643
rect 24869 33541 24903 33575
rect 17693 33473 17727 33507
rect 18981 33473 19015 33507
rect 20177 33473 20211 33507
rect 20361 33473 20395 33507
rect 21833 33473 21867 33507
rect 22201 33473 22235 33507
rect 23029 33473 23063 33507
rect 23890 33473 23924 33507
rect 25145 33473 25179 33507
rect 25789 33473 25823 33507
rect 25973 33473 26007 33507
rect 26985 33473 27019 33507
rect 27905 33473 27939 33507
rect 28089 33473 28123 33507
rect 28917 33473 28951 33507
rect 29009 33473 29043 33507
rect 29193 33473 29227 33507
rect 29285 33473 29319 33507
rect 29745 33473 29779 33507
rect 30021 33473 30055 33507
rect 30665 33473 30699 33507
rect 30849 33473 30883 33507
rect 47869 33473 47903 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 17785 33405 17819 33439
rect 19257 33405 19291 33439
rect 23305 33405 23339 33439
rect 24409 33405 24443 33439
rect 24961 33405 24995 33439
rect 27261 33405 27295 33439
rect 27997 33405 28031 33439
rect 29929 33405 29963 33439
rect 22845 33337 22879 33371
rect 24317 33337 24351 33371
rect 25329 33337 25363 33371
rect 27077 33337 27111 33371
rect 30205 33337 30239 33371
rect 31033 33337 31067 33371
rect 17693 33269 17727 33303
rect 19349 33269 19383 33303
rect 22201 33269 22235 33303
rect 23213 33269 23247 33303
rect 25145 33269 25179 33303
rect 25789 33269 25823 33303
rect 30021 33269 30055 33303
rect 30849 33269 30883 33303
rect 48053 33269 48087 33303
rect 17417 33065 17451 33099
rect 21649 33065 21683 33099
rect 23397 33065 23431 33099
rect 24409 33065 24443 33099
rect 24869 33065 24903 33099
rect 25973 33065 26007 33099
rect 17785 32997 17819 33031
rect 20637 32997 20671 33031
rect 29009 32997 29043 33031
rect 1409 32929 1443 32963
rect 19533 32929 19567 32963
rect 23213 32929 23247 32963
rect 24777 32929 24811 32963
rect 25605 32929 25639 32963
rect 30389 32929 30423 32963
rect 30665 32929 30699 32963
rect 16681 32861 16715 32895
rect 16957 32861 16991 32895
rect 17601 32861 17635 32895
rect 17877 32861 17911 32895
rect 18337 32861 18371 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 20637 32861 20671 32895
rect 20913 32861 20947 32895
rect 22201 32861 22235 32895
rect 22385 32861 22419 32895
rect 23121 32861 23155 32895
rect 23397 32861 23431 32895
rect 24685 32861 24719 32895
rect 24961 32861 24995 32895
rect 25145 32861 25179 32895
rect 25789 32861 25823 32895
rect 26065 32861 26099 32895
rect 26525 32861 26559 32895
rect 26709 32861 26743 32895
rect 28641 32861 28675 32895
rect 28825 32861 28859 32895
rect 30297 32861 30331 32895
rect 31217 32861 31251 32895
rect 46305 32861 46339 32895
rect 1593 32793 1627 32827
rect 3249 32793 3283 32827
rect 16865 32793 16899 32827
rect 20821 32793 20855 32827
rect 21557 32793 21591 32827
rect 27997 32793 28031 32827
rect 28181 32793 28215 32827
rect 31493 32793 31527 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 16497 32725 16531 32759
rect 18705 32725 18739 32759
rect 22293 32725 22327 32759
rect 23581 32725 23615 32759
rect 26617 32725 26651 32759
rect 32965 32725 32999 32759
rect 17233 32521 17267 32555
rect 19257 32521 19291 32555
rect 25237 32521 25271 32555
rect 27629 32521 27663 32555
rect 31585 32521 31619 32555
rect 47685 32521 47719 32555
rect 2053 32453 2087 32487
rect 16037 32453 16071 32487
rect 16865 32453 16899 32487
rect 16957 32453 16991 32487
rect 25078 32453 25112 32487
rect 27261 32453 27295 32487
rect 15301 32385 15335 32419
rect 15945 32385 15979 32419
rect 16129 32385 16163 32419
rect 16681 32385 16715 32419
rect 17049 32385 17083 32419
rect 17785 32385 17819 32419
rect 18061 32385 18095 32419
rect 18245 32385 18279 32419
rect 18889 32385 18923 32419
rect 19073 32385 19107 32419
rect 20177 32385 20211 32419
rect 24317 32385 24351 32419
rect 24961 32385 24995 32419
rect 25789 32385 25823 32419
rect 26985 32385 27019 32419
rect 27078 32385 27112 32419
rect 27353 32385 27387 32419
rect 27491 32385 27525 32419
rect 28641 32385 28675 32419
rect 28825 32385 28859 32419
rect 30941 32385 30975 32419
rect 31034 32385 31068 32419
rect 31217 32385 31251 32419
rect 31309 32385 31343 32419
rect 31447 32385 31481 32419
rect 47041 32385 47075 32419
rect 47593 32385 47627 32419
rect 1869 32317 1903 32351
rect 3249 32317 3283 32351
rect 20453 32317 20487 32351
rect 24593 32317 24627 32351
rect 24869 32317 24903 32351
rect 26249 32317 26283 32351
rect 15393 32181 15427 32215
rect 18245 32181 18279 32215
rect 18429 32181 18463 32215
rect 25881 32181 25915 32215
rect 28733 32181 28767 32215
rect 1409 31977 1443 32011
rect 17233 31977 17267 32011
rect 18429 31977 18463 32011
rect 18521 31977 18555 32011
rect 19533 31977 19567 32011
rect 21281 31977 21315 32011
rect 28641 31977 28675 32011
rect 30849 31977 30883 32011
rect 16681 31909 16715 31943
rect 17969 31909 18003 31943
rect 22017 31909 22051 31943
rect 14933 31841 14967 31875
rect 15209 31841 15243 31875
rect 18337 31841 18371 31875
rect 19349 31841 19383 31875
rect 23397 31841 23431 31875
rect 47317 31841 47351 31875
rect 47593 31841 47627 31875
rect 1593 31773 1627 31807
rect 2329 31773 2363 31807
rect 2789 31773 2823 31807
rect 17233 31773 17267 31807
rect 17417 31773 17451 31807
rect 18245 31773 18279 31807
rect 18705 31773 18739 31807
rect 19257 31773 19291 31807
rect 19533 31773 19567 31807
rect 20637 31773 20671 31807
rect 20785 31773 20819 31807
rect 21102 31773 21136 31807
rect 21833 31773 21867 31807
rect 23213 31773 23247 31807
rect 24869 31773 24903 31807
rect 25237 31773 25271 31807
rect 27169 31773 27203 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 30849 31773 30883 31807
rect 31033 31773 31067 31807
rect 20913 31705 20947 31739
rect 21005 31705 21039 31739
rect 27905 31705 27939 31739
rect 28089 31705 28123 31739
rect 2881 31637 2915 31671
rect 19717 31637 19751 31671
rect 27261 31637 27295 31671
rect 17877 31433 17911 31467
rect 22293 31433 22327 31467
rect 2237 31365 2271 31399
rect 22201 31365 22235 31399
rect 2053 31297 2087 31331
rect 18061 31297 18095 31331
rect 18245 31297 18279 31331
rect 18337 31297 18371 31331
rect 20361 31297 20395 31331
rect 20545 31297 20579 31331
rect 20637 31297 20671 31331
rect 20729 31297 20763 31331
rect 22845 31297 22879 31331
rect 23029 31297 23063 31331
rect 23213 31297 23247 31331
rect 23949 31297 23983 31331
rect 25145 31297 25179 31331
rect 26249 31297 26283 31331
rect 26433 31297 26467 31331
rect 27537 31297 27571 31331
rect 30849 31297 30883 31331
rect 31033 31297 31067 31331
rect 31125 31297 31159 31331
rect 2789 31229 2823 31263
rect 23673 31229 23707 31263
rect 27813 31229 27847 31263
rect 20913 31093 20947 31127
rect 25237 31093 25271 31127
rect 26249 31093 26283 31127
rect 29285 31093 29319 31127
rect 30665 31093 30699 31127
rect 19625 30889 19659 30923
rect 23581 30889 23615 30923
rect 23765 30889 23799 30923
rect 26065 30889 26099 30923
rect 27537 30889 27571 30923
rect 29009 30889 29043 30923
rect 30573 30889 30607 30923
rect 21189 30753 21223 30787
rect 31033 30753 31067 30787
rect 31309 30753 31343 30787
rect 16129 30685 16163 30719
rect 17601 30685 17635 30719
rect 17693 30685 17727 30719
rect 18061 30685 18095 30719
rect 19257 30685 19291 30719
rect 21097 30685 21131 30719
rect 22661 30685 22695 30719
rect 27169 30685 27203 30719
rect 27353 30685 27387 30719
rect 28365 30685 28399 30719
rect 28513 30685 28547 30719
rect 28830 30685 28864 30719
rect 30021 30685 30055 30719
rect 30389 30685 30423 30719
rect 17785 30617 17819 30651
rect 17923 30617 17957 30651
rect 19441 30617 19475 30651
rect 23397 30617 23431 30651
rect 23581 30617 23615 30651
rect 24777 30617 24811 30651
rect 28641 30617 28675 30651
rect 28733 30617 28767 30651
rect 30205 30617 30239 30651
rect 30297 30617 30331 30651
rect 16221 30549 16255 30583
rect 17417 30549 17451 30583
rect 21465 30549 21499 30583
rect 22845 30549 22879 30583
rect 32781 30549 32815 30583
rect 17417 30345 17451 30379
rect 28549 30345 28583 30379
rect 31033 30345 31067 30379
rect 20085 30277 20119 30311
rect 23121 30277 23155 30311
rect 23581 30277 23615 30311
rect 29377 30277 29411 30311
rect 32321 30277 32355 30311
rect 15945 30209 15979 30243
rect 16957 30209 16991 30243
rect 18153 30209 18187 30243
rect 18245 30209 18279 30243
rect 18337 30209 18371 30243
rect 18521 30209 18555 30243
rect 18981 30209 19015 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 21189 30209 21223 30243
rect 23305 30209 23339 30243
rect 23489 30209 23523 30243
rect 24041 30209 24075 30243
rect 24409 30209 24443 30243
rect 24685 30209 24719 30243
rect 25605 30209 25639 30243
rect 25789 30209 25823 30243
rect 25881 30209 25915 30243
rect 27353 30209 27387 30243
rect 27905 30209 27939 30243
rect 28365 30209 28399 30243
rect 29561 30209 29595 30243
rect 29745 30209 29779 30243
rect 30665 30209 30699 30243
rect 32229 30209 32263 30243
rect 24501 30141 24535 30175
rect 25697 30141 25731 30175
rect 28181 30141 28215 30175
rect 30757 30141 30791 30175
rect 17325 30073 17359 30107
rect 27537 30073 27571 30107
rect 29101 30073 29135 30107
rect 16037 30005 16071 30039
rect 17877 30005 17911 30039
rect 19165 30005 19199 30039
rect 20177 30005 20211 30039
rect 20729 30005 20763 30039
rect 25421 30005 25455 30039
rect 16773 29801 16807 29835
rect 21649 29801 21683 29835
rect 25586 29801 25620 29835
rect 28365 29801 28399 29835
rect 32229 29801 32263 29835
rect 23489 29733 23523 29767
rect 24409 29733 24443 29767
rect 27813 29733 27847 29767
rect 15025 29665 15059 29699
rect 17693 29665 17727 29699
rect 17785 29665 17819 29699
rect 22753 29665 22787 29699
rect 25329 29665 25363 29699
rect 31493 29665 31527 29699
rect 47593 29665 47627 29699
rect 19441 29597 19475 29631
rect 19717 29597 19751 29631
rect 21281 29597 21315 29631
rect 21649 29597 21683 29631
rect 22293 29597 22327 29631
rect 22477 29597 22511 29631
rect 22661 29597 22695 29631
rect 23305 29597 23339 29631
rect 24685 29597 24719 29631
rect 28273 29597 28307 29631
rect 29561 29597 29595 29631
rect 30297 29597 30331 29631
rect 31309 29597 31343 29631
rect 31585 29597 31619 29631
rect 32137 29597 32171 29631
rect 47317 29597 47351 29631
rect 15301 29529 15335 29563
rect 19625 29529 19659 29563
rect 24409 29529 24443 29563
rect 27629 29529 27663 29563
rect 30481 29529 30515 29563
rect 17233 29461 17267 29495
rect 17601 29461 17635 29495
rect 19257 29461 19291 29495
rect 21833 29461 21867 29495
rect 24593 29461 24627 29495
rect 27077 29461 27111 29495
rect 29745 29461 29779 29495
rect 30665 29461 30699 29495
rect 31125 29461 31159 29495
rect 20545 29257 20579 29291
rect 23397 29257 23431 29291
rect 27169 29257 27203 29291
rect 31493 29257 31527 29291
rect 34345 29257 34379 29291
rect 27077 29189 27111 29223
rect 29837 29189 29871 29223
rect 15945 29121 15979 29155
rect 18797 29121 18831 29155
rect 21833 29121 21867 29155
rect 22005 29119 22039 29153
rect 22385 29121 22419 29155
rect 23029 29121 23063 29155
rect 23213 29121 23247 29155
rect 24685 29121 24719 29155
rect 28089 29121 28123 29155
rect 30941 29121 30975 29155
rect 31217 29121 31251 29155
rect 19073 29053 19107 29087
rect 22109 29053 22143 29087
rect 22201 29053 22235 29087
rect 32597 29053 32631 29087
rect 32873 29053 32907 29087
rect 15761 28985 15795 29019
rect 22569 28985 22603 29019
rect 24869 28985 24903 29019
rect 28273 28985 28307 29019
rect 29929 28917 29963 28951
rect 31309 28917 31343 28951
rect 15564 28713 15598 28747
rect 27077 28713 27111 28747
rect 30665 28713 30699 28747
rect 31125 28713 31159 28747
rect 32781 28713 32815 28747
rect 33425 28713 33459 28747
rect 17049 28645 17083 28679
rect 15301 28577 15335 28611
rect 20085 28577 20119 28611
rect 21557 28577 21591 28611
rect 30849 28577 30883 28611
rect 32321 28577 32355 28611
rect 32413 28577 32447 28611
rect 19809 28509 19843 28543
rect 22201 28509 22235 28543
rect 23581 28509 23615 28543
rect 23765 28509 23799 28543
rect 24777 28509 24811 28543
rect 24961 28509 24995 28543
rect 25145 28509 25179 28543
rect 25973 28509 26007 28543
rect 26985 28509 27019 28543
rect 27813 28509 27847 28543
rect 28549 28509 28583 28543
rect 29653 28509 29687 28543
rect 29745 28509 29779 28543
rect 30941 28509 30975 28543
rect 32045 28509 32079 28543
rect 32229 28509 32263 28543
rect 32597 28509 32631 28543
rect 33333 28509 33367 28543
rect 22017 28441 22051 28475
rect 25053 28441 25087 28475
rect 25789 28441 25823 28475
rect 30665 28441 30699 28475
rect 22385 28373 22419 28407
rect 23765 28373 23799 28407
rect 25329 28373 25363 28407
rect 26157 28373 26191 28407
rect 27905 28373 27939 28407
rect 28733 28373 28767 28407
rect 29929 28373 29963 28407
rect 19993 28169 20027 28203
rect 20821 28169 20855 28203
rect 24501 28169 24535 28203
rect 24961 28169 24995 28203
rect 28641 28169 28675 28203
rect 29653 28169 29687 28203
rect 13737 28101 13771 28135
rect 22293 28101 22327 28135
rect 22385 28101 22419 28135
rect 23121 28101 23155 28135
rect 24041 28101 24075 28135
rect 36461 28101 36495 28135
rect 37473 28101 37507 28135
rect 8401 28033 8435 28067
rect 13553 28033 13587 28067
rect 13829 28033 13863 28067
rect 14289 28033 14323 28067
rect 15025 28033 15059 28067
rect 15209 28033 15243 28067
rect 19901 28033 19935 28067
rect 20729 28033 20763 28067
rect 22201 28033 22235 28067
rect 22569 28033 22603 28067
rect 22661 28033 22695 28067
rect 23397 28033 23431 28067
rect 24317 28033 24351 28067
rect 25237 28033 25271 28067
rect 25421 28033 25455 28067
rect 25697 28033 25731 28067
rect 26341 28033 26375 28067
rect 28582 28033 28616 28067
rect 29101 28033 29135 28067
rect 29561 28033 29595 28067
rect 30389 28033 30423 28067
rect 30481 28033 30515 28067
rect 30665 28033 30699 28067
rect 30767 28055 30801 28089
rect 31217 28033 31251 28067
rect 31401 28033 31435 28067
rect 32781 28033 32815 28067
rect 36369 28033 36403 28067
rect 8585 27965 8619 27999
rect 8861 27965 8895 27999
rect 23213 27965 23247 27999
rect 24225 27965 24259 27999
rect 29009 27965 29043 27999
rect 37289 27965 37323 27999
rect 39129 27965 39163 27999
rect 13553 27897 13587 27931
rect 14473 27897 14507 27931
rect 23581 27897 23615 27931
rect 15025 27829 15059 27863
rect 22017 27829 22051 27863
rect 23121 27829 23155 27863
rect 24317 27829 24351 27863
rect 25329 27829 25363 27863
rect 25513 27829 25547 27863
rect 26157 27829 26191 27863
rect 28457 27829 28491 27863
rect 30205 27829 30239 27863
rect 31217 27829 31251 27863
rect 31585 27829 31619 27863
rect 32873 27829 32907 27863
rect 8309 27625 8343 27659
rect 14920 27625 14954 27659
rect 25684 27625 25718 27659
rect 30389 27625 30423 27659
rect 37289 27625 37323 27659
rect 21741 27557 21775 27591
rect 24409 27557 24443 27591
rect 9413 27489 9447 27523
rect 23213 27489 23247 27523
rect 27169 27489 27203 27523
rect 28365 27489 28399 27523
rect 32229 27489 32263 27523
rect 8217 27421 8251 27455
rect 8953 27421 8987 27455
rect 14657 27421 14691 27455
rect 16865 27421 16899 27455
rect 19533 27421 19567 27455
rect 19625 27421 19659 27455
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 21005 27421 21039 27455
rect 21097 27399 21131 27433
rect 21741 27421 21775 27455
rect 21925 27421 21959 27455
rect 22937 27421 22971 27455
rect 23029 27421 23063 27455
rect 24685 27421 24719 27455
rect 25421 27421 25455 27455
rect 28089 27421 28123 27455
rect 28181 27421 28215 27455
rect 28457 27421 28491 27455
rect 30205 27421 30239 27455
rect 9137 27353 9171 27387
rect 13369 27353 13403 27387
rect 17049 27353 17083 27387
rect 18705 27353 18739 27387
rect 20821 27353 20855 27387
rect 23213 27353 23247 27387
rect 24409 27353 24443 27387
rect 24593 27353 24627 27387
rect 30021 27353 30055 27387
rect 32505 27353 32539 27387
rect 13461 27285 13495 27319
rect 16405 27285 16439 27319
rect 19257 27285 19291 27319
rect 20913 27285 20947 27319
rect 27905 27285 27939 27319
rect 33977 27285 34011 27319
rect 8309 27081 8343 27115
rect 14289 27081 14323 27115
rect 14473 27081 14507 27115
rect 15945 27081 15979 27115
rect 17141 27081 17175 27115
rect 13921 27013 13955 27047
rect 14933 27013 14967 27047
rect 15133 27013 15167 27047
rect 18889 27013 18923 27047
rect 22293 27013 22327 27047
rect 22477 27013 22511 27047
rect 27077 27013 27111 27047
rect 28181 27013 28215 27047
rect 32873 27013 32907 27047
rect 8217 26945 8251 26979
rect 9045 26945 9079 26979
rect 14105 26945 14139 26979
rect 14197 26945 14231 26979
rect 15761 26945 15795 26979
rect 17049 26945 17083 26979
rect 22109 26945 22143 26979
rect 22937 26945 22971 26979
rect 23213 26945 23247 26979
rect 26985 26945 27019 26979
rect 32137 26945 32171 26979
rect 32321 26945 32355 26979
rect 32413 26945 32447 26979
rect 32689 26945 32723 26979
rect 11529 26877 11563 26911
rect 11805 26877 11839 26911
rect 18613 26877 18647 26911
rect 23029 26877 23063 26911
rect 27905 26877 27939 26911
rect 29653 26877 29687 26911
rect 32505 26877 32539 26911
rect 15301 26809 15335 26843
rect 23397 26809 23431 26843
rect 8861 26741 8895 26775
rect 13277 26741 13311 26775
rect 15117 26741 15151 26775
rect 20361 26741 20395 26775
rect 22937 26741 22971 26775
rect 11713 26537 11747 26571
rect 29653 26537 29687 26571
rect 30389 26537 30423 26571
rect 31125 26537 31159 26571
rect 16129 26469 16163 26503
rect 16681 26469 16715 26503
rect 19901 26469 19935 26503
rect 21741 26469 21775 26503
rect 27905 26469 27939 26503
rect 8953 26401 8987 26435
rect 11529 26401 11563 26435
rect 12725 26401 12759 26435
rect 21189 26401 21223 26435
rect 22569 26401 22603 26435
rect 22845 26401 22879 26435
rect 24593 26401 24627 26435
rect 28365 26401 28399 26435
rect 28549 26401 28583 26435
rect 32137 26401 32171 26435
rect 11437 26333 11471 26367
rect 13001 26333 13035 26367
rect 14381 26333 14415 26367
rect 16589 26333 16623 26367
rect 19809 26333 19843 26367
rect 21097 26333 21131 26367
rect 21281 26333 21315 26367
rect 21741 26333 21775 26367
rect 22017 26333 22051 26367
rect 24777 26333 24811 26367
rect 25421 26333 25455 26367
rect 25605 26333 25639 26367
rect 27169 26333 27203 26367
rect 27353 26333 27387 26367
rect 27445 26333 27479 26367
rect 29561 26333 29595 26367
rect 30205 26333 30239 26367
rect 30941 26333 30975 26367
rect 31769 26333 31803 26367
rect 31953 26333 31987 26367
rect 32045 26333 32079 26367
rect 32321 26333 32355 26367
rect 9229 26265 9263 26299
rect 14657 26265 14691 26299
rect 21925 26265 21959 26299
rect 26985 26265 27019 26299
rect 28273 26265 28307 26299
rect 10701 26197 10735 26231
rect 24961 26197 24995 26231
rect 25513 26197 25547 26231
rect 32505 26197 32539 26231
rect 8861 25993 8895 26027
rect 10057 25993 10091 26027
rect 11621 25993 11655 26027
rect 12817 25993 12851 26027
rect 13737 25993 13771 26027
rect 13829 25993 13863 26027
rect 14013 25993 14047 26027
rect 14749 25993 14783 26027
rect 15853 25993 15887 26027
rect 31401 25993 31435 26027
rect 11713 25925 11747 25959
rect 12357 25925 12391 25959
rect 14841 25925 14875 25959
rect 21189 25925 21223 25959
rect 32505 25925 32539 25959
rect 8493 25857 8527 25891
rect 9965 25857 9999 25891
rect 11529 25857 11563 25891
rect 11805 25857 11839 25891
rect 12541 25857 12575 25891
rect 12909 25857 12943 25891
rect 13645 25857 13679 25891
rect 14473 25857 14507 25891
rect 14933 25857 14967 25891
rect 15761 25857 15795 25891
rect 21097 25857 21131 25891
rect 24685 25857 24719 25891
rect 24869 25857 24903 25891
rect 24961 25857 24995 25891
rect 25237 25857 25271 25891
rect 25881 25857 25915 25891
rect 26065 25857 26099 25891
rect 26985 25857 27019 25891
rect 28733 25857 28767 25891
rect 30113 25857 30147 25891
rect 30849 25857 30883 25891
rect 31125 25857 31159 25891
rect 8585 25789 8619 25823
rect 12633 25789 12667 25823
rect 13001 25789 13035 25823
rect 16681 25789 16715 25823
rect 16865 25789 16899 25823
rect 18521 25789 18555 25823
rect 21833 25789 21867 25823
rect 22109 25789 22143 25823
rect 23581 25789 23615 25823
rect 25053 25789 25087 25823
rect 32229 25789 32263 25823
rect 13461 25721 13495 25755
rect 26249 25721 26283 25755
rect 28917 25721 28951 25755
rect 30297 25721 30331 25755
rect 25421 25653 25455 25687
rect 25973 25653 26007 25687
rect 27077 25653 27111 25687
rect 31217 25653 31251 25687
rect 33977 25653 34011 25687
rect 47777 25653 47811 25687
rect 11437 25449 11471 25483
rect 12449 25449 12483 25483
rect 14381 25449 14415 25483
rect 16865 25449 16899 25483
rect 22109 25449 22143 25483
rect 27813 25449 27847 25483
rect 30665 25449 30699 25483
rect 30849 25449 30883 25483
rect 31401 25449 31435 25483
rect 33241 25449 33275 25483
rect 27077 25381 27111 25415
rect 9505 25313 9539 25347
rect 25605 25313 25639 25347
rect 46305 25313 46339 25347
rect 1409 25245 1443 25279
rect 9229 25245 9263 25279
rect 9413 25245 9447 25279
rect 9965 25245 9999 25279
rect 10609 25245 10643 25279
rect 10793 25245 10827 25279
rect 11345 25245 11379 25279
rect 12357 25245 12391 25279
rect 14381 25245 14415 25279
rect 16773 25245 16807 25279
rect 17693 25245 17727 25279
rect 18337 25245 18371 25279
rect 18521 25245 18555 25279
rect 19257 25245 19291 25279
rect 21465 25245 21499 25279
rect 21558 25245 21592 25279
rect 21741 25245 21775 25279
rect 21930 25245 21964 25279
rect 24685 25245 24719 25279
rect 25329 25245 25363 25279
rect 29561 25245 29595 25279
rect 29745 25245 29779 25279
rect 30573 25245 30607 25279
rect 30665 25245 30699 25279
rect 31585 25245 31619 25279
rect 31769 25245 31803 25279
rect 31861 25245 31895 25279
rect 33149 25245 33183 25279
rect 1685 25177 1719 25211
rect 10701 25177 10735 25211
rect 18429 25177 18463 25211
rect 21833 25177 21867 25211
rect 27721 25177 27755 25211
rect 30389 25177 30423 25211
rect 46489 25177 46523 25211
rect 48145 25177 48179 25211
rect 9045 25109 9079 25143
rect 10057 25109 10091 25143
rect 17785 25109 17819 25143
rect 19349 25109 19383 25143
rect 24777 25109 24811 25143
rect 29929 25109 29963 25143
rect 24041 24905 24075 24939
rect 27169 24905 27203 24939
rect 28457 24905 28491 24939
rect 14381 24837 14415 24871
rect 24409 24837 24443 24871
rect 24527 24837 24561 24871
rect 25513 24837 25547 24871
rect 26341 24837 26375 24871
rect 7757 24769 7791 24803
rect 10241 24769 10275 24803
rect 12633 24769 12667 24803
rect 12817 24769 12851 24803
rect 14013 24769 14047 24803
rect 22661 24769 22695 24803
rect 24225 24769 24259 24803
rect 24317 24769 24351 24803
rect 24685 24769 24719 24803
rect 25329 24769 25363 24803
rect 25605 24769 25639 24803
rect 26065 24769 26099 24803
rect 26985 24769 27019 24803
rect 28273 24769 28307 24803
rect 29745 24769 29779 24803
rect 29837 24769 29871 24803
rect 30113 24769 30147 24803
rect 30849 24769 30883 24803
rect 32229 24769 32263 24803
rect 46857 24769 46891 24803
rect 47593 24769 47627 24803
rect 47685 24769 47719 24803
rect 7941 24701 7975 24735
rect 8309 24701 8343 24735
rect 16773 24701 16807 24735
rect 17049 24701 17083 24735
rect 18981 24701 19015 24735
rect 19257 24701 19291 24735
rect 26157 24701 26191 24735
rect 26341 24701 26375 24735
rect 29561 24701 29595 24735
rect 31125 24701 31159 24735
rect 10057 24565 10091 24599
rect 12725 24565 12759 24599
rect 18521 24565 18555 24599
rect 20729 24565 20763 24599
rect 22845 24565 22879 24599
rect 25145 24565 25179 24599
rect 30021 24565 30055 24599
rect 30665 24565 30699 24599
rect 31033 24565 31067 24599
rect 32321 24565 32355 24599
rect 46949 24565 46983 24599
rect 8217 24361 8251 24395
rect 10701 24361 10735 24395
rect 11713 24361 11747 24395
rect 19257 24361 19291 24395
rect 20637 24361 20671 24395
rect 26157 24361 26191 24395
rect 28733 24361 28767 24395
rect 30573 24361 30607 24395
rect 32873 24361 32907 24395
rect 11161 24293 11195 24327
rect 8953 24225 8987 24259
rect 9229 24225 9263 24259
rect 12633 24225 12667 24259
rect 14289 24225 14323 24259
rect 17417 24225 17451 24259
rect 20085 24225 20119 24259
rect 24409 24225 24443 24259
rect 27261 24225 27295 24259
rect 30205 24225 30239 24259
rect 31125 24225 31159 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 8125 24157 8159 24191
rect 11437 24157 11471 24191
rect 12725 24157 12759 24191
rect 14565 24157 14599 24191
rect 15577 24157 15611 24191
rect 18153 24157 18187 24191
rect 18337 24157 18371 24191
rect 19349 24157 19383 24191
rect 19993 24157 20027 24191
rect 20177 24157 20211 24191
rect 20637 24157 20671 24191
rect 20821 24157 20855 24191
rect 26985 24157 27019 24191
rect 30297 24157 30331 24191
rect 46305 24157 46339 24191
rect 15761 24089 15795 24123
rect 18521 24089 18555 24123
rect 24685 24089 24719 24123
rect 31401 24089 31435 24123
rect 11345 24021 11379 24055
rect 11529 24021 11563 24055
rect 13093 24021 13127 24055
rect 1961 23817 1995 23851
rect 14933 23817 14967 23851
rect 15761 23817 15795 23851
rect 17049 23817 17083 23851
rect 17877 23817 17911 23851
rect 18905 23817 18939 23851
rect 19073 23817 19107 23851
rect 26341 23817 26375 23851
rect 11713 23749 11747 23783
rect 13461 23749 13495 23783
rect 18705 23749 18739 23783
rect 24133 23749 24167 23783
rect 1869 23681 1903 23715
rect 9321 23681 9355 23715
rect 9505 23681 9539 23715
rect 9965 23681 9999 23715
rect 10609 23681 10643 23715
rect 10701 23681 10735 23715
rect 10977 23681 11011 23715
rect 11805 23681 11839 23715
rect 11897 23681 11931 23715
rect 15577 23681 15611 23715
rect 17049 23681 17083 23715
rect 17785 23681 17819 23715
rect 17969 23681 18003 23715
rect 19625 23681 19659 23715
rect 19717 23681 19751 23715
rect 20453 23681 20487 23715
rect 22293 23681 22327 23715
rect 24685 23681 24719 23715
rect 25605 23681 25639 23715
rect 26249 23681 26283 23715
rect 28181 23681 28215 23715
rect 30573 23681 30607 23715
rect 30665 23681 30699 23715
rect 30941 23681 30975 23715
rect 31401 23681 31435 23715
rect 31585 23681 31619 23715
rect 47777 23681 47811 23715
rect 10793 23613 10827 23647
rect 13185 23613 13219 23647
rect 22477 23613 22511 23647
rect 28457 23613 28491 23647
rect 29929 23613 29963 23647
rect 46213 23613 46247 23647
rect 46489 23613 46523 23647
rect 10977 23545 11011 23579
rect 11529 23545 11563 23579
rect 24869 23545 24903 23579
rect 9321 23477 9355 23511
rect 10057 23477 10091 23511
rect 12081 23477 12115 23511
rect 18889 23477 18923 23511
rect 19901 23477 19935 23511
rect 20637 23477 20671 23511
rect 25697 23477 25731 23511
rect 30389 23477 30423 23511
rect 30849 23477 30883 23511
rect 31493 23477 31527 23511
rect 13093 23273 13127 23307
rect 15761 23273 15795 23307
rect 19809 23273 19843 23307
rect 23029 23273 23063 23307
rect 27997 23273 28031 23307
rect 28641 23273 28675 23307
rect 29561 23273 29595 23307
rect 30573 23273 30607 23307
rect 29929 23205 29963 23239
rect 9781 23137 9815 23171
rect 19257 23137 19291 23171
rect 25329 23137 25363 23171
rect 45017 23137 45051 23171
rect 46857 23137 46891 23171
rect 9505 23069 9539 23103
rect 13001 23069 13035 23103
rect 14105 23069 14139 23103
rect 15669 23069 15703 23103
rect 16957 23069 16991 23103
rect 17601 23069 17635 23103
rect 19533 23069 19567 23103
rect 20729 23069 20763 23103
rect 22937 23069 22971 23103
rect 25053 23069 25087 23103
rect 26249 23069 26283 23103
rect 27077 23069 27111 23103
rect 27905 23069 27939 23103
rect 28549 23069 28583 23103
rect 29745 23069 29779 23103
rect 30021 23069 30055 23103
rect 30481 23069 30515 23103
rect 30665 23069 30699 23103
rect 45293 23069 45327 23103
rect 46305 23069 46339 23103
rect 19625 23001 19659 23035
rect 21005 23001 21039 23035
rect 26617 23001 26651 23035
rect 46489 23001 46523 23035
rect 11253 22933 11287 22967
rect 14289 22933 14323 22967
rect 16957 22933 16991 22967
rect 17693 22933 17727 22967
rect 19441 22933 19475 22967
rect 22477 22933 22511 22967
rect 27169 22933 27203 22967
rect 9781 22729 9815 22763
rect 14013 22729 14047 22763
rect 20821 22729 20855 22763
rect 21925 22729 21959 22763
rect 47685 22729 47719 22763
rect 19901 22661 19935 22695
rect 24869 22661 24903 22695
rect 27169 22661 27203 22695
rect 45385 22661 45419 22695
rect 9689 22593 9723 22627
rect 12633 22593 12667 22627
rect 13921 22593 13955 22627
rect 15025 22593 15059 22627
rect 16681 22593 16715 22627
rect 19073 22593 19107 22627
rect 20085 22593 20119 22627
rect 20177 22593 20211 22627
rect 20821 22593 20855 22627
rect 21833 22593 21867 22627
rect 22017 22593 22051 22627
rect 23029 22593 23063 22627
rect 25329 22593 25363 22627
rect 43453 22593 43487 22627
rect 43729 22593 43763 22627
rect 47593 22593 47627 22627
rect 12725 22525 12759 22559
rect 16957 22525 16991 22559
rect 18429 22525 18463 22559
rect 19165 22525 19199 22559
rect 23213 22525 23247 22559
rect 25697 22525 25731 22559
rect 26985 22525 27019 22559
rect 27629 22525 27663 22559
rect 44281 22525 44315 22559
rect 45201 22525 45235 22559
rect 46581 22525 46615 22559
rect 19441 22457 19475 22491
rect 19901 22457 19935 22491
rect 13001 22389 13035 22423
rect 15117 22389 15151 22423
rect 23213 22185 23247 22219
rect 10885 22049 10919 22083
rect 15025 22049 15059 22083
rect 26065 22049 26099 22083
rect 45293 22049 45327 22083
rect 46857 22049 46891 22083
rect 14841 21981 14875 22015
rect 16681 21981 16715 22015
rect 19257 21981 19291 22015
rect 21557 21981 21591 22015
rect 23121 21981 23155 22015
rect 25053 21981 25087 22015
rect 25881 21981 25915 22015
rect 44189 21981 44223 22015
rect 44281 21981 44315 22015
rect 45017 21981 45051 22015
rect 46305 21981 46339 22015
rect 11069 21913 11103 21947
rect 12725 21913 12759 21947
rect 19441 21913 19475 21947
rect 21097 21913 21131 21947
rect 27721 21913 27755 21947
rect 46489 21913 46523 21947
rect 21649 21845 21683 21879
rect 25145 21845 25179 21879
rect 43821 21845 43855 21879
rect 44465 21845 44499 21879
rect 15393 21641 15427 21675
rect 21925 21641 21959 21675
rect 47685 21641 47719 21675
rect 13277 21573 13311 21607
rect 25697 21573 25731 21607
rect 42901 21573 42935 21607
rect 7941 21505 7975 21539
rect 10425 21505 10459 21539
rect 11529 21505 11563 21539
rect 12173 21505 12207 21539
rect 12357 21505 12391 21539
rect 15301 21505 15335 21539
rect 17969 21505 18003 21539
rect 20269 21505 20303 21539
rect 21833 21505 21867 21539
rect 23121 21505 23155 21539
rect 26157 21505 26191 21539
rect 42809 21505 42843 21539
rect 42993 21505 43027 21539
rect 44465 21505 44499 21539
rect 44557 21505 44591 21539
rect 45937 21505 45971 21539
rect 46121 21505 46155 21539
rect 47593 21505 47627 21539
rect 8125 21437 8159 21471
rect 9137 21437 9171 21471
rect 13001 21437 13035 21471
rect 14749 21437 14783 21471
rect 18153 21437 18187 21471
rect 18429 21437 18463 21471
rect 23857 21437 23891 21471
rect 24041 21437 24075 21471
rect 46857 21437 46891 21471
rect 20361 21369 20395 21403
rect 44741 21369 44775 21403
rect 10241 21301 10275 21335
rect 11621 21301 11655 21335
rect 12173 21301 12207 21335
rect 23305 21301 23339 21335
rect 26341 21301 26375 21335
rect 9045 21097 9079 21131
rect 11989 21097 12023 21131
rect 13093 21097 13127 21131
rect 19349 21097 19383 21131
rect 23765 21097 23799 21131
rect 43729 21097 43763 21131
rect 45661 21097 45695 21131
rect 20913 21029 20947 21063
rect 23121 21029 23155 21063
rect 10241 20961 10275 20995
rect 10517 20961 10551 20995
rect 20453 20961 20487 20995
rect 21373 20961 21407 20995
rect 21649 20961 21683 20995
rect 26617 20961 26651 20995
rect 29745 20961 29779 20995
rect 48145 20961 48179 20995
rect 8953 20893 8987 20927
rect 9597 20893 9631 20927
rect 13093 20893 13127 20927
rect 14105 20893 14139 20927
rect 16773 20893 16807 20927
rect 19257 20893 19291 20927
rect 20545 20893 20579 20927
rect 23673 20893 23707 20927
rect 24777 20893 24811 20927
rect 26157 20893 26191 20927
rect 29561 20893 29595 20927
rect 43637 20893 43671 20927
rect 43821 20893 43855 20927
rect 44281 20893 44315 20927
rect 44465 20893 44499 20927
rect 45293 20893 45327 20927
rect 46305 20893 46339 20927
rect 25421 20825 25455 20859
rect 26341 20825 26375 20859
rect 31401 20825 31435 20859
rect 45477 20825 45511 20859
rect 46489 20825 46523 20859
rect 9689 20757 9723 20791
rect 14289 20757 14323 20791
rect 16865 20757 16899 20791
rect 44465 20757 44499 20791
rect 13093 20553 13127 20587
rect 13921 20553 13955 20587
rect 20177 20553 20211 20587
rect 22109 20553 22143 20587
rect 27077 20553 27111 20587
rect 47685 20553 47719 20587
rect 7481 20485 7515 20519
rect 8217 20485 8251 20519
rect 11529 20485 11563 20519
rect 12725 20485 12759 20519
rect 12941 20485 12975 20519
rect 16865 20485 16899 20519
rect 19993 20485 20027 20519
rect 27813 20485 27847 20519
rect 45385 20485 45419 20519
rect 7389 20417 7423 20451
rect 11713 20417 11747 20451
rect 11805 20417 11839 20451
rect 13829 20417 13863 20451
rect 15761 20417 15795 20451
rect 20085 20417 20119 20451
rect 22017 20417 22051 20451
rect 23489 20417 23523 20451
rect 24777 20417 24811 20451
rect 26157 20417 26191 20451
rect 26249 20417 26283 20451
rect 26985 20417 27019 20451
rect 30389 20417 30423 20451
rect 39129 20417 39163 20451
rect 47593 20417 47627 20451
rect 8033 20349 8067 20383
rect 8585 20349 8619 20383
rect 16681 20349 16715 20383
rect 17141 20349 17175 20383
rect 23765 20349 23799 20383
rect 24961 20349 24995 20383
rect 27629 20349 27663 20383
rect 29009 20349 29043 20383
rect 39313 20349 39347 20383
rect 39589 20349 39623 20383
rect 44281 20349 44315 20383
rect 45201 20349 45235 20383
rect 47041 20349 47075 20383
rect 11529 20281 11563 20315
rect 19809 20281 19843 20315
rect 44557 20281 44591 20315
rect 12909 20213 12943 20247
rect 15945 20213 15979 20247
rect 20361 20213 20395 20247
rect 26433 20213 26467 20247
rect 30481 20213 30515 20247
rect 44741 20213 44775 20247
rect 9768 20009 9802 20043
rect 11713 20009 11747 20043
rect 26617 20009 26651 20043
rect 11253 19873 11287 19907
rect 19533 19873 19567 19907
rect 30481 19873 30515 19907
rect 40601 19873 40635 19907
rect 44373 19873 44407 19907
rect 45477 19873 45511 19907
rect 45569 19873 45603 19907
rect 46489 19873 46523 19907
rect 2053 19805 2087 19839
rect 9505 19805 9539 19839
rect 11894 19805 11928 19839
rect 12265 19805 12299 19839
rect 12357 19805 12391 19839
rect 14105 19805 14139 19839
rect 15301 19805 15335 19839
rect 17785 19805 17819 19839
rect 19257 19805 19291 19839
rect 21557 19805 21591 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 25145 19805 25179 19839
rect 26249 19805 26283 19839
rect 26433 19805 26467 19839
rect 27445 19805 27479 19839
rect 27629 19805 27663 19839
rect 28273 19805 28307 19839
rect 30297 19805 30331 19839
rect 43821 19805 43855 19839
rect 44097 19805 44131 19839
rect 45017 19805 45051 19839
rect 45201 19805 45235 19839
rect 46305 19805 46339 19839
rect 15577 19737 15611 19771
rect 25513 19737 25547 19771
rect 27721 19737 27755 19771
rect 32137 19737 32171 19771
rect 40785 19737 40819 19771
rect 42441 19737 42475 19771
rect 48145 19737 48179 19771
rect 11897 19669 11931 19703
rect 14289 19669 14323 19703
rect 17049 19669 17083 19703
rect 17877 19669 17911 19703
rect 21005 19669 21039 19703
rect 21649 19669 21683 19703
rect 24593 19669 24627 19703
rect 28365 19669 28399 19703
rect 10885 19465 10919 19499
rect 11897 19465 11931 19499
rect 16773 19465 16807 19499
rect 21189 19465 21223 19499
rect 28089 19465 28123 19499
rect 40785 19465 40819 19499
rect 11529 19397 11563 19431
rect 11745 19397 11779 19431
rect 17877 19397 17911 19431
rect 21833 19397 21867 19431
rect 23029 19397 23063 19431
rect 22063 19363 22097 19397
rect 1777 19329 1811 19363
rect 10793 19329 10827 19363
rect 12357 19329 12391 19363
rect 12541 19329 12575 19363
rect 15761 19329 15795 19363
rect 16681 19329 16715 19363
rect 17693 19329 17727 19363
rect 20170 19329 20204 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 25237 19329 25271 19363
rect 25329 19329 25363 19363
rect 25973 19329 26007 19363
rect 27721 19329 27755 19363
rect 28641 19329 28675 19363
rect 28917 19329 28951 19363
rect 29745 19329 29779 19363
rect 40693 19329 40727 19363
rect 43913 19329 43947 19363
rect 44097 19329 44131 19363
rect 45017 19329 45051 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 15853 19261 15887 19295
rect 18245 19261 18279 19295
rect 20269 19261 20303 19295
rect 20545 19261 20579 19295
rect 22937 19261 22971 19295
rect 23765 19261 23799 19295
rect 26065 19261 26099 19295
rect 26341 19261 26375 19295
rect 27813 19261 27847 19295
rect 29377 19261 29411 19295
rect 44005 19261 44039 19295
rect 44741 19261 44775 19295
rect 45569 19261 45603 19295
rect 47777 19261 47811 19295
rect 16129 19193 16163 19227
rect 22201 19193 22235 19227
rect 30021 19193 30055 19227
rect 11713 19125 11747 19159
rect 12357 19125 12391 19159
rect 21005 19125 21039 19159
rect 22017 19125 22051 19159
rect 47041 19125 47075 19159
rect 2329 18921 2363 18955
rect 11989 18921 12023 18955
rect 12173 18921 12207 18955
rect 14289 18921 14323 18955
rect 15761 18921 15795 18955
rect 19441 18921 19475 18955
rect 22293 18921 22327 18955
rect 27997 18921 28031 18955
rect 31953 18921 31987 18955
rect 44281 18921 44315 18955
rect 14473 18853 14507 18887
rect 23857 18853 23891 18887
rect 27813 18853 27847 18887
rect 43361 18853 43395 18887
rect 45109 18853 45143 18887
rect 12909 18785 12943 18819
rect 23489 18785 23523 18819
rect 26065 18785 26099 18819
rect 28457 18785 28491 18819
rect 46305 18785 46339 18819
rect 48145 18785 48179 18819
rect 2237 18717 2271 18751
rect 11069 18717 11103 18751
rect 13369 18717 13403 18751
rect 14933 18717 14967 18751
rect 15669 18717 15703 18751
rect 17601 18717 17635 18751
rect 19349 18717 19383 18751
rect 20545 18717 20579 18751
rect 23673 18717 23707 18751
rect 24501 18717 24535 18751
rect 26157 18717 26191 18751
rect 27537 18717 27571 18751
rect 28641 18717 28675 18751
rect 28917 18717 28951 18751
rect 30113 18717 30147 18751
rect 31033 18717 31067 18751
rect 43269 18717 43303 18751
rect 43545 18717 43579 18751
rect 44189 18717 44223 18751
rect 44373 18717 44407 18751
rect 45017 18717 45051 18751
rect 45201 18717 45235 18751
rect 11805 18649 11839 18683
rect 12021 18649 12055 18683
rect 12725 18649 12759 18683
rect 14105 18649 14139 18683
rect 18245 18649 18279 18683
rect 20821 18649 20855 18683
rect 25237 18649 25271 18683
rect 29009 18649 29043 18683
rect 46489 18649 46523 18683
rect 11161 18581 11195 18615
rect 13461 18581 13495 18615
rect 14305 18581 14339 18615
rect 15117 18581 15151 18615
rect 26525 18581 26559 18615
rect 1961 18377 1995 18411
rect 19901 18377 19935 18411
rect 20545 18377 20579 18411
rect 47685 18377 47719 18411
rect 12909 18309 12943 18343
rect 16037 18309 16071 18343
rect 16865 18309 16899 18343
rect 27629 18309 27663 18343
rect 46305 18309 46339 18343
rect 1869 18241 1903 18275
rect 11713 18241 11747 18275
rect 11897 18241 11931 18275
rect 11989 18241 12023 18275
rect 15945 18241 15979 18275
rect 16681 18241 16715 18275
rect 19073 18241 19107 18275
rect 19809 18241 19843 18275
rect 20453 18241 20487 18275
rect 20637 18241 20671 18275
rect 23305 18241 23339 18275
rect 25789 18241 25823 18275
rect 27353 18241 27387 18275
rect 27445 18241 27479 18275
rect 28089 18241 28123 18275
rect 44189 18241 44223 18275
rect 44649 18241 44683 18275
rect 44925 18241 44959 18275
rect 45937 18241 45971 18275
rect 46121 18241 46155 18275
rect 47041 18241 47075 18275
rect 47593 18241 47627 18275
rect 8585 18173 8619 18207
rect 8769 18173 8803 18207
rect 9045 18173 9079 18207
rect 12633 18173 12667 18207
rect 14381 18173 14415 18207
rect 18521 18173 18555 18207
rect 19165 18173 19199 18207
rect 23489 18173 23523 18207
rect 25145 18173 25179 18207
rect 28273 18173 28307 18207
rect 29929 18173 29963 18207
rect 45293 18173 45327 18207
rect 11713 18105 11747 18139
rect 45385 18105 45419 18139
rect 25881 18037 25915 18071
rect 46857 18037 46891 18071
rect 12633 17833 12667 17867
rect 16681 17833 16715 17867
rect 23489 17833 23523 17867
rect 28089 17833 28123 17867
rect 44465 17833 44499 17867
rect 45293 17833 45327 17867
rect 8309 17765 8343 17799
rect 9045 17697 9079 17731
rect 9505 17697 9539 17731
rect 10241 17697 10275 17731
rect 17969 17697 18003 17731
rect 25878 17697 25912 17731
rect 26157 17697 26191 17731
rect 2145 17629 2179 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 9965 17629 9999 17663
rect 12633 17629 12667 17663
rect 14105 17629 14139 17663
rect 16589 17629 16623 17663
rect 17509 17629 17543 17663
rect 19257 17629 19291 17663
rect 19993 17629 20027 17663
rect 20821 17629 20855 17663
rect 20913 17629 20947 17663
rect 21465 17629 21499 17663
rect 22293 17629 22327 17663
rect 23397 17629 23431 17663
rect 25697 17629 25731 17663
rect 27997 17629 28031 17663
rect 44097 17629 44131 17663
rect 44281 17629 44315 17663
rect 45017 17629 45051 17663
rect 46305 17629 46339 17663
rect 45201 17561 45235 17595
rect 46489 17561 46523 17595
rect 48145 17561 48179 17595
rect 2237 17493 2271 17527
rect 11713 17493 11747 17527
rect 14289 17493 14323 17527
rect 19441 17493 19475 17527
rect 20177 17493 20211 17527
rect 21649 17493 21683 17527
rect 22385 17493 22419 17527
rect 10609 17289 10643 17323
rect 44373 17289 44407 17323
rect 47685 17289 47719 17323
rect 1961 17221 1995 17255
rect 23029 17221 23063 17255
rect 7941 17153 7975 17187
rect 10517 17153 10551 17187
rect 14197 17153 14231 17187
rect 14933 17153 14967 17187
rect 15669 17153 15703 17187
rect 16773 17153 16807 17187
rect 17601 17153 17635 17187
rect 22017 17153 22051 17187
rect 26985 17153 27019 17187
rect 44281 17153 44315 17187
rect 44465 17153 44499 17187
rect 47041 17153 47075 17187
rect 47593 17153 47627 17187
rect 1777 17085 1811 17119
rect 2789 17085 2823 17119
rect 8125 17085 8159 17119
rect 8401 17085 8435 17119
rect 17785 17085 17819 17119
rect 19257 17085 19291 17119
rect 19533 17085 19567 17119
rect 21281 17085 21315 17119
rect 22845 17085 22879 17119
rect 24685 17085 24719 17119
rect 27169 17085 27203 17119
rect 28825 17085 28859 17119
rect 14381 16949 14415 16983
rect 14933 16949 14967 16983
rect 15761 16949 15795 16983
rect 16865 16949 16899 16983
rect 21833 16949 21867 16983
rect 2053 16745 2087 16779
rect 8217 16745 8251 16779
rect 13553 16745 13587 16779
rect 14657 16609 14691 16643
rect 14933 16609 14967 16643
rect 16405 16609 16439 16643
rect 16865 16609 16899 16643
rect 17049 16609 17083 16643
rect 46305 16609 46339 16643
rect 8125 16541 8159 16575
rect 11253 16541 11287 16575
rect 11989 16541 12023 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 13001 16541 13035 16575
rect 19257 16541 19291 16575
rect 20821 16541 20855 16575
rect 21925 16541 21959 16575
rect 22661 16541 22695 16575
rect 27353 16541 27387 16575
rect 11345 16473 11379 16507
rect 18705 16473 18739 16507
rect 20085 16473 20119 16507
rect 21373 16473 21407 16507
rect 46489 16473 46523 16507
rect 48145 16473 48179 16507
rect 11805 16405 11839 16439
rect 13185 16405 13219 16439
rect 13277 16405 13311 16439
rect 13369 16405 13403 16439
rect 22109 16405 22143 16439
rect 22753 16405 22787 16439
rect 27537 16405 27571 16439
rect 13277 16201 13311 16235
rect 46765 16201 46799 16235
rect 11805 16133 11839 16167
rect 13829 16133 13863 16167
rect 17141 16133 17175 16167
rect 17877 16133 17911 16167
rect 22109 16133 22143 16167
rect 11529 16065 11563 16099
rect 13737 16065 13771 16099
rect 14381 16065 14415 16099
rect 17049 16065 17083 16099
rect 19993 16065 20027 16099
rect 21833 16065 21867 16099
rect 24041 16065 24075 16099
rect 25421 16065 25455 16099
rect 46673 16065 46707 16099
rect 47777 16065 47811 16099
rect 14657 15997 14691 16031
rect 16129 15997 16163 16031
rect 17693 15997 17727 16031
rect 19533 15997 19567 16031
rect 20361 15997 20395 16031
rect 23581 15861 23615 15895
rect 24133 15861 24167 15895
rect 25513 15861 25547 15895
rect 13369 15657 13403 15691
rect 15945 15657 15979 15691
rect 20269 15657 20303 15691
rect 14657 15589 14691 15623
rect 15117 15589 15151 15623
rect 14105 15521 14139 15555
rect 22017 15521 22051 15555
rect 25513 15521 25547 15555
rect 27169 15521 27203 15555
rect 2053 15453 2087 15487
rect 14289 15453 14323 15487
rect 15117 15453 15151 15487
rect 15393 15453 15427 15487
rect 15853 15453 15887 15487
rect 19441 15453 19475 15487
rect 20177 15453 20211 15487
rect 21097 15453 21131 15487
rect 22109 15453 22143 15487
rect 22937 15453 22971 15487
rect 25329 15453 25363 15487
rect 13185 15385 13219 15419
rect 14473 15385 14507 15419
rect 18245 15385 18279 15419
rect 21281 15385 21315 15419
rect 13385 15317 13419 15351
rect 13553 15317 13587 15351
rect 14381 15317 14415 15351
rect 15301 15317 15335 15351
rect 18337 15317 18371 15351
rect 19625 15317 19659 15351
rect 21465 15317 21499 15351
rect 22477 15317 22511 15351
rect 23029 15317 23063 15351
rect 15025 15113 15059 15147
rect 24409 15113 24443 15147
rect 21189 15045 21223 15079
rect 22937 15045 22971 15079
rect 1777 14977 1811 15011
rect 13185 14977 13219 15011
rect 13277 14977 13311 15011
rect 14105 14977 14139 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 18337 14977 18371 15011
rect 21097 14977 21131 15011
rect 21281 14977 21315 15011
rect 21833 14977 21867 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22661 14977 22695 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 14013 14909 14047 14943
rect 18613 14909 18647 14943
rect 14473 14841 14507 14875
rect 13461 14773 13495 14807
rect 2237 14569 2271 14603
rect 17877 14501 17911 14535
rect 20729 14433 20763 14467
rect 20913 14433 20947 14467
rect 2145 14365 2179 14399
rect 17509 14365 17543 14399
rect 20085 14365 20119 14399
rect 20821 14365 20855 14399
rect 21005 14365 21039 14399
rect 17325 14297 17359 14331
rect 17693 14297 17727 14331
rect 17601 14229 17635 14263
rect 19901 14229 19935 14263
rect 20545 14229 20579 14263
rect 17141 14025 17175 14059
rect 17877 14025 17911 14059
rect 18981 14025 19015 14059
rect 20177 14025 20211 14059
rect 22385 14025 22419 14059
rect 16773 13957 16807 13991
rect 16989 13957 17023 13991
rect 17969 13957 18003 13991
rect 18797 13957 18831 13991
rect 15853 13889 15887 13923
rect 17785 13889 17819 13923
rect 18889 13889 18923 13923
rect 20729 13889 20763 13923
rect 22201 13889 22235 13923
rect 17601 13821 17635 13855
rect 18153 13821 18187 13855
rect 18613 13821 18647 13855
rect 19165 13821 19199 13855
rect 19717 13821 19751 13855
rect 20085 13753 20119 13787
rect 16037 13685 16071 13719
rect 16957 13685 16991 13719
rect 20821 13685 20855 13719
rect 22109 13481 22143 13515
rect 19809 13413 19843 13447
rect 13277 13345 13311 13379
rect 13553 13345 13587 13379
rect 14381 13345 14415 13379
rect 19349 13345 19383 13379
rect 20361 13345 20395 13379
rect 13185 13277 13219 13311
rect 14105 13277 14139 13311
rect 16405 13277 16439 13311
rect 19441 13277 19475 13311
rect 16681 13209 16715 13243
rect 20637 13209 20671 13243
rect 15853 13141 15887 13175
rect 18153 13141 18187 13175
rect 14105 12937 14139 12971
rect 14749 12937 14783 12971
rect 16865 12937 16899 12971
rect 17601 12937 17635 12971
rect 18245 12937 18279 12971
rect 20913 12937 20947 12971
rect 21925 12937 21959 12971
rect 17417 12869 17451 12903
rect 1409 12801 1443 12835
rect 14105 12801 14139 12835
rect 14657 12801 14691 12835
rect 16681 12801 16715 12835
rect 17693 12801 17727 12835
rect 18153 12801 18187 12835
rect 19165 12801 19199 12835
rect 21833 12801 21867 12835
rect 19441 12733 19475 12767
rect 1593 12597 1627 12631
rect 17417 12597 17451 12631
rect 47777 12597 47811 12631
rect 16957 12393 16991 12427
rect 19533 12393 19567 12427
rect 20269 12393 20303 12427
rect 46305 12257 46339 12291
rect 48145 12257 48179 12291
rect 14749 12189 14783 12223
rect 16957 12189 16991 12223
rect 17141 12189 17175 12223
rect 19441 12189 19475 12223
rect 20177 12189 20211 12223
rect 46489 12121 46523 12155
rect 14841 12053 14875 12087
rect 47685 11849 47719 11883
rect 16773 11781 16807 11815
rect 16973 11781 17007 11815
rect 14197 11713 14231 11747
rect 15853 11713 15887 11747
rect 17601 11713 17635 11747
rect 47593 11713 47627 11747
rect 14013 11509 14047 11543
rect 16037 11509 16071 11543
rect 16957 11509 16991 11543
rect 17141 11509 17175 11543
rect 17693 11509 17727 11543
rect 16037 11169 16071 11203
rect 46305 11169 46339 11203
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 18245 11101 18279 11135
rect 19257 11101 19291 11135
rect 15485 11033 15519 11067
rect 16313 11033 16347 11067
rect 18337 11033 18371 11067
rect 19349 11033 19383 11067
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 14289 10965 14323 10999
rect 17785 10965 17819 10999
rect 15577 10761 15611 10795
rect 46857 10761 46891 10795
rect 14105 10693 14139 10727
rect 13829 10625 13863 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 46765 10625 46799 10659
rect 47777 10625 47811 10659
rect 17141 10557 17175 10591
rect 18153 10557 18187 10591
rect 17417 10489 17451 10523
rect 19625 10421 19659 10455
rect 46305 10421 46339 10455
rect 17693 10217 17727 10251
rect 15393 10081 15427 10115
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 17969 10013 18003 10047
rect 15577 9945 15611 9979
rect 17233 9945 17267 9979
rect 17693 9945 17727 9979
rect 17877 9945 17911 9979
rect 46489 9945 46523 9979
rect 16983 9673 17017 9707
rect 16773 9605 16807 9639
rect 18705 9605 18739 9639
rect 47685 9605 47719 9639
rect 17601 9537 17635 9571
rect 18889 9537 18923 9571
rect 19441 9537 19475 9571
rect 46213 9537 46247 9571
rect 47593 9537 47627 9571
rect 19625 9469 19659 9503
rect 21281 9469 21315 9503
rect 46489 9469 46523 9503
rect 17141 9401 17175 9435
rect 16957 9333 16991 9367
rect 17693 9333 17727 9367
rect 15485 9129 15519 9163
rect 19349 9129 19383 9163
rect 16589 8993 16623 9027
rect 18245 8993 18279 9027
rect 46489 8993 46523 9027
rect 46949 8993 46983 9027
rect 15393 8925 15427 8959
rect 19257 8925 19291 8959
rect 46305 8925 46339 8959
rect 16773 8857 16807 8891
rect 17233 8517 17267 8551
rect 47777 8517 47811 8551
rect 14197 8449 14231 8483
rect 19349 8449 19383 8483
rect 14381 8381 14415 8415
rect 14657 8381 14691 8415
rect 17049 8381 17083 8415
rect 17509 8381 17543 8415
rect 19441 8313 19475 8347
rect 47961 8313 47995 8347
rect 14381 8041 14415 8075
rect 16313 8041 16347 8075
rect 16865 7905 16899 7939
rect 17049 7905 17083 7939
rect 18061 7905 18095 7939
rect 46305 7905 46339 7939
rect 48053 7905 48087 7939
rect 14289 7837 14323 7871
rect 16221 7837 16255 7871
rect 46489 7769 46523 7803
rect 44833 7429 44867 7463
rect 17233 7361 17267 7395
rect 48145 7361 48179 7395
rect 17417 7293 17451 7327
rect 17969 7293 18003 7327
rect 44741 7293 44775 7327
rect 45201 7293 45235 7327
rect 47961 7225 47995 7259
rect 17509 6953 17543 6987
rect 47317 6817 47351 6851
rect 47593 6817 47627 6851
rect 17417 6749 17451 6783
rect 48145 6273 48179 6307
rect 47961 6069 47995 6103
rect 47317 5729 47351 5763
rect 20821 5661 20855 5695
rect 47593 5661 47627 5695
rect 20913 5525 20947 5559
rect 45477 5253 45511 5287
rect 45569 5253 45603 5287
rect 18613 5185 18647 5219
rect 19533 5185 19567 5219
rect 20177 5185 20211 5219
rect 20821 5185 20855 5219
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 47869 5185 47903 5219
rect 45753 5117 45787 5151
rect 18705 4981 18739 5015
rect 19625 4981 19659 5015
rect 20269 4981 20303 5015
rect 20913 4981 20947 5015
rect 21925 4981 21959 5015
rect 22569 4981 22603 5015
rect 48053 4981 48087 5015
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 21649 4777 21683 4811
rect 22293 4777 22327 4811
rect 15301 4641 15335 4675
rect 45845 4641 45879 4675
rect 47041 4641 47075 4675
rect 9505 4573 9539 4607
rect 18429 4573 18463 4607
rect 19257 4573 19291 4607
rect 20269 4573 20303 4607
rect 20913 4573 20947 4607
rect 21557 4573 21591 4607
rect 22201 4573 22235 4607
rect 22845 4573 22879 4607
rect 23489 4573 23523 4607
rect 39865 4573 39899 4607
rect 42717 4573 42751 4607
rect 45385 4573 45419 4607
rect 15485 4505 15519 4539
rect 17141 4505 17175 4539
rect 46029 4505 46063 4539
rect 18521 4437 18555 4471
rect 19349 4437 19383 4471
rect 22937 4437 22971 4471
rect 23581 4437 23615 4471
rect 39957 4437 39991 4471
rect 42809 4437 42843 4471
rect 18245 4233 18279 4267
rect 20177 4233 20211 4267
rect 22845 4233 22879 4267
rect 33241 4233 33275 4267
rect 39405 4233 39439 4267
rect 23673 4165 23707 4199
rect 24593 4165 24627 4199
rect 46673 4165 46707 4199
rect 47777 4165 47811 4199
rect 8493 4097 8527 4131
rect 9137 4097 9171 4131
rect 11529 4097 11563 4131
rect 13645 4097 13679 4131
rect 18153 4097 18187 4131
rect 18797 4097 18831 4131
rect 18889 4097 18923 4131
rect 19441 4097 19475 4131
rect 20085 4097 20119 4131
rect 21097 4097 21131 4131
rect 22753 4097 22787 4131
rect 25329 4097 25363 4131
rect 33149 4097 33183 4131
rect 39313 4097 39347 4131
rect 39957 4097 39991 4131
rect 41245 4097 41279 4131
rect 45937 4097 45971 4131
rect 1961 4029 1995 4063
rect 2145 4029 2179 4063
rect 2973 4029 3007 4063
rect 9321 4029 9355 4063
rect 10241 4029 10275 4063
rect 19533 4029 19567 4063
rect 21189 4029 21223 4063
rect 23581 4029 23615 4063
rect 29469 4029 29503 4063
rect 29653 4029 29687 4063
rect 31309 4029 31343 4063
rect 41061 4029 41095 4063
rect 43085 4029 43119 4063
rect 43269 4029 43303 4063
rect 44189 4029 44223 4063
rect 48053 4029 48087 4063
rect 46857 3961 46891 3995
rect 8585 3893 8619 3927
rect 11621 3893 11655 3927
rect 13737 3893 13771 3927
rect 22293 3893 22327 3927
rect 25421 3893 25455 3927
rect 40049 3893 40083 3927
rect 41705 3893 41739 3927
rect 42625 3893 42659 3927
rect 46029 3893 46063 3927
rect 2881 3689 2915 3723
rect 3985 3689 4019 3723
rect 10149 3689 10183 3723
rect 17233 3689 17267 3723
rect 19349 3689 19383 3723
rect 39221 3689 39255 3723
rect 10885 3553 10919 3587
rect 11161 3553 11195 3587
rect 27169 3553 27203 3587
rect 27353 3553 27387 3587
rect 27629 3553 27663 3587
rect 33241 3553 33275 3587
rect 39865 3553 39899 3587
rect 40325 3553 40359 3587
rect 42625 3553 42659 3587
rect 42809 3553 42843 3587
rect 43177 3553 43211 3587
rect 45201 3553 45235 3587
rect 46305 3553 46339 3587
rect 46489 3553 46523 3587
rect 1685 3485 1719 3519
rect 2145 3485 2179 3519
rect 2789 3485 2823 3519
rect 5273 3485 5307 3519
rect 5917 3485 5951 3519
rect 8217 3485 8251 3519
rect 9137 3485 9171 3519
rect 10057 3485 10091 3519
rect 10701 3485 10735 3519
rect 14289 3485 14323 3519
rect 17141 3485 17175 3519
rect 17785 3485 17819 3519
rect 18429 3485 18463 3519
rect 19257 3485 19291 3519
rect 20085 3485 20119 3519
rect 22385 3485 22419 3519
rect 23029 3485 23063 3519
rect 23121 3485 23155 3519
rect 23673 3485 23707 3519
rect 25145 3485 25179 3519
rect 35909 3485 35943 3519
rect 39129 3485 39163 3519
rect 45661 3485 45695 3519
rect 5365 3417 5399 3451
rect 6101 3417 6135 3451
rect 7757 3417 7791 3451
rect 20269 3417 20303 3451
rect 21925 3417 21959 3451
rect 36093 3417 36127 3451
rect 37749 3417 37783 3451
rect 40049 3417 40083 3451
rect 48145 3417 48179 3451
rect 2237 3349 2271 3383
rect 8309 3349 8343 3383
rect 17877 3349 17911 3383
rect 18521 3349 18555 3383
rect 22477 3349 22511 3383
rect 23765 3349 23799 3383
rect 45753 3349 45787 3383
rect 18889 3145 18923 3179
rect 36185 3145 36219 3179
rect 39589 3145 39623 3179
rect 41521 3145 41555 3179
rect 1961 3077 1995 3111
rect 8125 3077 8159 3111
rect 13737 3077 13771 3111
rect 19625 3077 19659 3111
rect 21005 3077 21039 3111
rect 22201 3077 22235 3111
rect 24777 3077 24811 3111
rect 33241 3077 33275 3111
rect 42625 3077 42659 3111
rect 44281 3077 44315 3111
rect 45385 3077 45419 3111
rect 1777 3009 1811 3043
rect 6561 3009 6595 3043
rect 7941 3009 7975 3043
rect 10977 3009 11011 3043
rect 13553 3009 13587 3043
rect 17877 3009 17911 3043
rect 18797 3009 18831 3043
rect 19533 3009 19567 3043
rect 20361 3009 20395 3043
rect 20913 3009 20947 3043
rect 22017 3009 22051 3043
rect 24593 3009 24627 3043
rect 33057 3009 33091 3043
rect 36369 3009 36403 3043
rect 39129 3009 39163 3043
rect 40325 3009 40359 3043
rect 41429 3009 41463 3043
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 47777 3009 47811 3043
rect 2237 2941 2271 2975
rect 8401 2941 8435 2975
rect 14197 2941 14231 2975
rect 17785 2941 17819 2975
rect 18245 2941 18279 2975
rect 22569 2941 22603 2975
rect 25145 2941 25179 2975
rect 33517 2941 33551 2975
rect 38945 2941 38979 2975
rect 40049 2941 40083 2975
rect 47041 2941 47075 2975
rect 47961 2873 47995 2907
rect 7297 2805 7331 2839
rect 18613 2601 18647 2635
rect 19349 2601 19383 2635
rect 23029 2601 23063 2635
rect 25513 2601 25547 2635
rect 26341 2601 26375 2635
rect 45477 2601 45511 2635
rect 20545 2533 20579 2567
rect 27629 2533 27663 2567
rect 38393 2533 38427 2567
rect 40509 2533 40543 2567
rect 47961 2533 47995 2567
rect 5273 2465 5307 2499
rect 6561 2465 6595 2499
rect 7389 2465 7423 2499
rect 15577 2465 15611 2499
rect 25053 2465 25087 2499
rect 28733 2465 28767 2499
rect 30021 2465 30055 2499
rect 46213 2465 46247 2499
rect 2697 2397 2731 2431
rect 4997 2397 5031 2431
rect 8953 2397 8987 2431
rect 15301 2397 15335 2431
rect 18521 2397 18555 2431
rect 19257 2397 19291 2431
rect 21281 2397 21315 2431
rect 22017 2397 22051 2431
rect 23121 2397 23155 2431
rect 25697 2397 25731 2431
rect 29745 2397 29779 2431
rect 35541 2397 35575 2431
rect 35817 2397 35851 2431
rect 41061 2397 41095 2431
rect 41337 2397 41371 2431
rect 43637 2397 43671 2431
rect 43913 2397 43947 2431
rect 46489 2397 46523 2431
rect 1869 2329 1903 2363
rect 6745 2329 6779 2363
rect 17141 2329 17175 2363
rect 20361 2329 20395 2363
rect 21097 2329 21131 2363
rect 24869 2329 24903 2363
rect 26249 2329 26283 2363
rect 27445 2329 27479 2363
rect 28549 2329 28583 2363
rect 38209 2329 38243 2363
rect 40325 2329 40359 2363
rect 45385 2329 45419 2363
rect 47777 2329 47811 2363
rect 2145 2261 2179 2295
rect 2881 2261 2915 2295
rect 9137 2261 9171 2295
rect 17233 2261 17267 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 19334 47132 19340 47184
rect 19392 47172 19398 47184
rect 19429 47175 19487 47181
rect 19429 47172 19441 47175
rect 19392 47144 19441 47172
rect 19392 47132 19398 47144
rect 19429 47141 19441 47144
rect 19475 47141 19487 47175
rect 19429 47135 19487 47141
rect 29362 47132 29368 47184
rect 29420 47172 29426 47184
rect 29917 47175 29975 47181
rect 29917 47172 29929 47175
rect 29420 47144 29929 47172
rect 29420 47132 29426 47144
rect 29917 47141 29929 47144
rect 29963 47141 29975 47175
rect 29917 47135 29975 47141
rect 47854 47132 47860 47184
rect 47912 47172 47918 47184
rect 47949 47175 48007 47181
rect 47949 47172 47961 47175
rect 47912 47144 47961 47172
rect 47912 47132 47918 47144
rect 47949 47141 47961 47144
rect 47995 47141 48007 47175
rect 47949 47135 48007 47141
rect 13814 47064 13820 47116
rect 13872 47104 13878 47116
rect 14093 47107 14151 47113
rect 14093 47104 14105 47107
rect 13872 47076 14105 47104
rect 13872 47064 13878 47076
rect 14093 47073 14105 47076
rect 14139 47073 14151 47107
rect 14093 47067 14151 47073
rect 16945 47107 17003 47113
rect 16945 47073 16957 47107
rect 16991 47104 17003 47107
rect 22094 47104 22100 47116
rect 16991 47076 22100 47104
rect 16991 47073 17003 47076
rect 16945 47067 17003 47073
rect 22094 47064 22100 47076
rect 22152 47064 22158 47116
rect 30742 47104 30748 47116
rect 30703 47076 30748 47104
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 43162 47104 43168 47116
rect 43123 47076 43168 47104
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 2130 47036 2136 47048
rect 2091 47008 2136 47036
rect 2130 46996 2136 47008
rect 2188 46996 2194 47048
rect 2774 46996 2780 47048
rect 2832 47036 2838 47048
rect 2961 47039 3019 47045
rect 2961 47036 2973 47039
rect 2832 47008 2973 47036
rect 2832 46996 2838 47008
rect 2961 47005 2973 47008
rect 3007 47005 3019 47039
rect 2961 46999 3019 47005
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6825 47039 6883 47045
rect 6825 47036 6837 47039
rect 5868 47008 6837 47036
rect 5868 46996 5874 47008
rect 6825 47005 6837 47008
rect 6871 47005 6883 47039
rect 6825 46999 6883 47005
rect 7098 46996 7104 47048
rect 7156 47036 7162 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7156 47008 7757 47036
rect 7156 46996 7162 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 7745 46999 7803 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9401 47039 9459 47045
rect 9401 47036 9413 47039
rect 9088 47008 9413 47036
rect 9088 46996 9094 47008
rect 9401 47005 9413 47008
rect 9447 47005 9459 47039
rect 11606 47036 11612 47048
rect 11567 47008 11612 47036
rect 9401 46999 9459 47005
rect 11606 46996 11612 47008
rect 11664 46996 11670 47048
rect 12250 46996 12256 47048
rect 12308 47036 12314 47048
rect 12345 47039 12403 47045
rect 12345 47036 12357 47039
rect 12308 47008 12357 47036
rect 12308 46996 12314 47008
rect 12345 47005 12357 47008
rect 12391 47005 12403 47039
rect 12345 46999 12403 47005
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 14366 47036 14372 47048
rect 14327 47008 14372 47036
rect 13081 46999 13139 47005
rect 14366 46996 14372 47008
rect 14424 46996 14430 47048
rect 16482 46996 16488 47048
rect 16540 47036 16546 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16540 47008 16681 47036
rect 16540 46996 16546 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 19245 46999 19303 47005
rect 19426 46996 19432 47048
rect 19484 47036 19490 47048
rect 20257 47039 20315 47045
rect 20257 47036 20269 47039
rect 19484 47008 20269 47036
rect 19484 46996 19490 47008
rect 20257 47005 20269 47008
rect 20303 47005 20315 47039
rect 20898 47036 20904 47048
rect 20859 47008 20904 47036
rect 20257 46999 20315 47005
rect 20898 46996 20904 47008
rect 20956 46996 20962 47048
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21008 47008 22017 47036
rect 2498 46968 2504 46980
rect 2459 46940 2504 46968
rect 2498 46928 2504 46940
rect 2556 46928 2562 46980
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 7834 46928 7840 46980
rect 7892 46968 7898 46980
rect 7929 46971 7987 46977
rect 7929 46968 7941 46971
rect 7892 46940 7941 46968
rect 7892 46928 7898 46940
rect 7929 46937 7941 46940
rect 7975 46937 7987 46971
rect 7929 46931 7987 46937
rect 9490 46928 9496 46980
rect 9548 46968 9554 46980
rect 9585 46971 9643 46977
rect 9585 46968 9597 46971
rect 9548 46940 9597 46968
rect 9548 46928 9554 46940
rect 9585 46937 9597 46940
rect 9631 46937 9643 46971
rect 9585 46931 9643 46937
rect 11698 46928 11704 46980
rect 11756 46968 11762 46980
rect 11793 46971 11851 46977
rect 11793 46968 11805 46971
rect 11756 46940 11805 46968
rect 11756 46928 11762 46940
rect 11793 46937 11805 46940
rect 11839 46937 11851 46971
rect 11793 46931 11851 46937
rect 12434 46928 12440 46980
rect 12492 46968 12498 46980
rect 12529 46971 12587 46977
rect 12529 46968 12541 46971
rect 12492 46940 12541 46968
rect 12492 46928 12498 46940
rect 12529 46937 12541 46940
rect 12575 46937 12587 46971
rect 12529 46931 12587 46937
rect 13449 46971 13507 46977
rect 13449 46937 13461 46971
rect 13495 46968 13507 46971
rect 15838 46968 15844 46980
rect 13495 46940 15844 46968
rect 13495 46937 13507 46940
rect 13449 46931 13507 46937
rect 15838 46928 15844 46940
rect 15896 46928 15902 46980
rect 3142 46900 3148 46912
rect 3103 46872 3148 46900
rect 3142 46860 3148 46872
rect 3200 46860 3206 46912
rect 6914 46860 6920 46912
rect 6972 46900 6978 46912
rect 6972 46872 7017 46900
rect 6972 46860 6978 46872
rect 15286 46860 15292 46912
rect 15344 46900 15350 46912
rect 16482 46900 16488 46912
rect 15344 46872 16488 46900
rect 15344 46860 15350 46872
rect 16482 46860 16488 46872
rect 16540 46860 16546 46912
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 21008 46900 21036 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 24578 46996 24584 47048
rect 24636 47036 24642 47048
rect 24765 47039 24823 47045
rect 24765 47036 24777 47039
rect 24636 47008 24777 47036
rect 24636 46996 24642 47008
rect 24765 47005 24777 47008
rect 24811 47005 24823 47039
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 24765 46999 24823 47005
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28629 47039 28687 47045
rect 28629 47036 28641 47039
rect 28408 47008 28641 47036
rect 28408 46996 28414 47008
rect 28629 47005 28641 47008
rect 28675 47005 28687 47039
rect 28629 46999 28687 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 31021 47039 31079 47045
rect 31021 47005 31033 47039
rect 31067 47036 31079 47039
rect 31110 47036 31116 47048
rect 31067 47008 31116 47036
rect 31067 47005 31079 47008
rect 31021 46999 31079 47005
rect 31110 46996 31116 47008
rect 31168 46996 31174 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38381 47039 38439 47045
rect 38381 47036 38393 47039
rect 38160 47008 38393 47036
rect 38160 46996 38166 47008
rect 38381 47005 38393 47008
rect 38427 47005 38439 47039
rect 41874 47036 41880 47048
rect 41835 47008 41880 47036
rect 38381 46999 38439 47005
rect 41874 46996 41880 47008
rect 41932 46996 41938 47048
rect 42610 47036 42616 47048
rect 42571 47008 42616 47036
rect 42610 46996 42616 47008
rect 42668 46996 42674 47048
rect 45186 47036 45192 47048
rect 45147 47008 45192 47036
rect 45186 46996 45192 47008
rect 45244 46996 45250 47048
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 21818 46900 21824 46912
rect 20036 46872 21036 46900
rect 21779 46872 21824 46900
rect 20036 46860 20042 46872
rect 21818 46860 21824 46872
rect 21876 46860 21882 46912
rect 28258 46860 28264 46912
rect 28316 46900 28322 46912
rect 28445 46903 28503 46909
rect 28445 46900 28457 46903
rect 28316 46872 28457 46900
rect 28316 46860 28322 46872
rect 28445 46869 28457 46872
rect 28491 46869 28503 46903
rect 28445 46863 28503 46869
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 42797 46971 42855 46977
rect 42797 46937 42809 46971
rect 42843 46968 42855 46971
rect 42886 46968 42892 46980
rect 42843 46940 42892 46968
rect 42843 46937 42855 46940
rect 42797 46931 42855 46937
rect 42886 46928 42892 46940
rect 42944 46928 42950 46980
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 39356 46872 40356 46900
rect 39356 46860 39362 46872
rect 46382 46860 46388 46912
rect 46440 46900 46446 46912
rect 47118 46900 47124 46912
rect 46440 46872 47124 46900
rect 46440 46860 46446 46872
rect 47118 46860 47124 46872
rect 47176 46860 47182 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 6886 46668 26234 46696
rect 1854 46628 1860 46640
rect 1815 46600 1860 46628
rect 1854 46588 1860 46600
rect 1912 46588 1918 46640
rect 3142 46588 3148 46640
rect 3200 46628 3206 46640
rect 6886 46628 6914 46668
rect 3200 46600 6914 46628
rect 26206 46628 26234 46668
rect 28445 46631 28503 46637
rect 28445 46628 28457 46631
rect 26206 46600 28457 46628
rect 3200 46588 3206 46600
rect 28445 46597 28457 46600
rect 28491 46597 28503 46631
rect 28445 46591 28503 46597
rect 30101 46631 30159 46637
rect 30101 46597 30113 46631
rect 30147 46628 30159 46631
rect 30147 46600 35894 46628
rect 30147 46597 30159 46600
rect 30101 46591 30159 46597
rect 19426 46560 19432 46572
rect 19387 46532 19432 46560
rect 19426 46520 19432 46532
rect 19484 46520 19490 46572
rect 24578 46560 24584 46572
rect 24539 46532 24584 46560
rect 24578 46520 24584 46532
rect 24636 46520 24642 46572
rect 28258 46560 28264 46572
rect 28219 46532 28264 46560
rect 28258 46520 28264 46532
rect 28316 46520 28322 46572
rect 3421 46495 3479 46501
rect 3421 46461 3433 46495
rect 3467 46461 3479 46495
rect 3421 46455 3479 46461
rect 3605 46495 3663 46501
rect 3605 46461 3617 46495
rect 3651 46492 3663 46495
rect 3878 46492 3884 46504
rect 3651 46464 3884 46492
rect 3651 46461 3663 46464
rect 3605 46455 3663 46461
rect 3436 46424 3464 46455
rect 3878 46452 3884 46464
rect 3936 46452 3942 46504
rect 3970 46452 3976 46504
rect 4028 46492 4034 46504
rect 4157 46495 4215 46501
rect 4157 46492 4169 46495
rect 4028 46464 4169 46492
rect 4028 46452 4034 46464
rect 4157 46461 4169 46464
rect 4203 46461 4215 46495
rect 4157 46455 4215 46461
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46461 11759 46495
rect 11701 46455 11759 46461
rect 11977 46495 12035 46501
rect 11977 46461 11989 46495
rect 12023 46461 12035 46495
rect 13814 46492 13820 46504
rect 13775 46464 13820 46492
rect 11977 46455 12035 46461
rect 4614 46424 4620 46436
rect 3436 46396 4620 46424
rect 4614 46384 4620 46396
rect 4672 46384 4678 46436
rect 11238 46384 11244 46436
rect 11296 46424 11302 46436
rect 11716 46424 11744 46455
rect 11296 46396 11744 46424
rect 11296 46384 11302 46396
rect 2133 46359 2191 46365
rect 2133 46325 2145 46359
rect 2179 46356 2191 46359
rect 2590 46356 2596 46368
rect 2179 46328 2596 46356
rect 2179 46325 2191 46328
rect 2133 46319 2191 46325
rect 2590 46316 2596 46328
rect 2648 46316 2654 46368
rect 2866 46356 2872 46368
rect 2827 46328 2872 46356
rect 2866 46316 2872 46328
rect 2924 46316 2930 46368
rect 10962 46316 10968 46368
rect 11020 46356 11026 46368
rect 11992 46356 12020 46455
rect 13814 46452 13820 46464
rect 13872 46452 13878 46504
rect 13998 46492 14004 46504
rect 13959 46464 14004 46492
rect 13998 46452 14004 46464
rect 14056 46452 14062 46504
rect 14182 46452 14188 46504
rect 14240 46492 14246 46504
rect 14277 46495 14335 46501
rect 14277 46492 14289 46495
rect 14240 46464 14289 46492
rect 14240 46452 14246 46464
rect 14277 46461 14289 46464
rect 14323 46461 14335 46495
rect 14277 46455 14335 46461
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46492 19671 46495
rect 20162 46492 20168 46504
rect 19659 46464 20168 46492
rect 19659 46461 19671 46464
rect 19613 46455 19671 46461
rect 20162 46452 20168 46464
rect 20220 46452 20226 46504
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 32585 46455 32643 46461
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 32272 46396 32628 46424
rect 35866 46424 35894 46600
rect 38378 46588 38384 46640
rect 38436 46628 38442 46640
rect 45922 46628 45928 46640
rect 38436 46600 45928 46628
rect 38436 46588 38442 46600
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 41708 46569 41736 46600
rect 45922 46588 45928 46600
rect 45980 46588 45986 46640
rect 41693 46563 41751 46569
rect 41693 46529 41705 46563
rect 41739 46529 41751 46563
rect 41693 46523 41751 46529
rect 41874 46520 41880 46572
rect 41932 46560 41938 46572
rect 42429 46563 42487 46569
rect 42429 46560 42441 46563
rect 41932 46532 42441 46560
rect 41932 46520 41938 46532
rect 42429 46529 42441 46532
rect 42475 46529 42487 46563
rect 42429 46523 42487 46529
rect 47857 46563 47915 46569
rect 47857 46529 47869 46563
rect 47903 46560 47915 46563
rect 47946 46560 47952 46572
rect 47903 46532 47952 46560
rect 47903 46529 47915 46532
rect 47857 46523 47915 46529
rect 47946 46520 47952 46532
rect 48004 46520 48010 46572
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41785 46495 41843 46501
rect 41785 46461 41797 46495
rect 41831 46492 41843 46495
rect 42613 46495 42671 46501
rect 42613 46492 42625 46495
rect 41831 46464 42625 46492
rect 41831 46461 41843 46464
rect 41785 46455 41843 46461
rect 42613 46461 42625 46464
rect 42659 46461 42671 46495
rect 42613 46455 42671 46461
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46290 46492 46296 46504
rect 45419 46464 46296 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 35866 46396 41460 46424
rect 32272 46384 32278 46396
rect 11020 46328 12020 46356
rect 11020 46316 11026 46328
rect 33778 46316 33784 46368
rect 33836 46356 33842 46368
rect 39942 46356 39948 46368
rect 33836 46328 39948 46356
rect 33836 46316 33842 46328
rect 39942 46316 39948 46328
rect 40000 46316 40006 46368
rect 41233 46359 41291 46365
rect 41233 46325 41245 46359
rect 41279 46356 41291 46359
rect 41322 46356 41328 46368
rect 41279 46328 41328 46356
rect 41279 46325 41291 46328
rect 41233 46319 41291 46325
rect 41322 46316 41328 46328
rect 41380 46316 41386 46368
rect 41432 46356 41460 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 42576 46396 42932 46424
rect 45204 46424 45232 46455
rect 46290 46452 46296 46464
rect 46348 46452 46354 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 47762 46424 47768 46436
rect 45204 46396 47768 46424
rect 42576 46384 42582 46396
rect 47762 46384 47768 46396
rect 47820 46384 47826 46436
rect 43530 46356 43536 46368
rect 41432 46328 43536 46356
rect 43530 46316 43536 46328
rect 43588 46316 43594 46368
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3878 46152 3884 46164
rect 3839 46124 3884 46152
rect 3878 46112 3884 46124
rect 3936 46112 3942 46164
rect 4614 46152 4620 46164
rect 4575 46124 4620 46152
rect 4614 46112 4620 46124
rect 4672 46112 4678 46164
rect 11238 46152 11244 46164
rect 11199 46124 11244 46152
rect 11238 46112 11244 46124
rect 11296 46112 11302 46164
rect 13814 46112 13820 46164
rect 13872 46152 13878 46164
rect 14277 46155 14335 46161
rect 14277 46152 14289 46155
rect 13872 46124 14289 46152
rect 13872 46112 13878 46124
rect 14277 46121 14289 46124
rect 14323 46121 14335 46155
rect 20162 46152 20168 46164
rect 20123 46124 20168 46152
rect 14277 46115 14335 46121
rect 20162 46112 20168 46124
rect 20220 46112 20226 46164
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 20717 46019 20775 46025
rect 20717 45985 20729 46019
rect 20763 46016 20775 46019
rect 20898 46016 20904 46028
rect 20763 45988 20904 46016
rect 20763 45985 20775 45988
rect 20717 45979 20775 45985
rect 20898 45976 20904 45988
rect 20956 45976 20962 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25498 46016 25504 46028
rect 25271 45988 25504 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 41322 46016 41328 46028
rect 41283 45988 41328 46016
rect 41322 45976 41328 45988
rect 41380 45976 41386 46028
rect 41966 46016 41972 46028
rect 41927 45988 41972 46016
rect 41966 45976 41972 45988
rect 42024 45976 42030 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 2869 45951 2927 45957
rect 2869 45917 2881 45951
rect 2915 45948 2927 45951
rect 3789 45951 3847 45957
rect 3789 45948 3801 45951
rect 2915 45920 3801 45948
rect 2915 45917 2927 45920
rect 2869 45911 2927 45917
rect 3789 45917 3801 45920
rect 3835 45917 3847 45951
rect 3789 45911 3847 45917
rect 11149 45951 11207 45957
rect 11149 45917 11161 45951
rect 11195 45948 11207 45951
rect 20070 45948 20076 45960
rect 11195 45920 16574 45948
rect 20031 45920 20076 45948
rect 11195 45917 11207 45920
rect 11149 45911 11207 45917
rect 3804 45880 3832 45911
rect 16546 45880 16574 45920
rect 20070 45908 20076 45920
rect 20128 45908 20134 45960
rect 24118 45908 24124 45960
rect 24176 45948 24182 45960
rect 24581 45951 24639 45957
rect 24581 45948 24593 45951
rect 24176 45920 24593 45948
rect 24176 45908 24182 45920
rect 24581 45917 24593 45920
rect 24627 45917 24639 45951
rect 38194 45948 38200 45960
rect 38107 45920 38200 45948
rect 24581 45911 24639 45917
rect 38194 45908 38200 45920
rect 38252 45948 38258 45960
rect 38378 45948 38384 45960
rect 38252 45920 38384 45948
rect 38252 45908 38258 45920
rect 38378 45908 38384 45920
rect 38436 45908 38442 45960
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43901 45951 43959 45957
rect 43901 45948 43913 45951
rect 43864 45920 43913 45948
rect 43864 45908 43870 45920
rect 43901 45917 43913 45920
rect 43947 45917 43959 45951
rect 43901 45911 43959 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45948 45707 45951
rect 45738 45948 45744 45960
rect 45695 45920 45744 45948
rect 45695 45917 45707 45920
rect 45649 45911 45707 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 45830 45908 45836 45960
rect 45888 45948 45894 45960
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45888 45920 46305 45948
rect 45888 45908 45894 45920
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 20714 45880 20720 45892
rect 3804 45852 6914 45880
rect 16546 45852 20720 45880
rect 2958 45812 2964 45824
rect 2919 45784 2964 45812
rect 2958 45772 2964 45784
rect 3016 45772 3022 45824
rect 6886 45812 6914 45852
rect 20714 45840 20720 45852
rect 20772 45840 20778 45892
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 41506 45880 41512 45892
rect 41467 45852 41512 45880
rect 41506 45840 41512 45852
rect 41564 45840 41570 45892
rect 46474 45880 46480 45892
rect 46435 45852 46480 45880
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 25314 45812 25320 45824
rect 6886 45784 25320 45812
rect 25314 45772 25320 45784
rect 25372 45772 25378 45824
rect 44082 45812 44088 45824
rect 44043 45784 44088 45812
rect 44082 45772 44088 45784
rect 44140 45772 44146 45824
rect 45554 45772 45560 45824
rect 45612 45812 45618 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 45612 45784 45753 45812
rect 45612 45772 45618 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45741 45775 45799 45781
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 13817 45611 13875 45617
rect 13817 45577 13829 45611
rect 13863 45608 13875 45611
rect 13998 45608 14004 45620
rect 13863 45580 14004 45608
rect 13863 45577 13875 45580
rect 13817 45571 13875 45577
rect 13998 45568 14004 45580
rect 14056 45568 14062 45620
rect 20898 45608 20904 45620
rect 20859 45580 20904 45608
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 25406 45608 25412 45620
rect 25367 45580 25412 45608
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 32217 45611 32275 45617
rect 32217 45577 32229 45611
rect 32263 45608 32275 45611
rect 32306 45608 32312 45620
rect 32263 45580 32312 45608
rect 32263 45577 32275 45580
rect 32217 45571 32275 45577
rect 32306 45568 32312 45580
rect 32364 45568 32370 45620
rect 41506 45608 41512 45620
rect 41467 45580 41512 45608
rect 41506 45568 41512 45580
rect 41564 45568 41570 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45646 45608 45652 45620
rect 45152 45580 45652 45608
rect 45152 45568 45158 45580
rect 45646 45568 45652 45580
rect 45704 45568 45710 45620
rect 2225 45543 2283 45549
rect 2225 45509 2237 45543
rect 2271 45540 2283 45543
rect 2958 45540 2964 45552
rect 2271 45512 2964 45540
rect 2271 45509 2283 45512
rect 2225 45503 2283 45509
rect 2958 45500 2964 45512
rect 3016 45500 3022 45552
rect 20714 45500 20720 45552
rect 20772 45540 20778 45552
rect 24118 45540 24124 45552
rect 20772 45512 24124 45540
rect 20772 45500 20778 45512
rect 13722 45472 13728 45484
rect 13683 45444 13728 45472
rect 13722 45432 13728 45444
rect 13780 45432 13786 45484
rect 20824 45481 20852 45512
rect 24118 45500 24124 45512
rect 24176 45500 24182 45552
rect 42886 45540 42892 45552
rect 42847 45512 42892 45540
rect 42886 45500 42892 45512
rect 42944 45500 42950 45552
rect 43901 45543 43959 45549
rect 43901 45509 43913 45543
rect 43947 45540 43959 45543
rect 44174 45540 44180 45552
rect 43947 45512 44180 45540
rect 43947 45509 43959 45512
rect 43901 45503 43959 45509
rect 44174 45500 44180 45512
rect 44232 45500 44238 45552
rect 45370 45500 45376 45552
rect 45428 45540 45434 45552
rect 46937 45543 46995 45549
rect 46937 45540 46949 45543
rect 45428 45512 46949 45540
rect 45428 45500 45434 45512
rect 46937 45509 46949 45512
rect 46983 45509 46995 45543
rect 46937 45503 46995 45509
rect 47118 45500 47124 45552
rect 47176 45540 47182 45552
rect 47949 45543 48007 45549
rect 47949 45540 47961 45543
rect 47176 45512 47961 45540
rect 47176 45500 47182 45512
rect 47949 45509 47961 45512
rect 47995 45509 48007 45543
rect 47949 45503 48007 45509
rect 20809 45475 20867 45481
rect 20809 45441 20821 45475
rect 20855 45472 20867 45475
rect 25314 45472 25320 45484
rect 20855 45444 20889 45472
rect 25275 45444 25320 45472
rect 20855 45441 20867 45444
rect 20809 45435 20867 45441
rect 25314 45432 25320 45444
rect 25372 45432 25378 45484
rect 32122 45472 32128 45484
rect 32083 45444 32128 45472
rect 32122 45432 32128 45444
rect 32180 45432 32186 45484
rect 41417 45475 41475 45481
rect 41417 45441 41429 45475
rect 41463 45472 41475 45475
rect 42794 45472 42800 45484
rect 41463 45444 42800 45472
rect 41463 45441 41475 45444
rect 41417 45435 41475 45441
rect 42794 45432 42800 45444
rect 42852 45432 42858 45484
rect 46658 45432 46664 45484
rect 46716 45472 46722 45484
rect 46845 45475 46903 45481
rect 46845 45472 46857 45475
rect 46716 45444 46857 45472
rect 46716 45432 46722 45444
rect 46845 45441 46857 45444
rect 46891 45441 46903 45475
rect 46845 45435 46903 45441
rect 2041 45407 2099 45413
rect 2041 45373 2053 45407
rect 2087 45404 2099 45407
rect 2866 45404 2872 45416
rect 2087 45376 2872 45404
rect 2087 45373 2099 45376
rect 2041 45367 2099 45373
rect 2866 45364 2872 45376
rect 2924 45364 2930 45416
rect 3050 45404 3056 45416
rect 3011 45376 3056 45404
rect 3050 45364 3056 45376
rect 3108 45364 3114 45416
rect 20070 45364 20076 45416
rect 20128 45404 20134 45416
rect 20128 45376 40724 45404
rect 20128 45364 20134 45376
rect 13722 45296 13728 45348
rect 13780 45336 13786 45348
rect 37182 45336 37188 45348
rect 13780 45308 37188 45336
rect 13780 45296 13786 45308
rect 37182 45296 37188 45308
rect 37240 45296 37246 45348
rect 40696 45336 40724 45376
rect 44450 45364 44456 45416
rect 44508 45404 44514 45416
rect 44545 45407 44603 45413
rect 44545 45404 44557 45407
rect 44508 45376 44557 45404
rect 44508 45364 44514 45376
rect 44545 45373 44557 45376
rect 44591 45373 44603 45407
rect 44545 45367 44603 45373
rect 44729 45407 44787 45413
rect 44729 45373 44741 45407
rect 44775 45404 44787 45407
rect 45094 45404 45100 45416
rect 44775 45376 45100 45404
rect 44775 45373 44787 45376
rect 44729 45367 44787 45373
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45646 45404 45652 45416
rect 45607 45376 45652 45404
rect 45646 45364 45652 45376
rect 45704 45364 45710 45416
rect 46658 45336 46664 45348
rect 40696 45308 46664 45336
rect 46658 45296 46664 45308
rect 46716 45296 46722 45348
rect 43990 45268 43996 45280
rect 43951 45240 43996 45268
rect 43990 45228 43996 45240
rect 44048 45228 44054 45280
rect 47210 45228 47216 45280
rect 47268 45268 47274 45280
rect 48041 45271 48099 45277
rect 48041 45268 48053 45271
rect 47268 45240 48053 45268
rect 47268 45228 47274 45240
rect 48041 45237 48053 45240
rect 48087 45237 48099 45271
rect 48041 45231 48099 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 42610 45024 42616 45076
rect 42668 45064 42674 45076
rect 42889 45067 42947 45073
rect 42889 45064 42901 45067
rect 42668 45036 42901 45064
rect 42668 45024 42674 45036
rect 42889 45033 42901 45036
rect 42935 45033 42947 45067
rect 44450 45064 44456 45076
rect 44411 45036 44456 45064
rect 42889 45027 42947 45033
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 46474 45064 46480 45076
rect 45787 45036 46480 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 46474 45024 46480 45036
rect 46532 45024 46538 45076
rect 42794 44956 42800 45008
rect 42852 44996 42858 45008
rect 47394 44996 47400 45008
rect 42852 44968 47400 44996
rect 42852 44956 42858 44968
rect 47394 44956 47400 44968
rect 47452 44956 47458 45008
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 44910 44820 44916 44872
rect 44968 44860 44974 44872
rect 45005 44863 45063 44869
rect 45005 44860 45017 44863
rect 44968 44832 45017 44860
rect 44968 44820 44974 44832
rect 45005 44829 45017 44832
rect 45051 44829 45063 44863
rect 45646 44860 45652 44872
rect 45607 44832 45652 44860
rect 45005 44823 45063 44829
rect 45646 44820 45652 44832
rect 45704 44820 45710 44872
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 46934 44792 46940 44804
rect 46523 44764 46940 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 46934 44752 46940 44764
rect 46992 44752 46998 44804
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 46290 44520 46296 44532
rect 46251 44492 46296 44520
rect 46290 44480 46296 44492
rect 46348 44480 46354 44532
rect 46934 44520 46940 44532
rect 46895 44492 46940 44520
rect 46934 44480 46940 44492
rect 46992 44480 46998 44532
rect 45646 44412 45652 44464
rect 45704 44452 45710 44464
rect 45704 44424 46244 44452
rect 45704 44412 45710 44424
rect 45097 44387 45155 44393
rect 45097 44353 45109 44387
rect 45143 44384 45155 44387
rect 45186 44384 45192 44396
rect 45143 44356 45192 44384
rect 45143 44353 45155 44356
rect 45097 44347 45155 44353
rect 45186 44344 45192 44356
rect 45244 44344 45250 44396
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46216 44393 46244 44424
rect 46201 44387 46259 44393
rect 46201 44353 46213 44387
rect 46247 44353 46259 44387
rect 46201 44347 46259 44353
rect 46845 44387 46903 44393
rect 46845 44353 46857 44387
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 37182 44276 37188 44328
rect 37240 44316 37246 44328
rect 46860 44316 46888 44347
rect 37240 44288 46888 44316
rect 37240 44276 37246 44288
rect 25314 44140 25320 44192
rect 25372 44180 25378 44192
rect 25866 44180 25872 44192
rect 25372 44152 25872 44180
rect 25372 44140 25378 44152
rect 25866 44140 25872 44152
rect 25924 44140 25930 44192
rect 47670 44180 47676 44192
rect 47631 44152 47676 44180
rect 47670 44140 47676 44152
rect 47728 44140 47734 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 47670 43840 47676 43852
rect 46523 43812 47676 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 47670 43800 47676 43812
rect 47728 43800 47734 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1854 43296 1860 43308
rect 1815 43268 1860 43296
rect 1854 43256 1860 43268
rect 1912 43256 1918 43308
rect 25498 43256 25504 43308
rect 25556 43296 25562 43308
rect 25869 43299 25927 43305
rect 25869 43296 25881 43299
rect 25556 43268 25881 43296
rect 25556 43256 25562 43268
rect 25869 43265 25881 43268
rect 25915 43296 25927 43299
rect 32122 43296 32128 43308
rect 25915 43268 32128 43296
rect 25915 43265 25927 43268
rect 25869 43259 25927 43265
rect 32122 43256 32128 43268
rect 32180 43256 32186 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47762 43296 47768 43308
rect 47723 43268 47768 43296
rect 47762 43256 47768 43268
rect 47820 43256 47826 43308
rect 1946 43092 1952 43104
rect 1907 43064 1952 43092
rect 1946 43052 1952 43064
rect 2004 43052 2010 43104
rect 25958 43092 25964 43104
rect 25919 43064 25964 43092
rect 25958 43052 25964 43064
rect 26016 43052 26022 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 25958 42752 25964 42764
rect 25919 42724 25964 42752
rect 25958 42712 25964 42724
rect 26016 42712 26022 42764
rect 27617 42755 27675 42761
rect 27617 42721 27629 42755
rect 27663 42752 27675 42755
rect 33778 42752 33784 42764
rect 27663 42724 33784 42752
rect 27663 42721 27675 42724
rect 27617 42715 27675 42721
rect 33778 42712 33784 42724
rect 33836 42712 33842 42764
rect 25222 42644 25228 42696
rect 25280 42684 25286 42696
rect 25777 42687 25835 42693
rect 25777 42684 25789 42687
rect 25280 42656 25789 42684
rect 25280 42644 25286 42656
rect 25777 42653 25789 42656
rect 25823 42653 25835 42687
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 25777 42647 25835 42653
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 25222 42344 25228 42356
rect 25183 42316 25228 42344
rect 25222 42304 25228 42316
rect 25280 42304 25286 42356
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 25133 42211 25191 42217
rect 25133 42177 25145 42211
rect 25179 42208 25191 42211
rect 25314 42208 25320 42220
rect 25179 42180 25320 42208
rect 25179 42177 25191 42180
rect 25133 42171 25191 42177
rect 25314 42168 25320 42180
rect 25372 42168 25378 42220
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47029 42171 47087 42177
rect 47394 42168 47400 42220
rect 47452 42208 47458 42220
rect 47581 42211 47639 42217
rect 47581 42208 47593 42211
rect 47452 42180 47593 42208
rect 47452 42168 47458 42180
rect 47581 42177 47593 42180
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 1636 41228 2237 41256
rect 1636 41216 1642 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 2225 41219 2283 41225
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46845 41259 46903 41265
rect 46845 41256 46857 41259
rect 46532 41228 46857 41256
rect 46532 41216 46538 41228
rect 46845 41225 46857 41228
rect 46891 41225 46903 41259
rect 46845 41219 46903 41225
rect 2130 41120 2136 41132
rect 2091 41092 2136 41120
rect 2130 41080 2136 41092
rect 2188 41080 2194 41132
rect 45830 41080 45836 41132
rect 45888 41120 45894 41132
rect 46753 41123 46811 41129
rect 46753 41120 46765 41123
rect 45888 41092 46765 41120
rect 45888 41080 45894 41092
rect 46753 41089 46765 41092
rect 46799 41089 46811 41123
rect 47946 41120 47952 41132
rect 47907 41092 47952 41120
rect 46753 41083 46811 41089
rect 47946 41080 47952 41092
rect 48004 41080 48010 41132
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 45526 40956 48145 40984
rect 43714 40876 43720 40928
rect 43772 40916 43778 40928
rect 45526 40916 45554 40956
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 43772 40888 45554 40916
rect 43772 40876 43778 40888
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 47670 40712 47676 40724
rect 47631 40684 47676 40712
rect 47670 40672 47676 40684
rect 47728 40672 47734 40724
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2041 40443 2099 40449
rect 2041 40409 2053 40443
rect 2087 40440 2099 40443
rect 2406 40440 2412 40452
rect 2087 40412 2412 40440
rect 2087 40409 2099 40412
rect 2041 40403 2099 40409
rect 2406 40400 2412 40412
rect 2464 40400 2470 40452
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 46348 39800 47777 39828
rect 46348 39788 46354 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 46934 39352 46940 39364
rect 46523 39324 46940 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 46934 39312 46940 39324
rect 46992 39312 46998 39364
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 46934 39080 46940 39092
rect 46895 39052 46940 39080
rect 46934 39040 46940 39052
rect 46992 39040 46998 39092
rect 46106 38904 46112 38956
rect 46164 38944 46170 38956
rect 46845 38947 46903 38953
rect 46845 38944 46857 38947
rect 46164 38916 46857 38944
rect 46164 38904 46170 38916
rect 46845 38913 46857 38916
rect 46891 38913 46903 38947
rect 47762 38944 47768 38956
rect 47723 38916 47768 38944
rect 46845 38907 46903 38913
rect 47762 38904 47768 38916
rect 47820 38904 47826 38956
rect 47762 38700 47768 38752
rect 47820 38740 47826 38752
rect 47857 38743 47915 38749
rect 47857 38740 47869 38743
rect 47820 38712 47869 38740
rect 47820 38700 47826 38712
rect 47857 38709 47869 38712
rect 47903 38709 47915 38743
rect 47857 38703 47915 38709
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 47670 38264 47676 38276
rect 46523 38236 47676 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 47670 38224 47676 38236
rect 47728 38224 47734 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 47670 37992 47676 38004
rect 47631 37964 47676 37992
rect 47670 37952 47676 37964
rect 47728 37952 47734 38004
rect 25130 37884 25136 37936
rect 25188 37884 25194 37936
rect 19426 37816 19432 37868
rect 19484 37856 19490 37868
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19484 37828 19625 37856
rect 19484 37816 19490 37828
rect 19613 37825 19625 37828
rect 19659 37825 19671 37859
rect 19613 37819 19671 37825
rect 32122 37816 32128 37868
rect 32180 37856 32186 37868
rect 47581 37859 47639 37865
rect 47581 37856 47593 37859
rect 32180 37828 47593 37856
rect 32180 37816 32186 37828
rect 47581 37825 47593 37828
rect 47627 37825 47639 37859
rect 47581 37819 47639 37825
rect 24397 37791 24455 37797
rect 24397 37757 24409 37791
rect 24443 37757 24455 37791
rect 24397 37751 24455 37757
rect 24673 37791 24731 37797
rect 24673 37757 24685 37791
rect 24719 37788 24731 37791
rect 25038 37788 25044 37800
rect 24719 37760 25044 37788
rect 24719 37757 24731 37760
rect 24673 37751 24731 37757
rect 19429 37655 19487 37661
rect 19429 37621 19441 37655
rect 19475 37652 19487 37655
rect 19518 37652 19524 37664
rect 19475 37624 19524 37652
rect 19475 37621 19487 37624
rect 19429 37615 19487 37621
rect 19518 37612 19524 37624
rect 19576 37612 19582 37664
rect 24412 37652 24440 37751
rect 25038 37748 25044 37760
rect 25096 37748 25102 37800
rect 26234 37720 26240 37732
rect 26068 37692 26240 37720
rect 26068 37652 26096 37692
rect 26234 37680 26240 37692
rect 26292 37680 26298 37732
rect 24412 37624 26096 37652
rect 26142 37612 26148 37664
rect 26200 37652 26206 37664
rect 26200 37624 26245 37652
rect 26200 37612 26206 37624
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 25038 37448 25044 37460
rect 24999 37420 25044 37448
rect 25038 37408 25044 37420
rect 25096 37408 25102 37460
rect 46290 37408 46296 37460
rect 46348 37448 46354 37460
rect 47673 37451 47731 37457
rect 47673 37448 47685 37451
rect 46348 37420 47685 37448
rect 46348 37408 46354 37420
rect 47673 37417 47685 37420
rect 47719 37417 47731 37451
rect 47673 37411 47731 37417
rect 19518 37312 19524 37324
rect 19479 37284 19524 37312
rect 19518 37272 19524 37284
rect 19576 37272 19582 37324
rect 26329 37315 26387 37321
rect 26329 37281 26341 37315
rect 26375 37312 26387 37315
rect 27246 37312 27252 37324
rect 26375 37284 27016 37312
rect 27207 37284 27252 37312
rect 26375 37281 26387 37284
rect 26329 37275 26387 37281
rect 19242 37244 19248 37256
rect 19203 37216 19248 37244
rect 19242 37204 19248 37216
rect 19300 37204 19306 37256
rect 22738 37244 22744 37256
rect 22699 37216 22744 37244
rect 22738 37204 22744 37216
rect 22796 37204 22802 37256
rect 26988 37253 27016 37284
rect 27246 37272 27252 37284
rect 27304 37272 27310 37324
rect 45554 37312 45560 37324
rect 27540 37284 45560 37312
rect 23569 37247 23627 37253
rect 23569 37244 23581 37247
rect 22940 37216 23581 37244
rect 21174 37176 21180 37188
rect 20746 37148 21180 37176
rect 21174 37136 21180 37148
rect 21232 37136 21238 37188
rect 20254 37068 20260 37120
rect 20312 37108 20318 37120
rect 20993 37111 21051 37117
rect 20993 37108 21005 37111
rect 20312 37080 21005 37108
rect 20312 37068 20318 37080
rect 20993 37077 21005 37080
rect 21039 37077 21051 37111
rect 20993 37071 21051 37077
rect 22462 37068 22468 37120
rect 22520 37108 22526 37120
rect 22940 37117 22968 37216
rect 23569 37213 23581 37216
rect 23615 37213 23627 37247
rect 23569 37207 23627 37213
rect 25225 37247 25283 37253
rect 25225 37213 25237 37247
rect 25271 37244 25283 37247
rect 26973 37247 27031 37253
rect 25271 37216 26648 37244
rect 25271 37213 25283 37216
rect 25225 37207 25283 37213
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22520 37080 22937 37108
rect 22520 37068 22526 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 23658 37108 23664 37120
rect 23619 37080 23664 37108
rect 22925 37071 22983 37077
rect 23658 37068 23664 37080
rect 23716 37068 23722 37120
rect 26620 37117 26648 37216
rect 26973 37213 26985 37247
rect 27019 37244 27031 37247
rect 27540 37244 27568 37284
rect 45554 37272 45560 37284
rect 45612 37272 45618 37324
rect 27019 37216 27568 37244
rect 27019 37213 27031 37216
rect 26973 37207 27031 37213
rect 26605 37111 26663 37117
rect 26605 37077 26617 37111
rect 26651 37077 26663 37111
rect 26605 37071 26663 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27120 37080 27165 37108
rect 27120 37068 27126 37080
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 19429 36907 19487 36913
rect 19429 36873 19441 36907
rect 19475 36904 19487 36907
rect 20349 36907 20407 36913
rect 20349 36904 20361 36907
rect 19475 36876 20361 36904
rect 19475 36873 19487 36876
rect 19429 36867 19487 36873
rect 20349 36873 20361 36876
rect 20395 36873 20407 36907
rect 21174 36904 21180 36916
rect 21135 36876 21180 36904
rect 20349 36867 20407 36873
rect 21174 36864 21180 36876
rect 21232 36864 21238 36916
rect 27246 36904 27252 36916
rect 22480 36876 27252 36904
rect 20257 36839 20315 36845
rect 20257 36805 20269 36839
rect 20303 36836 20315 36839
rect 21818 36836 21824 36848
rect 20303 36808 21824 36836
rect 20303 36805 20315 36808
rect 20257 36799 20315 36805
rect 21818 36796 21824 36808
rect 21876 36796 21882 36848
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36768 19119 36771
rect 20162 36768 20168 36780
rect 19107 36740 20168 36768
rect 19107 36737 19119 36740
rect 19061 36731 19119 36737
rect 20162 36728 20168 36740
rect 20220 36728 20226 36780
rect 21082 36768 21088 36780
rect 21043 36740 21088 36768
rect 21082 36728 21088 36740
rect 21140 36728 21146 36780
rect 19153 36703 19211 36709
rect 19153 36669 19165 36703
rect 19199 36700 19211 36703
rect 20438 36700 20444 36712
rect 19199 36672 20444 36700
rect 19199 36669 19211 36672
rect 19153 36663 19211 36669
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 20533 36703 20591 36709
rect 20533 36669 20545 36703
rect 20579 36700 20591 36703
rect 22480 36700 22508 36876
rect 27246 36864 27252 36876
rect 27304 36864 27310 36916
rect 23658 36796 23664 36848
rect 23716 36796 23722 36848
rect 25222 36728 25228 36780
rect 25280 36768 25286 36780
rect 25317 36771 25375 36777
rect 25317 36768 25329 36771
rect 25280 36740 25329 36768
rect 25280 36728 25286 36740
rect 25317 36737 25329 36740
rect 25363 36768 25375 36771
rect 26142 36768 26148 36780
rect 25363 36740 26148 36768
rect 25363 36737 25375 36740
rect 25317 36731 25375 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 20579 36672 22508 36700
rect 20579 36669 20591 36672
rect 20533 36663 20591 36669
rect 22554 36660 22560 36712
rect 22612 36700 22618 36712
rect 22649 36703 22707 36709
rect 22649 36700 22661 36703
rect 22612 36672 22661 36700
rect 22612 36660 22618 36672
rect 22649 36669 22661 36672
rect 22695 36669 22707 36703
rect 22922 36700 22928 36712
rect 22883 36672 22928 36700
rect 22649 36663 22707 36669
rect 22922 36660 22928 36672
rect 22980 36660 22986 36712
rect 24854 36660 24860 36712
rect 24912 36700 24918 36712
rect 25409 36703 25467 36709
rect 25409 36700 25421 36703
rect 24912 36672 25421 36700
rect 24912 36660 24918 36672
rect 25409 36669 25421 36672
rect 25455 36669 25467 36703
rect 25409 36663 25467 36669
rect 25685 36703 25743 36709
rect 25685 36669 25697 36703
rect 25731 36700 25743 36703
rect 27062 36700 27068 36712
rect 25731 36672 27068 36700
rect 25731 36669 25743 36672
rect 25685 36663 25743 36669
rect 27062 36660 27068 36672
rect 27120 36660 27126 36712
rect 19889 36567 19947 36573
rect 19889 36533 19901 36567
rect 19935 36564 19947 36567
rect 20162 36564 20168 36576
rect 19935 36536 20168 36564
rect 19935 36533 19947 36536
rect 19889 36527 19947 36533
rect 20162 36524 20168 36536
rect 20220 36524 20226 36576
rect 24397 36567 24455 36573
rect 24397 36533 24409 36567
rect 24443 36564 24455 36567
rect 24946 36564 24952 36576
rect 24443 36536 24952 36564
rect 24443 36533 24455 36536
rect 24397 36527 24455 36533
rect 24946 36524 24952 36536
rect 25004 36524 25010 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 19426 36320 19432 36372
rect 19484 36360 19490 36372
rect 19705 36363 19763 36369
rect 19705 36360 19717 36363
rect 19484 36332 19717 36360
rect 19484 36320 19490 36332
rect 19705 36329 19717 36332
rect 19751 36329 19763 36363
rect 19705 36323 19763 36329
rect 22741 36363 22799 36369
rect 22741 36329 22753 36363
rect 22787 36360 22799 36363
rect 22922 36360 22928 36372
rect 22787 36332 22928 36360
rect 22787 36329 22799 36332
rect 22741 36323 22799 36329
rect 22922 36320 22928 36332
rect 22980 36320 22986 36372
rect 24489 36363 24547 36369
rect 24489 36329 24501 36363
rect 24535 36360 24547 36363
rect 25130 36360 25136 36372
rect 24535 36332 25136 36360
rect 24535 36329 24547 36332
rect 24489 36323 24547 36329
rect 25130 36320 25136 36332
rect 25188 36320 25194 36372
rect 12434 36252 12440 36304
rect 12492 36292 12498 36304
rect 23109 36295 23167 36301
rect 23109 36292 23121 36295
rect 12492 36264 23121 36292
rect 12492 36252 12498 36264
rect 23109 36261 23121 36264
rect 23155 36261 23167 36295
rect 23109 36255 23167 36261
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 20162 36224 20168 36236
rect 20123 36196 20168 36224
rect 20162 36184 20168 36196
rect 20220 36184 20226 36236
rect 20349 36227 20407 36233
rect 20349 36193 20361 36227
rect 20395 36224 20407 36227
rect 20395 36196 22094 36224
rect 20395 36193 20407 36196
rect 20349 36187 20407 36193
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36156 20131 36159
rect 20254 36156 20260 36168
rect 20119 36128 20260 36156
rect 20119 36125 20131 36128
rect 20073 36119 20131 36125
rect 20254 36116 20260 36128
rect 20312 36116 20318 36168
rect 22066 36156 22094 36196
rect 22462 36184 22468 36236
rect 22520 36224 22526 36236
rect 22520 36196 24440 36224
rect 22520 36184 22526 36196
rect 22830 36156 22836 36168
rect 22066 36128 22836 36156
rect 22830 36116 22836 36128
rect 22888 36116 22894 36168
rect 22925 36159 22983 36165
rect 22925 36125 22937 36159
rect 22971 36125 22983 36159
rect 23198 36156 23204 36168
rect 23159 36128 23204 36156
rect 22925 36119 22983 36125
rect 1581 36091 1639 36097
rect 1581 36057 1593 36091
rect 1627 36088 1639 36091
rect 2222 36088 2228 36100
rect 1627 36060 2228 36088
rect 1627 36057 1639 36060
rect 1581 36051 1639 36057
rect 2222 36048 2228 36060
rect 2280 36048 2286 36100
rect 22940 36020 22968 36119
rect 23198 36116 23204 36128
rect 23256 36116 23262 36168
rect 24412 36165 24440 36196
rect 24397 36159 24455 36165
rect 24397 36125 24409 36159
rect 24443 36125 24455 36159
rect 24397 36119 24455 36125
rect 24394 36020 24400 36032
rect 22940 35992 24400 36020
rect 24394 35980 24400 35992
rect 24452 35980 24458 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 19978 35708 19984 35760
rect 20036 35748 20042 35760
rect 23198 35748 23204 35760
rect 20036 35720 23204 35748
rect 20036 35708 20042 35720
rect 23198 35708 23204 35720
rect 23256 35708 23262 35760
rect 1394 35640 1400 35692
rect 1452 35680 1458 35692
rect 2041 35683 2099 35689
rect 2041 35680 2053 35683
rect 1452 35652 2053 35680
rect 1452 35640 1458 35652
rect 2041 35649 2053 35652
rect 2087 35649 2099 35683
rect 2041 35643 2099 35649
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 22462 35680 22468 35692
rect 21140 35652 22468 35680
rect 21140 35640 21146 35652
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 23753 35683 23811 35689
rect 23753 35649 23765 35683
rect 23799 35649 23811 35683
rect 26970 35680 26976 35692
rect 23753 35643 23811 35649
rect 23952 35652 26976 35680
rect 15838 35572 15844 35624
rect 15896 35612 15902 35624
rect 22738 35612 22744 35624
rect 15896 35584 22744 35612
rect 15896 35572 15902 35584
rect 22738 35572 22744 35584
rect 22796 35612 22802 35624
rect 23768 35612 23796 35643
rect 22796 35584 23796 35612
rect 22796 35572 22802 35584
rect 9490 35504 9496 35556
rect 9548 35544 9554 35556
rect 23952 35553 23980 35652
rect 26970 35640 26976 35652
rect 27028 35680 27034 35692
rect 27157 35683 27215 35689
rect 27157 35680 27169 35683
rect 27028 35652 27169 35680
rect 27028 35640 27034 35652
rect 27157 35649 27169 35652
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 29638 35640 29644 35692
rect 29696 35640 29702 35692
rect 26234 35572 26240 35624
rect 26292 35612 26298 35624
rect 27522 35612 27528 35624
rect 26292 35584 27528 35612
rect 26292 35572 26298 35584
rect 27522 35572 27528 35584
rect 27580 35612 27586 35624
rect 28261 35615 28319 35621
rect 28261 35612 28273 35615
rect 27580 35584 28273 35612
rect 27580 35572 27586 35584
rect 28261 35581 28273 35584
rect 28307 35581 28319 35615
rect 28261 35575 28319 35581
rect 28537 35615 28595 35621
rect 28537 35581 28549 35615
rect 28583 35612 28595 35615
rect 28994 35612 29000 35624
rect 28583 35584 29000 35612
rect 28583 35581 28595 35584
rect 28537 35575 28595 35581
rect 28994 35572 29000 35584
rect 29052 35572 29058 35624
rect 23937 35547 23995 35553
rect 9548 35516 23888 35544
rect 9548 35504 9554 35516
rect 7834 35436 7840 35488
rect 7892 35476 7898 35488
rect 18138 35476 18144 35488
rect 7892 35448 18144 35476
rect 7892 35436 7898 35448
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 22462 35436 22468 35488
rect 22520 35476 22526 35488
rect 22557 35479 22615 35485
rect 22557 35476 22569 35479
rect 22520 35448 22569 35476
rect 22520 35436 22526 35448
rect 22557 35445 22569 35448
rect 22603 35445 22615 35479
rect 23860 35476 23888 35516
rect 23937 35513 23949 35547
rect 23983 35513 23995 35547
rect 23937 35507 23995 35513
rect 27080 35516 28396 35544
rect 27080 35476 27108 35516
rect 23860 35448 27108 35476
rect 22557 35439 22615 35445
rect 27154 35436 27160 35488
rect 27212 35476 27218 35488
rect 27249 35479 27307 35485
rect 27249 35476 27261 35479
rect 27212 35448 27261 35476
rect 27212 35436 27218 35448
rect 27249 35445 27261 35448
rect 27295 35445 27307 35479
rect 28368 35476 28396 35516
rect 28626 35476 28632 35488
rect 28368 35448 28632 35476
rect 27249 35439 27307 35445
rect 28626 35436 28632 35448
rect 28684 35436 28690 35488
rect 30006 35476 30012 35488
rect 29967 35448 30012 35476
rect 30006 35436 30012 35448
rect 30064 35436 30070 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 19705 35275 19763 35281
rect 19705 35241 19717 35275
rect 19751 35272 19763 35275
rect 20254 35272 20260 35284
rect 19751 35244 20260 35272
rect 19751 35241 19763 35244
rect 19705 35235 19763 35241
rect 20254 35232 20260 35244
rect 20312 35232 20318 35284
rect 24946 35272 24952 35284
rect 24907 35244 24952 35272
rect 24946 35232 24952 35244
rect 25004 35232 25010 35284
rect 26970 35232 26976 35284
rect 27028 35272 27034 35284
rect 29638 35272 29644 35284
rect 27028 35244 28488 35272
rect 29599 35244 29644 35272
rect 27028 35232 27034 35244
rect 18693 35207 18751 35213
rect 18693 35173 18705 35207
rect 18739 35204 18751 35207
rect 19058 35204 19064 35216
rect 18739 35176 19064 35204
rect 18739 35173 18751 35176
rect 18693 35167 18751 35173
rect 19058 35164 19064 35176
rect 19116 35204 19122 35216
rect 19116 35176 19656 35204
rect 19116 35164 19122 35176
rect 16945 35139 17003 35145
rect 16945 35136 16957 35139
rect 14752 35108 16957 35136
rect 14752 35080 14780 35108
rect 16945 35105 16957 35108
rect 16991 35136 17003 35139
rect 19242 35136 19248 35148
rect 16991 35108 19248 35136
rect 16991 35105 17003 35108
rect 16945 35099 17003 35105
rect 19242 35096 19248 35108
rect 19300 35096 19306 35148
rect 19628 35145 19656 35176
rect 19613 35139 19671 35145
rect 19613 35105 19625 35139
rect 19659 35105 19671 35139
rect 19613 35099 19671 35105
rect 21450 35096 21456 35148
rect 21508 35136 21514 35148
rect 21545 35139 21603 35145
rect 21545 35136 21557 35139
rect 21508 35108 21557 35136
rect 21508 35096 21514 35108
rect 21545 35105 21557 35108
rect 21591 35136 21603 35139
rect 22554 35136 22560 35148
rect 21591 35108 22560 35136
rect 21591 35105 21603 35108
rect 21545 35099 21603 35105
rect 22554 35096 22560 35108
rect 22612 35136 22618 35148
rect 23014 35136 23020 35148
rect 22612 35108 23020 35136
rect 22612 35096 22618 35108
rect 23014 35096 23020 35108
rect 23072 35096 23078 35148
rect 25133 35139 25191 35145
rect 25133 35105 25145 35139
rect 25179 35136 25191 35139
rect 26142 35136 26148 35148
rect 25179 35108 26004 35136
rect 26103 35108 26148 35136
rect 25179 35105 25191 35108
rect 25133 35099 25191 35105
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 2133 35071 2191 35077
rect 2133 35037 2145 35071
rect 2179 35068 2191 35071
rect 2314 35068 2320 35080
rect 2179 35040 2320 35068
rect 2179 35037 2191 35040
rect 2133 35031 2191 35037
rect 2314 35028 2320 35040
rect 2372 35028 2378 35080
rect 14734 35068 14740 35080
rect 14695 35040 14740 35068
rect 14734 35028 14740 35040
rect 14792 35028 14798 35080
rect 19521 35071 19579 35077
rect 19521 35037 19533 35071
rect 19567 35068 19579 35071
rect 20622 35068 20628 35080
rect 19567 35040 20628 35068
rect 19567 35037 19579 35040
rect 19521 35031 19579 35037
rect 20622 35028 20628 35040
rect 20680 35028 20686 35080
rect 20901 35071 20959 35077
rect 20901 35037 20913 35071
rect 20947 35068 20959 35071
rect 21082 35068 21088 35080
rect 20947 35040 21088 35068
rect 20947 35037 20959 35040
rect 20901 35031 20959 35037
rect 21082 35028 21088 35040
rect 21140 35028 21146 35080
rect 25222 35068 25228 35080
rect 25183 35040 25228 35068
rect 25222 35028 25228 35040
rect 25280 35028 25286 35080
rect 25976 35068 26004 35108
rect 26142 35096 26148 35108
rect 26200 35096 26206 35148
rect 26421 35139 26479 35145
rect 26421 35105 26433 35139
rect 26467 35136 26479 35139
rect 27614 35136 27620 35148
rect 26467 35108 27620 35136
rect 26467 35105 26479 35108
rect 26421 35099 26479 35105
rect 27614 35096 27620 35108
rect 27672 35096 27678 35148
rect 28460 35068 28488 35244
rect 29638 35232 29644 35244
rect 29696 35232 29702 35284
rect 29549 35071 29607 35077
rect 29549 35068 29561 35071
rect 25976 35040 26188 35068
rect 28460 35040 29561 35068
rect 15010 35000 15016 35012
rect 14971 34972 15016 35000
rect 15010 34960 15016 34972
rect 15068 34960 15074 35012
rect 16390 35000 16396 35012
rect 16238 34972 16396 35000
rect 16390 34960 16396 34972
rect 16448 34960 16454 35012
rect 17221 35003 17279 35009
rect 17221 34969 17233 35003
rect 17267 34969 17279 35003
rect 17221 34963 17279 34969
rect 1397 34935 1455 34941
rect 1397 34901 1409 34935
rect 1443 34932 1455 34935
rect 1486 34932 1492 34944
rect 1443 34904 1492 34932
rect 1443 34901 1455 34904
rect 1397 34895 1455 34901
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 16485 34935 16543 34941
rect 16485 34901 16497 34935
rect 16531 34932 16543 34935
rect 17126 34932 17132 34944
rect 16531 34904 17132 34932
rect 16531 34901 16543 34904
rect 16485 34895 16543 34901
rect 17126 34892 17132 34904
rect 17184 34892 17190 34944
rect 17236 34932 17264 34963
rect 17678 34960 17684 35012
rect 17736 34960 17742 35012
rect 20162 35000 20168 35012
rect 19812 34972 20168 35000
rect 19812 34932 19840 34972
rect 20162 34960 20168 34972
rect 20220 34960 20226 35012
rect 21818 35000 21824 35012
rect 21779 34972 21824 35000
rect 21818 34960 21824 34972
rect 21876 34960 21882 35012
rect 22462 34960 22468 35012
rect 22520 34960 22526 35012
rect 24946 35000 24952 35012
rect 24859 34972 24952 35000
rect 24946 34960 24952 34972
rect 25004 35000 25010 35012
rect 25958 35000 25964 35012
rect 25004 34972 25964 35000
rect 25004 34960 25010 34972
rect 25958 34960 25964 34972
rect 26016 34960 26022 35012
rect 26160 34944 26188 35040
rect 29549 35037 29561 35040
rect 29595 35068 29607 35071
rect 31113 35071 31171 35077
rect 31113 35068 31125 35071
rect 29595 35040 31125 35068
rect 29595 35037 29607 35040
rect 29549 35031 29607 35037
rect 31113 35037 31125 35040
rect 31159 35068 31171 35071
rect 31754 35068 31760 35080
rect 31159 35040 31760 35068
rect 31159 35037 31171 35040
rect 31113 35031 31171 35037
rect 31754 35028 31760 35040
rect 31812 35028 31818 35080
rect 47302 35068 47308 35080
rect 47263 35040 47308 35068
rect 47302 35028 47308 35040
rect 47360 35028 47366 35080
rect 47486 35028 47492 35080
rect 47544 35068 47550 35080
rect 47581 35071 47639 35077
rect 47581 35068 47593 35071
rect 47544 35040 47593 35068
rect 47544 35028 47550 35040
rect 47581 35037 47593 35040
rect 47627 35037 47639 35071
rect 47581 35031 47639 35037
rect 27154 34960 27160 35012
rect 27212 34960 27218 35012
rect 17236 34904 19840 34932
rect 19889 34935 19947 34941
rect 19889 34901 19901 34935
rect 19935 34932 19947 34935
rect 20346 34932 20352 34944
rect 19935 34904 20352 34932
rect 19935 34901 19947 34904
rect 19889 34895 19947 34901
rect 20346 34892 20352 34904
rect 20404 34892 20410 34944
rect 20990 34932 20996 34944
rect 20951 34904 20996 34932
rect 20990 34892 20996 34904
rect 21048 34892 21054 34944
rect 23290 34932 23296 34944
rect 23251 34904 23296 34932
rect 23290 34892 23296 34904
rect 23348 34892 23354 34944
rect 25406 34932 25412 34944
rect 25367 34904 25412 34932
rect 25406 34892 25412 34904
rect 25464 34892 25470 34944
rect 26142 34932 26148 34944
rect 26055 34904 26148 34932
rect 26142 34892 26148 34904
rect 26200 34932 26206 34944
rect 27893 34935 27951 34941
rect 27893 34932 27905 34935
rect 26200 34904 27905 34932
rect 26200 34892 26206 34904
rect 27893 34901 27905 34904
rect 27939 34901 27951 34935
rect 31202 34932 31208 34944
rect 31163 34904 31208 34932
rect 27893 34895 27951 34901
rect 31202 34892 31208 34904
rect 31260 34892 31266 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 17129 34731 17187 34737
rect 17129 34697 17141 34731
rect 17175 34728 17187 34731
rect 17678 34728 17684 34740
rect 17175 34700 17684 34728
rect 17175 34697 17187 34700
rect 17129 34691 17187 34697
rect 17678 34688 17684 34700
rect 17736 34688 17742 34740
rect 18509 34731 18567 34737
rect 18509 34728 18521 34731
rect 17788 34700 18521 34728
rect 15010 34620 15016 34672
rect 15068 34660 15074 34672
rect 17788 34660 17816 34700
rect 18509 34697 18521 34700
rect 18555 34697 18567 34731
rect 18509 34691 18567 34697
rect 19168 34700 21772 34728
rect 18046 34660 18052 34672
rect 15068 34632 17816 34660
rect 17880 34632 18052 34660
rect 15068 34620 15074 34632
rect 15838 34592 15844 34604
rect 15799 34564 15844 34592
rect 15838 34552 15844 34564
rect 15896 34552 15902 34604
rect 16114 34552 16120 34604
rect 16172 34592 16178 34604
rect 17037 34595 17095 34601
rect 17037 34592 17049 34595
rect 16172 34564 17049 34592
rect 16172 34552 16178 34564
rect 17037 34561 17049 34564
rect 17083 34561 17095 34595
rect 17037 34555 17095 34561
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34592 17831 34595
rect 17880 34592 17908 34632
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 19168 34660 19196 34700
rect 19978 34660 19984 34672
rect 18248 34632 19196 34660
rect 17819 34564 17908 34592
rect 17957 34595 18015 34601
rect 17819 34561 17831 34564
rect 17773 34555 17831 34561
rect 17957 34561 17969 34595
rect 18003 34592 18015 34595
rect 18248 34592 18276 34632
rect 18003 34564 18276 34592
rect 18325 34595 18383 34601
rect 18003 34561 18015 34564
rect 17957 34555 18015 34561
rect 18325 34561 18337 34595
rect 18371 34561 18383 34595
rect 18966 34592 18972 34604
rect 18927 34564 18972 34592
rect 18325 34555 18383 34561
rect 17126 34484 17132 34536
rect 17184 34524 17190 34536
rect 18049 34527 18107 34533
rect 18049 34524 18061 34527
rect 17184 34496 18061 34524
rect 17184 34484 17190 34496
rect 17972 34468 18000 34496
rect 18049 34493 18061 34496
rect 18095 34493 18107 34527
rect 18049 34487 18107 34493
rect 18138 34484 18144 34536
rect 18196 34524 18202 34536
rect 18340 34524 18368 34555
rect 18966 34552 18972 34564
rect 19024 34552 19030 34604
rect 19168 34601 19196 34632
rect 19536 34632 19984 34660
rect 19536 34604 19564 34632
rect 19978 34620 19984 34632
rect 20036 34620 20042 34672
rect 20254 34620 20260 34672
rect 20312 34660 20318 34672
rect 21744 34660 21772 34700
rect 21818 34688 21824 34740
rect 21876 34728 21882 34740
rect 22557 34731 22615 34737
rect 22557 34728 22569 34731
rect 21876 34700 22569 34728
rect 21876 34688 21882 34700
rect 22557 34697 22569 34700
rect 22603 34697 22615 34731
rect 22557 34691 22615 34697
rect 23106 34688 23112 34740
rect 23164 34728 23170 34740
rect 26050 34728 26056 34740
rect 23164 34700 26056 34728
rect 23164 34688 23170 34700
rect 26050 34688 26056 34700
rect 26108 34728 26114 34740
rect 28810 34728 28816 34740
rect 26108 34700 28816 34728
rect 26108 34688 26114 34700
rect 28810 34688 28816 34700
rect 28868 34688 28874 34740
rect 28994 34728 29000 34740
rect 28955 34700 29000 34728
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 24762 34660 24768 34672
rect 20312 34632 20668 34660
rect 21744 34632 24768 34660
rect 20312 34620 20318 34632
rect 19153 34595 19211 34601
rect 19153 34561 19165 34595
rect 19199 34561 19211 34595
rect 19153 34555 19211 34561
rect 19260 34564 19472 34592
rect 18196 34496 18241 34524
rect 18340 34496 19012 34524
rect 18196 34484 18202 34496
rect 17954 34416 17960 34468
rect 18012 34416 18018 34468
rect 16025 34391 16083 34397
rect 16025 34357 16037 34391
rect 16071 34388 16083 34391
rect 16114 34388 16120 34400
rect 16071 34360 16120 34388
rect 16071 34357 16083 34360
rect 16025 34351 16083 34357
rect 16114 34348 16120 34360
rect 16172 34348 16178 34400
rect 18984 34388 19012 34496
rect 19058 34484 19064 34536
rect 19116 34524 19122 34536
rect 19260 34533 19288 34564
rect 19245 34527 19303 34533
rect 19245 34524 19257 34527
rect 19116 34496 19257 34524
rect 19116 34484 19122 34496
rect 19245 34493 19257 34496
rect 19291 34493 19303 34527
rect 19245 34487 19303 34493
rect 19337 34527 19395 34533
rect 19337 34493 19349 34527
rect 19383 34493 19395 34527
rect 19444 34524 19472 34564
rect 19518 34552 19524 34604
rect 19576 34592 19582 34604
rect 19705 34595 19763 34601
rect 19576 34564 19669 34592
rect 19576 34552 19582 34564
rect 19705 34561 19717 34595
rect 19751 34592 19763 34595
rect 20162 34592 20168 34604
rect 19751 34564 20168 34592
rect 19751 34561 19763 34564
rect 19705 34555 19763 34561
rect 20162 34552 20168 34564
rect 20220 34552 20226 34604
rect 20349 34595 20407 34601
rect 20349 34561 20361 34595
rect 20395 34561 20407 34595
rect 20349 34555 20407 34561
rect 20364 34524 20392 34555
rect 20438 34552 20444 34604
rect 20496 34592 20502 34604
rect 20640 34601 20668 34632
rect 20533 34595 20591 34601
rect 20533 34592 20545 34595
rect 20496 34564 20545 34592
rect 20496 34552 20502 34564
rect 20533 34561 20545 34564
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20625 34595 20683 34601
rect 20625 34561 20637 34595
rect 20671 34561 20683 34595
rect 21818 34592 21824 34604
rect 21779 34564 21824 34592
rect 20625 34555 20683 34561
rect 21818 34552 21824 34564
rect 21876 34552 21882 34604
rect 22008 34601 22036 34632
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 27065 34663 27123 34669
rect 27065 34660 27077 34663
rect 25714 34632 27077 34660
rect 27065 34629 27077 34632
rect 27111 34629 27123 34663
rect 27065 34623 27123 34629
rect 27522 34620 27528 34672
rect 27580 34660 27586 34672
rect 27580 34632 29868 34660
rect 27580 34620 27586 34632
rect 22005 34595 22063 34601
rect 22005 34561 22017 34595
rect 22051 34561 22063 34595
rect 22186 34592 22192 34604
rect 22147 34564 22192 34592
rect 22005 34555 22063 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22373 34595 22431 34601
rect 22373 34561 22385 34595
rect 22419 34592 22431 34595
rect 22922 34592 22928 34604
rect 22419 34564 22928 34592
rect 22419 34561 22431 34564
rect 22373 34555 22431 34561
rect 22922 34552 22928 34564
rect 22980 34552 22986 34604
rect 23014 34552 23020 34604
rect 23072 34592 23078 34604
rect 24213 34595 24271 34601
rect 24213 34592 24225 34595
rect 23072 34564 24225 34592
rect 23072 34552 23078 34564
rect 24213 34561 24225 34564
rect 24259 34561 24271 34595
rect 26970 34592 26976 34604
rect 26931 34564 26976 34592
rect 24213 34555 24271 34561
rect 26970 34552 26976 34564
rect 27028 34552 27034 34604
rect 28261 34595 28319 34601
rect 28261 34561 28273 34595
rect 28307 34561 28319 34595
rect 28442 34592 28448 34604
rect 28403 34564 28448 34592
rect 28261 34555 28319 34561
rect 19444 34496 20392 34524
rect 22097 34527 22155 34533
rect 19337 34487 19395 34493
rect 22097 34493 22109 34527
rect 22143 34524 22155 34527
rect 23290 34524 23296 34536
rect 22143 34496 23296 34524
rect 22143 34493 22155 34496
rect 22097 34487 22155 34493
rect 19352 34456 19380 34487
rect 23290 34484 23296 34496
rect 23348 34484 23354 34536
rect 24486 34524 24492 34536
rect 24447 34496 24492 34524
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 28276 34524 28304 34555
rect 28442 34552 28448 34564
rect 28500 34552 28506 34604
rect 28626 34592 28632 34604
rect 28587 34564 28632 34592
rect 28626 34552 28632 34564
rect 28684 34552 28690 34604
rect 28810 34592 28816 34604
rect 28771 34564 28816 34592
rect 28810 34552 28816 34564
rect 28868 34552 28874 34604
rect 29840 34601 29868 34632
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 31202 34552 31208 34604
rect 31260 34552 31266 34604
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 28537 34527 28595 34533
rect 28276 34496 28488 34524
rect 20438 34456 20444 34468
rect 19352 34428 20444 34456
rect 20438 34416 20444 34428
rect 20496 34416 20502 34468
rect 25958 34456 25964 34468
rect 25919 34428 25964 34456
rect 25958 34416 25964 34428
rect 26016 34416 26022 34468
rect 28460 34456 28488 34496
rect 28537 34493 28549 34527
rect 28583 34524 28595 34527
rect 29730 34524 29736 34536
rect 28583 34496 29736 34524
rect 28583 34493 28595 34496
rect 28537 34487 28595 34493
rect 29730 34484 29736 34496
rect 29788 34484 29794 34536
rect 30098 34524 30104 34536
rect 30059 34496 30104 34524
rect 30098 34484 30104 34496
rect 30156 34484 30162 34536
rect 28994 34456 29000 34468
rect 28460 34428 29000 34456
rect 28994 34416 29000 34428
rect 29052 34416 29058 34468
rect 19518 34388 19524 34400
rect 18984 34360 19524 34388
rect 19518 34348 19524 34360
rect 19576 34348 19582 34400
rect 20162 34388 20168 34400
rect 20123 34360 20168 34388
rect 20162 34348 20168 34360
rect 20220 34348 20226 34400
rect 29730 34348 29736 34400
rect 29788 34388 29794 34400
rect 30190 34388 30196 34400
rect 29788 34360 30196 34388
rect 29788 34348 29794 34360
rect 30190 34348 30196 34360
rect 30248 34388 30254 34400
rect 31573 34391 31631 34397
rect 31573 34388 31585 34391
rect 30248 34360 31585 34388
rect 30248 34348 30254 34360
rect 31573 34357 31585 34360
rect 31619 34357 31631 34391
rect 47946 34388 47952 34400
rect 47907 34360 47952 34388
rect 31573 34351 31631 34357
rect 47946 34348 47952 34360
rect 48004 34348 48010 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 16390 34184 16396 34196
rect 16351 34156 16396 34184
rect 16390 34144 16396 34156
rect 16448 34144 16454 34196
rect 24486 34144 24492 34196
rect 24544 34184 24550 34196
rect 25225 34187 25283 34193
rect 25225 34184 25237 34187
rect 24544 34156 25237 34184
rect 24544 34144 24550 34156
rect 25225 34153 25237 34156
rect 25271 34153 25283 34187
rect 25225 34147 25283 34153
rect 28721 34187 28779 34193
rect 28721 34153 28733 34187
rect 28767 34153 28779 34187
rect 28994 34184 29000 34196
rect 28955 34156 29000 34184
rect 28721 34147 28779 34153
rect 24762 34076 24768 34128
rect 24820 34116 24826 34128
rect 27801 34119 27859 34125
rect 27801 34116 27813 34119
rect 24820 34088 27813 34116
rect 24820 34076 24826 34088
rect 27801 34085 27813 34088
rect 27847 34116 27859 34119
rect 28442 34116 28448 34128
rect 27847 34088 28448 34116
rect 27847 34085 27859 34088
rect 27801 34079 27859 34085
rect 28442 34076 28448 34088
rect 28500 34076 28506 34128
rect 28534 34076 28540 34128
rect 28592 34116 28598 34128
rect 28736 34116 28764 34147
rect 28994 34144 29000 34156
rect 29052 34144 29058 34196
rect 29730 34144 29736 34196
rect 29788 34144 29794 34196
rect 30098 34144 30104 34196
rect 30156 34184 30162 34196
rect 30285 34187 30343 34193
rect 30285 34184 30297 34187
rect 30156 34156 30297 34184
rect 30156 34144 30162 34156
rect 30285 34153 30297 34156
rect 30331 34153 30343 34187
rect 30285 34147 30343 34153
rect 30650 34144 30656 34196
rect 30708 34184 30714 34196
rect 31113 34187 31171 34193
rect 31113 34184 31125 34187
rect 30708 34156 31125 34184
rect 30708 34144 30714 34156
rect 31113 34153 31125 34156
rect 31159 34153 31171 34187
rect 31113 34147 31171 34153
rect 29638 34116 29644 34128
rect 28592 34088 29644 34116
rect 28592 34076 28598 34088
rect 29638 34076 29644 34088
rect 29696 34076 29702 34128
rect 19334 34008 19340 34060
rect 19392 34048 19398 34060
rect 20165 34051 20223 34057
rect 20165 34048 20177 34051
rect 19392 34020 20177 34048
rect 19392 34008 19398 34020
rect 20165 34017 20177 34020
rect 20211 34048 20223 34051
rect 21450 34048 21456 34060
rect 20211 34020 21456 34048
rect 20211 34017 20223 34020
rect 20165 34011 20223 34017
rect 21450 34008 21456 34020
rect 21508 34008 21514 34060
rect 24946 34048 24952 34060
rect 24907 34020 24952 34048
rect 24946 34008 24952 34020
rect 25004 34048 25010 34060
rect 25222 34048 25228 34060
rect 25004 34020 25228 34048
rect 25004 34008 25010 34020
rect 25222 34008 25228 34020
rect 25280 34008 25286 34060
rect 28460 34048 28488 34076
rect 28721 34051 28779 34057
rect 28460 34020 28580 34048
rect 16114 33940 16120 33992
rect 16172 33980 16178 33992
rect 16301 33983 16359 33989
rect 16301 33980 16313 33983
rect 16172 33952 16313 33980
rect 16172 33940 16178 33952
rect 16301 33949 16313 33952
rect 16347 33949 16359 33983
rect 25038 33980 25044 33992
rect 24999 33952 25044 33980
rect 16301 33943 16359 33949
rect 25038 33940 25044 33952
rect 25096 33940 25102 33992
rect 25406 33940 25412 33992
rect 25464 33980 25470 33992
rect 25685 33983 25743 33989
rect 25685 33980 25697 33983
rect 25464 33952 25697 33980
rect 25464 33940 25470 33952
rect 25685 33949 25697 33952
rect 25731 33949 25743 33983
rect 25685 33943 25743 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33980 27675 33983
rect 27706 33980 27712 33992
rect 27663 33952 27712 33980
rect 27663 33949 27675 33952
rect 27617 33943 27675 33949
rect 27706 33940 27712 33952
rect 27764 33940 27770 33992
rect 28442 33980 28448 33992
rect 28403 33952 28448 33980
rect 28442 33940 28448 33952
rect 28500 33940 28506 33992
rect 20441 33915 20499 33921
rect 20441 33881 20453 33915
rect 20487 33912 20499 33915
rect 20714 33912 20720 33924
rect 20487 33884 20720 33912
rect 20487 33881 20499 33884
rect 20441 33875 20499 33881
rect 20714 33872 20720 33884
rect 20772 33872 20778 33924
rect 20990 33872 20996 33924
rect 21048 33872 21054 33924
rect 23382 33872 23388 33924
rect 23440 33912 23446 33924
rect 23440 33884 24716 33912
rect 23440 33872 23446 33884
rect 20622 33804 20628 33856
rect 20680 33844 20686 33856
rect 21910 33844 21916 33856
rect 20680 33816 21916 33844
rect 20680 33804 20686 33816
rect 21910 33804 21916 33816
rect 21968 33804 21974 33856
rect 23750 33804 23756 33856
rect 23808 33844 23814 33856
rect 24581 33847 24639 33853
rect 24581 33844 24593 33847
rect 23808 33816 24593 33844
rect 23808 33804 23814 33816
rect 24581 33813 24593 33816
rect 24627 33813 24639 33847
rect 24688 33844 24716 33884
rect 24762 33872 24768 33924
rect 24820 33912 24826 33924
rect 25869 33915 25927 33921
rect 25869 33912 25881 33915
rect 24820 33884 25881 33912
rect 24820 33872 24826 33884
rect 25869 33881 25881 33884
rect 25915 33912 25927 33915
rect 27890 33912 27896 33924
rect 25915 33884 27896 33912
rect 25915 33881 25927 33884
rect 25869 33875 25927 33881
rect 27890 33872 27896 33884
rect 27948 33872 27954 33924
rect 28552 33912 28580 34020
rect 28721 34017 28733 34051
rect 28767 34048 28779 34051
rect 29178 34048 29184 34060
rect 28767 34020 29184 34048
rect 28767 34017 28779 34020
rect 28721 34011 28779 34017
rect 29178 34008 29184 34020
rect 29236 34008 29242 34060
rect 29748 34048 29776 34144
rect 29819 34051 29877 34057
rect 29819 34048 29831 34051
rect 29748 34020 29831 34048
rect 29819 34017 29831 34020
rect 29865 34017 29877 34051
rect 29819 34011 29877 34017
rect 31018 34008 31024 34060
rect 31076 34048 31082 34060
rect 31205 34051 31263 34057
rect 31205 34048 31217 34051
rect 31076 34020 31217 34048
rect 31076 34008 31082 34020
rect 31205 34017 31217 34020
rect 31251 34017 31263 34051
rect 31205 34011 31263 34017
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34048 46351 34051
rect 47946 34048 47952 34060
rect 46339 34020 47952 34048
rect 46339 34017 46351 34020
rect 46293 34011 46351 34017
rect 47946 34008 47952 34020
rect 48004 34008 48010 34060
rect 29454 33940 29460 33992
rect 29512 33958 29518 33992
rect 29549 33961 29607 33967
rect 29549 33958 29561 33961
rect 29512 33940 29561 33958
rect 29472 33930 29561 33940
rect 29549 33927 29561 33930
rect 29595 33927 29607 33961
rect 29730 33940 29736 33992
rect 29788 33978 29794 33992
rect 29917 33983 29975 33989
rect 29788 33950 29831 33978
rect 29788 33940 29794 33950
rect 29917 33949 29929 33983
rect 29963 33958 29975 33983
rect 29963 33949 30052 33958
rect 29917 33943 30052 33949
rect 29932 33930 30052 33943
rect 30098 33940 30104 33992
rect 30156 33980 30162 33992
rect 30926 33980 30932 33992
rect 30156 33952 30201 33980
rect 30887 33952 30932 33980
rect 30156 33940 30162 33952
rect 30926 33940 30932 33952
rect 30984 33940 30990 33992
rect 31754 33980 31760 33992
rect 31715 33952 31760 33980
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 29270 33912 29276 33924
rect 28552 33884 29276 33912
rect 29270 33872 29276 33884
rect 29328 33872 29334 33924
rect 29549 33921 29607 33927
rect 30024 33912 30052 33930
rect 30024 33884 30696 33912
rect 26053 33847 26111 33853
rect 26053 33844 26065 33847
rect 24688 33816 26065 33844
rect 24581 33807 24639 33813
rect 26053 33813 26065 33816
rect 26099 33813 26111 33847
rect 26053 33807 26111 33813
rect 26970 33804 26976 33856
rect 27028 33844 27034 33856
rect 30558 33844 30564 33856
rect 27028 33816 30564 33844
rect 27028 33804 27034 33816
rect 30558 33804 30564 33816
rect 30616 33804 30622 33856
rect 30668 33853 30696 33884
rect 30742 33872 30748 33924
rect 30800 33912 30806 33924
rect 46477 33915 46535 33921
rect 30800 33884 30845 33912
rect 30800 33872 30806 33884
rect 46477 33881 46489 33915
rect 46523 33912 46535 33915
rect 47486 33912 47492 33924
rect 46523 33884 47492 33912
rect 46523 33881 46535 33884
rect 46477 33875 46535 33881
rect 47486 33872 47492 33884
rect 47544 33872 47550 33924
rect 48133 33915 48191 33921
rect 48133 33881 48145 33915
rect 48179 33881 48191 33915
rect 48133 33875 48191 33881
rect 30653 33847 30711 33853
rect 30653 33813 30665 33847
rect 30699 33844 30711 33847
rect 31662 33844 31668 33856
rect 30699 33816 31668 33844
rect 30699 33813 30711 33816
rect 30653 33807 30711 33813
rect 31662 33804 31668 33816
rect 31720 33804 31726 33856
rect 31849 33847 31907 33853
rect 31849 33813 31861 33847
rect 31895 33844 31907 33847
rect 31938 33844 31944 33856
rect 31895 33816 31944 33844
rect 31895 33813 31907 33816
rect 31849 33807 31907 33813
rect 31938 33804 31944 33816
rect 31996 33804 32002 33856
rect 45830 33804 45836 33856
rect 45888 33844 45894 33856
rect 48148 33844 48176 33875
rect 45888 33816 48176 33844
rect 45888 33804 45894 33816
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 18046 33640 18052 33652
rect 18007 33612 18052 33640
rect 18046 33600 18052 33612
rect 18104 33600 18110 33652
rect 18966 33600 18972 33652
rect 19024 33640 19030 33652
rect 19521 33643 19579 33649
rect 19521 33640 19533 33643
rect 19024 33612 19533 33640
rect 19024 33600 19030 33612
rect 19521 33609 19533 33612
rect 19567 33609 19579 33643
rect 20530 33640 20536 33652
rect 20491 33612 20536 33640
rect 19521 33603 19579 33609
rect 20530 33600 20536 33612
rect 20588 33600 20594 33652
rect 21818 33600 21824 33652
rect 21876 33640 21882 33652
rect 22373 33643 22431 33649
rect 22373 33640 22385 33643
rect 21876 33612 22385 33640
rect 21876 33600 21882 33612
rect 22373 33609 22385 33612
rect 22419 33609 22431 33643
rect 23750 33640 23756 33652
rect 22373 33603 22431 33609
rect 22940 33612 23428 33640
rect 23711 33612 23756 33640
rect 22940 33572 22968 33612
rect 23290 33572 23296 33584
rect 17696 33544 22968 33572
rect 23032 33544 23296 33572
rect 17696 33513 17724 33544
rect 17681 33507 17739 33513
rect 17681 33473 17693 33507
rect 17727 33473 17739 33507
rect 17681 33467 17739 33473
rect 18969 33507 19027 33513
rect 18969 33473 18981 33507
rect 19015 33504 19027 33507
rect 19518 33504 19524 33516
rect 19015 33476 19524 33504
rect 19015 33473 19027 33476
rect 18969 33467 19027 33473
rect 19518 33464 19524 33476
rect 19576 33464 19582 33516
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33504 20223 33507
rect 20254 33504 20260 33516
rect 20211 33476 20260 33504
rect 20211 33473 20223 33476
rect 20165 33467 20223 33473
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 20349 33510 20407 33513
rect 20349 33507 20484 33510
rect 20349 33473 20361 33507
rect 20395 33504 20484 33507
rect 20622 33504 20628 33516
rect 20395 33482 20628 33504
rect 20395 33473 20407 33482
rect 20456 33476 20628 33482
rect 20349 33467 20407 33473
rect 20622 33464 20628 33476
rect 20680 33504 20686 33516
rect 20806 33504 20812 33516
rect 20680 33476 20812 33504
rect 20680 33464 20686 33476
rect 20806 33464 20812 33476
rect 20864 33464 20870 33516
rect 21818 33504 21824 33516
rect 21731 33476 21824 33504
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2038 33436 2044 33448
rect 1719 33408 2044 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2038 33396 2044 33408
rect 2096 33396 2102 33448
rect 17770 33436 17776 33448
rect 17731 33408 17776 33436
rect 17770 33396 17776 33408
rect 17828 33396 17834 33448
rect 19245 33440 19303 33445
rect 19245 33439 19294 33440
rect 19245 33405 19257 33439
rect 19291 33405 19294 33439
rect 19245 33399 19294 33405
rect 19288 33388 19294 33399
rect 19346 33436 19352 33440
rect 20272 33436 20300 33464
rect 21744 33436 21772 33476
rect 21818 33464 21824 33476
rect 21876 33464 21882 33516
rect 22186 33504 22192 33516
rect 22147 33476 22192 33504
rect 22186 33464 22192 33476
rect 22244 33464 22250 33516
rect 23032 33513 23060 33544
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 23400 33572 23428 33612
rect 23750 33600 23756 33612
rect 23808 33600 23814 33652
rect 23934 33640 23940 33652
rect 23895 33612 23940 33640
rect 23934 33600 23940 33612
rect 23992 33600 23998 33652
rect 24412 33612 24992 33640
rect 24412 33572 24440 33612
rect 23400 33544 24440 33572
rect 23017 33507 23075 33513
rect 23017 33473 23029 33507
rect 23063 33473 23075 33507
rect 23017 33467 23075 33473
rect 23842 33464 23848 33516
rect 23900 33513 23906 33516
rect 23900 33507 23936 33513
rect 23924 33473 23936 33507
rect 23900 33467 23936 33473
rect 23900 33464 23906 33467
rect 19346 33408 19385 33436
rect 20272 33408 21772 33436
rect 19346 33388 19352 33408
rect 23198 33396 23204 33448
rect 23256 33436 23262 33448
rect 24412 33445 24440 33544
rect 24762 33532 24768 33584
rect 24820 33572 24826 33584
rect 24857 33575 24915 33581
rect 24857 33572 24869 33575
rect 24820 33544 24869 33572
rect 24820 33532 24826 33544
rect 24857 33541 24869 33544
rect 24903 33541 24915 33575
rect 24964 33572 24992 33612
rect 25038 33600 25044 33652
rect 25096 33640 25102 33652
rect 27249 33643 27307 33649
rect 27249 33640 27261 33643
rect 25096 33612 27261 33640
rect 25096 33600 25102 33612
rect 27249 33609 27261 33612
rect 27295 33609 27307 33643
rect 27249 33603 27307 33609
rect 28721 33643 28779 33649
rect 28721 33609 28733 33643
rect 28767 33640 28779 33643
rect 29454 33640 29460 33652
rect 28767 33612 29460 33640
rect 28767 33609 28779 33612
rect 28721 33603 28779 33609
rect 29454 33600 29460 33612
rect 29512 33600 29518 33652
rect 28810 33572 28816 33584
rect 24964 33544 28816 33572
rect 24857 33535 24915 33541
rect 28810 33532 28816 33544
rect 28868 33532 28874 33584
rect 29012 33544 30052 33572
rect 25133 33507 25191 33513
rect 24872 33476 25084 33504
rect 23293 33439 23351 33445
rect 23293 33436 23305 33439
rect 23256 33408 23305 33436
rect 23256 33396 23262 33408
rect 23293 33405 23305 33408
rect 23339 33405 23351 33439
rect 23293 33399 23351 33405
rect 24397 33439 24455 33445
rect 24397 33405 24409 33439
rect 24443 33405 24455 33439
rect 24397 33399 24455 33405
rect 22833 33371 22891 33377
rect 22833 33368 22845 33371
rect 22204 33340 22845 33368
rect 17678 33300 17684 33312
rect 17639 33272 17684 33300
rect 17678 33260 17684 33272
rect 17736 33260 17742 33312
rect 19337 33303 19395 33309
rect 19337 33269 19349 33303
rect 19383 33300 19395 33303
rect 20162 33300 20168 33312
rect 19383 33272 20168 33300
rect 19383 33269 19395 33272
rect 19337 33263 19395 33269
rect 20162 33260 20168 33272
rect 20220 33260 20226 33312
rect 22204 33309 22232 33340
rect 22833 33337 22845 33340
rect 22879 33337 22891 33371
rect 22833 33331 22891 33337
rect 23014 33328 23020 33380
rect 23072 33368 23078 33380
rect 24305 33371 24363 33377
rect 23072 33340 23520 33368
rect 23072 33328 23078 33340
rect 22189 33303 22247 33309
rect 22189 33269 22201 33303
rect 22235 33269 22247 33303
rect 22189 33263 22247 33269
rect 23106 33260 23112 33312
rect 23164 33300 23170 33312
rect 23201 33303 23259 33309
rect 23201 33300 23213 33303
rect 23164 33272 23213 33300
rect 23164 33260 23170 33272
rect 23201 33269 23213 33272
rect 23247 33300 23259 33303
rect 23382 33300 23388 33312
rect 23247 33272 23388 33300
rect 23247 33269 23259 33272
rect 23201 33263 23259 33269
rect 23382 33260 23388 33272
rect 23440 33260 23446 33312
rect 23492 33300 23520 33340
rect 24305 33337 24317 33371
rect 24351 33368 24363 33371
rect 24872 33368 24900 33476
rect 24949 33439 25007 33445
rect 24949 33405 24961 33439
rect 24995 33405 25007 33439
rect 24949 33399 25007 33405
rect 24351 33340 24900 33368
rect 24351 33337 24363 33340
rect 24305 33331 24363 33337
rect 24964 33300 24992 33399
rect 25056 33368 25084 33476
rect 25133 33473 25145 33507
rect 25179 33504 25191 33507
rect 25222 33504 25228 33516
rect 25179 33476 25228 33504
rect 25179 33473 25191 33476
rect 25133 33467 25191 33473
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25774 33504 25780 33516
rect 25332 33476 25780 33504
rect 25332 33377 25360 33476
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33504 26019 33507
rect 26142 33504 26148 33516
rect 26007 33476 26148 33504
rect 26007 33473 26019 33476
rect 25961 33467 26019 33473
rect 26142 33464 26148 33476
rect 26200 33464 26206 33516
rect 26970 33504 26976 33516
rect 26931 33476 26976 33504
rect 26970 33464 26976 33476
rect 27028 33464 27034 33516
rect 27890 33504 27896 33516
rect 27851 33476 27896 33504
rect 27890 33464 27896 33476
rect 27948 33464 27954 33516
rect 28074 33504 28080 33516
rect 28035 33476 28080 33504
rect 28074 33464 28080 33476
rect 28132 33464 28138 33516
rect 28442 33464 28448 33516
rect 28500 33504 28506 33516
rect 29012 33513 29040 33544
rect 28905 33507 28963 33513
rect 28905 33504 28917 33507
rect 28500 33476 28917 33504
rect 28500 33464 28506 33476
rect 28905 33473 28917 33476
rect 28951 33473 28963 33507
rect 28905 33467 28963 33473
rect 28997 33507 29055 33513
rect 28997 33473 29009 33507
rect 29043 33473 29055 33507
rect 28997 33467 29055 33473
rect 29181 33507 29239 33513
rect 29181 33473 29193 33507
rect 29227 33473 29239 33507
rect 29181 33467 29239 33473
rect 27249 33439 27307 33445
rect 27249 33405 27261 33439
rect 27295 33436 27307 33439
rect 27706 33436 27712 33448
rect 27295 33408 27712 33436
rect 27295 33405 27307 33408
rect 27249 33399 27307 33405
rect 27706 33396 27712 33408
rect 27764 33396 27770 33448
rect 27985 33439 28043 33445
rect 27985 33405 27997 33439
rect 28031 33436 28043 33439
rect 28644 33436 28856 33447
rect 29196 33436 29224 33467
rect 29270 33464 29276 33516
rect 29328 33504 29334 33516
rect 29730 33504 29736 33516
rect 29328 33476 29373 33504
rect 29691 33476 29736 33504
rect 29328 33464 29334 33476
rect 29730 33464 29736 33476
rect 29788 33464 29794 33516
rect 30024 33513 30052 33544
rect 30098 33532 30104 33584
rect 30156 33572 30162 33584
rect 30926 33572 30932 33584
rect 30156 33544 30932 33572
rect 30156 33532 30162 33544
rect 30009 33507 30067 33513
rect 30009 33473 30021 33507
rect 30055 33504 30067 33507
rect 30190 33504 30196 33516
rect 30055 33476 30196 33504
rect 30055 33473 30067 33476
rect 30009 33467 30067 33473
rect 30190 33464 30196 33476
rect 30248 33464 30254 33516
rect 30650 33504 30656 33516
rect 30611 33476 30656 33504
rect 30650 33464 30656 33476
rect 30708 33464 30714 33516
rect 30852 33513 30880 33544
rect 30926 33532 30932 33544
rect 30984 33532 30990 33584
rect 30837 33507 30895 33513
rect 30837 33473 30849 33507
rect 30883 33473 30895 33507
rect 47854 33504 47860 33516
rect 47815 33476 47860 33504
rect 30837 33467 30895 33473
rect 47854 33464 47860 33476
rect 47912 33464 47918 33516
rect 28031 33428 28948 33436
rect 29012 33428 29224 33436
rect 28031 33419 29224 33428
rect 28031 33408 28672 33419
rect 28828 33408 29224 33419
rect 29917 33439 29975 33445
rect 28031 33405 28043 33408
rect 27985 33399 28043 33405
rect 28920 33400 29040 33408
rect 29917 33405 29929 33439
rect 29963 33436 29975 33439
rect 30466 33436 30472 33448
rect 29963 33408 30472 33436
rect 29963 33405 29975 33408
rect 29917 33399 29975 33405
rect 25317 33371 25375 33377
rect 25317 33368 25329 33371
rect 25056 33340 25329 33368
rect 25317 33337 25329 33340
rect 25363 33337 25375 33371
rect 25317 33331 25375 33337
rect 27065 33371 27123 33377
rect 27065 33337 27077 33371
rect 27111 33368 27123 33371
rect 28000 33368 28028 33399
rect 30466 33396 30472 33408
rect 30524 33396 30530 33448
rect 27111 33340 28028 33368
rect 27111 33337 27123 33340
rect 27065 33331 27123 33337
rect 28442 33328 28448 33380
rect 28500 33368 28506 33380
rect 29454 33368 29460 33380
rect 28500 33340 29460 33368
rect 28500 33328 28506 33340
rect 29454 33328 29460 33340
rect 29512 33328 29518 33380
rect 30193 33371 30251 33377
rect 30193 33337 30205 33371
rect 30239 33368 30251 33371
rect 30239 33340 30328 33368
rect 30239 33337 30251 33340
rect 30193 33331 30251 33337
rect 30300 33312 30328 33340
rect 30374 33328 30380 33380
rect 30432 33368 30438 33380
rect 31021 33371 31079 33377
rect 31021 33368 31033 33371
rect 30432 33340 31033 33368
rect 30432 33328 30438 33340
rect 31021 33337 31033 33340
rect 31067 33337 31079 33371
rect 31021 33331 31079 33337
rect 25130 33300 25136 33312
rect 23492 33272 24992 33300
rect 25043 33272 25136 33300
rect 25130 33260 25136 33272
rect 25188 33300 25194 33312
rect 25590 33300 25596 33312
rect 25188 33272 25596 33300
rect 25188 33260 25194 33272
rect 25590 33260 25596 33272
rect 25648 33260 25654 33312
rect 25777 33303 25835 33309
rect 25777 33269 25789 33303
rect 25823 33300 25835 33303
rect 25866 33300 25872 33312
rect 25823 33272 25872 33300
rect 25823 33269 25835 33272
rect 25777 33263 25835 33269
rect 25866 33260 25872 33272
rect 25924 33260 25930 33312
rect 27890 33260 27896 33312
rect 27948 33300 27954 33312
rect 29546 33300 29552 33312
rect 27948 33272 29552 33300
rect 27948 33260 27954 33272
rect 29546 33260 29552 33272
rect 29604 33260 29610 33312
rect 30006 33260 30012 33312
rect 30064 33300 30070 33312
rect 30064 33272 30109 33300
rect 30064 33260 30070 33272
rect 30282 33260 30288 33312
rect 30340 33260 30346 33312
rect 30466 33260 30472 33312
rect 30524 33300 30530 33312
rect 30837 33303 30895 33309
rect 30837 33300 30849 33303
rect 30524 33272 30849 33300
rect 30524 33260 30530 33272
rect 30837 33269 30849 33272
rect 30883 33300 30895 33303
rect 30926 33300 30932 33312
rect 30883 33272 30932 33300
rect 30883 33269 30895 33272
rect 30837 33263 30895 33269
rect 30926 33260 30932 33272
rect 30984 33260 30990 33312
rect 44174 33260 44180 33312
rect 44232 33300 44238 33312
rect 48041 33303 48099 33309
rect 48041 33300 48053 33303
rect 44232 33272 48053 33300
rect 44232 33260 44238 33272
rect 48041 33269 48053 33272
rect 48087 33269 48099 33303
rect 48041 33263 48099 33269
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 17405 33099 17463 33105
rect 17405 33065 17417 33099
rect 17451 33096 17463 33099
rect 17678 33096 17684 33108
rect 17451 33068 17684 33096
rect 17451 33065 17463 33068
rect 17405 33059 17463 33065
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 21450 33056 21456 33108
rect 21508 33096 21514 33108
rect 21637 33099 21695 33105
rect 21637 33096 21649 33099
rect 21508 33068 21649 33096
rect 21508 33056 21514 33068
rect 21637 33065 21649 33068
rect 21683 33065 21695 33099
rect 21637 33059 21695 33065
rect 23385 33099 23443 33105
rect 23385 33065 23397 33099
rect 23431 33065 23443 33099
rect 24394 33096 24400 33108
rect 24355 33068 24400 33096
rect 23385 33059 23443 33065
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 15930 32988 15936 33040
rect 15988 33028 15994 33040
rect 17773 33031 17831 33037
rect 17773 33028 17785 33031
rect 15988 33000 17785 33028
rect 15988 32988 15994 33000
rect 17773 32997 17785 33000
rect 17819 33028 17831 33031
rect 20622 33028 20628 33040
rect 17819 33000 19334 33028
rect 20583 33000 20628 33028
rect 17819 32997 17831 33000
rect 17773 32991 17831 32997
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 17954 32960 17960 32972
rect 1397 32923 1455 32929
rect 17604 32932 17960 32960
rect 16666 32892 16672 32904
rect 16627 32864 16672 32892
rect 16666 32852 16672 32864
rect 16724 32852 16730 32904
rect 16942 32892 16948 32904
rect 16903 32864 16948 32892
rect 16942 32852 16948 32864
rect 17000 32852 17006 32904
rect 17604 32901 17632 32932
rect 17954 32920 17960 32932
rect 18012 32960 18018 32972
rect 18230 32960 18236 32972
rect 18012 32932 18236 32960
rect 18012 32920 18018 32932
rect 18230 32920 18236 32932
rect 18288 32960 18294 32972
rect 19306 32960 19334 33000
rect 20622 32988 20628 33000
rect 20680 32988 20686 33040
rect 23400 33028 23428 33059
rect 24394 33056 24400 33068
rect 24452 33056 24458 33108
rect 24854 33096 24860 33108
rect 24815 33068 24860 33096
rect 24854 33056 24860 33068
rect 24912 33056 24918 33108
rect 25774 33056 25780 33108
rect 25832 33096 25838 33108
rect 25961 33099 26019 33105
rect 25961 33096 25973 33099
rect 25832 33068 25973 33096
rect 25832 33056 25838 33068
rect 25961 33065 25973 33068
rect 26007 33065 26019 33099
rect 25961 33059 26019 33065
rect 25130 33028 25136 33040
rect 23400 33000 25136 33028
rect 25130 32988 25136 33000
rect 25188 32988 25194 33040
rect 19518 32960 19524 32972
rect 18288 32932 18552 32960
rect 19306 32932 19524 32960
rect 18288 32920 18294 32932
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 17865 32895 17923 32901
rect 17865 32861 17877 32895
rect 17911 32892 17923 32895
rect 18046 32892 18052 32904
rect 17911 32864 18052 32892
rect 17911 32861 17923 32864
rect 17865 32855 17923 32861
rect 1394 32784 1400 32836
rect 1452 32824 1458 32836
rect 1581 32827 1639 32833
rect 1581 32824 1593 32827
rect 1452 32796 1593 32824
rect 1452 32784 1458 32796
rect 1581 32793 1593 32796
rect 1627 32793 1639 32827
rect 3234 32824 3240 32836
rect 3195 32796 3240 32824
rect 1581 32787 1639 32793
rect 3234 32784 3240 32796
rect 3292 32784 3298 32836
rect 16850 32824 16856 32836
rect 16763 32796 16856 32824
rect 16850 32784 16856 32796
rect 16908 32824 16914 32836
rect 17880 32824 17908 32855
rect 18046 32852 18052 32864
rect 18104 32892 18110 32904
rect 18524 32901 18552 32932
rect 19518 32920 19524 32932
rect 19576 32920 19582 32972
rect 21634 32960 21640 32972
rect 20640 32932 21640 32960
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 18104 32864 18337 32892
rect 18104 32852 18110 32864
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 18325 32855 18383 32861
rect 18509 32895 18567 32901
rect 18509 32861 18521 32895
rect 18555 32861 18567 32895
rect 18509 32855 18567 32861
rect 18598 32852 18604 32904
rect 18656 32892 18662 32904
rect 20640 32901 20668 32932
rect 21634 32920 21640 32932
rect 21692 32920 21698 32972
rect 21910 32920 21916 32972
rect 21968 32960 21974 32972
rect 21968 32932 22416 32960
rect 21968 32920 21974 32932
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18656 32864 19257 32892
rect 18656 32852 18662 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 20625 32895 20683 32901
rect 20625 32861 20637 32895
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 20901 32895 20959 32901
rect 20901 32861 20913 32895
rect 20947 32861 20959 32895
rect 20901 32855 20959 32861
rect 16908 32796 17908 32824
rect 16908 32784 16914 32796
rect 20530 32784 20536 32836
rect 20588 32824 20594 32836
rect 20809 32827 20867 32833
rect 20809 32824 20821 32827
rect 20588 32796 20821 32824
rect 20588 32784 20594 32796
rect 20809 32793 20821 32796
rect 20855 32793 20867 32827
rect 20809 32787 20867 32793
rect 15194 32716 15200 32768
rect 15252 32756 15258 32768
rect 16485 32759 16543 32765
rect 16485 32756 16497 32759
rect 15252 32728 16497 32756
rect 15252 32716 15258 32728
rect 16485 32725 16497 32728
rect 16531 32725 16543 32759
rect 18690 32756 18696 32768
rect 18651 32728 18696 32756
rect 16485 32719 16543 32725
rect 18690 32716 18696 32728
rect 18748 32716 18754 32768
rect 20916 32756 20944 32855
rect 21818 32852 21824 32904
rect 21876 32892 21882 32904
rect 22189 32895 22247 32901
rect 22189 32892 22201 32895
rect 21876 32864 22201 32892
rect 21876 32852 21882 32864
rect 22189 32861 22201 32864
rect 22235 32861 22247 32895
rect 22189 32855 22247 32861
rect 22278 32852 22284 32904
rect 22336 32852 22342 32904
rect 22388 32901 22416 32932
rect 22738 32920 22744 32972
rect 22796 32960 22802 32972
rect 23014 32960 23020 32972
rect 22796 32932 23020 32960
rect 22796 32920 22802 32932
rect 23014 32920 23020 32932
rect 23072 32960 23078 32972
rect 23201 32963 23259 32969
rect 23201 32960 23213 32963
rect 23072 32932 23213 32960
rect 23072 32920 23078 32932
rect 23201 32929 23213 32932
rect 23247 32929 23259 32963
rect 23201 32923 23259 32929
rect 24765 32963 24823 32969
rect 24765 32929 24777 32963
rect 24811 32960 24823 32963
rect 25593 32963 25651 32969
rect 25593 32960 25605 32963
rect 24811 32932 25605 32960
rect 24811 32929 24823 32932
rect 24765 32923 24823 32929
rect 25593 32929 25605 32932
rect 25639 32929 25651 32963
rect 25976 32960 26004 33059
rect 29546 33056 29552 33108
rect 29604 33096 29610 33108
rect 30282 33096 30288 33108
rect 29604 33068 30288 33096
rect 29604 33056 29610 33068
rect 30282 33056 30288 33068
rect 30340 33056 30346 33108
rect 30650 33056 30656 33108
rect 30708 33056 30714 33108
rect 28997 33031 29055 33037
rect 28997 32997 29009 33031
rect 29043 33028 29055 33031
rect 29086 33028 29092 33040
rect 29043 33000 29092 33028
rect 29043 32997 29055 33000
rect 28997 32991 29055 32997
rect 29086 32988 29092 33000
rect 29144 33028 29150 33040
rect 30668 33028 30696 33056
rect 29144 33000 30696 33028
rect 29144 32988 29150 33000
rect 30392 32969 30420 33000
rect 30377 32963 30435 32969
rect 25976 32932 26556 32960
rect 25593 32923 25651 32929
rect 22373 32895 22431 32901
rect 22373 32861 22385 32895
rect 22419 32861 22431 32895
rect 23106 32892 23112 32904
rect 23067 32864 23112 32892
rect 22373 32855 22431 32861
rect 23106 32852 23112 32864
rect 23164 32852 23170 32904
rect 23290 32852 23296 32904
rect 23348 32892 23354 32904
rect 23385 32895 23443 32901
rect 23385 32892 23397 32895
rect 23348 32864 23397 32892
rect 23348 32852 23354 32864
rect 23385 32861 23397 32864
rect 23431 32861 23443 32895
rect 23385 32855 23443 32861
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24673 32895 24731 32901
rect 24673 32892 24685 32895
rect 23900 32864 24685 32892
rect 23900 32852 23906 32864
rect 24673 32861 24685 32864
rect 24719 32861 24731 32895
rect 24673 32855 24731 32861
rect 24949 32895 25007 32901
rect 24949 32861 24961 32895
rect 24995 32892 25007 32895
rect 25038 32892 25044 32904
rect 24995 32864 25044 32892
rect 24995 32861 25007 32864
rect 24949 32855 25007 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 21545 32827 21603 32833
rect 21545 32793 21557 32827
rect 21591 32824 21603 32827
rect 22296 32824 22324 32852
rect 21591 32796 22324 32824
rect 25148 32824 25176 32855
rect 25222 32852 25228 32904
rect 25280 32892 25286 32904
rect 25777 32895 25835 32901
rect 25777 32892 25789 32895
rect 25280 32864 25789 32892
rect 25280 32852 25286 32864
rect 25777 32861 25789 32864
rect 25823 32861 25835 32895
rect 25777 32855 25835 32861
rect 26053 32895 26111 32901
rect 26053 32861 26065 32895
rect 26099 32892 26111 32895
rect 26142 32892 26148 32904
rect 26099 32864 26148 32892
rect 26099 32861 26111 32864
rect 26053 32855 26111 32861
rect 26142 32852 26148 32864
rect 26200 32892 26206 32904
rect 26528 32901 26556 32932
rect 30377 32929 30389 32963
rect 30423 32929 30435 32963
rect 30650 32960 30656 32972
rect 30611 32932 30656 32960
rect 30377 32923 30435 32929
rect 30650 32920 30656 32932
rect 30708 32920 30714 32972
rect 26513 32895 26571 32901
rect 26200 32864 26464 32892
rect 26200 32852 26206 32864
rect 26326 32824 26332 32836
rect 25148 32796 26332 32824
rect 21591 32793 21603 32796
rect 21545 32787 21603 32793
rect 26326 32784 26332 32796
rect 26384 32784 26390 32836
rect 26436 32824 26464 32864
rect 26513 32861 26525 32895
rect 26559 32861 26571 32895
rect 26513 32855 26571 32861
rect 26697 32895 26755 32901
rect 26697 32861 26709 32895
rect 26743 32861 26755 32895
rect 26697 32855 26755 32861
rect 26712 32824 26740 32855
rect 28074 32852 28080 32904
rect 28132 32892 28138 32904
rect 28442 32892 28448 32904
rect 28132 32864 28448 32892
rect 28132 32852 28138 32864
rect 28442 32852 28448 32864
rect 28500 32892 28506 32904
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28500 32864 28641 32892
rect 28500 32852 28506 32864
rect 28629 32861 28641 32864
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 28994 32892 29000 32904
rect 28859 32864 29000 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 28994 32852 29000 32864
rect 29052 32892 29058 32904
rect 29730 32892 29736 32904
rect 29052 32864 29736 32892
rect 29052 32852 29058 32864
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 30285 32895 30343 32901
rect 30285 32861 30297 32895
rect 30331 32861 30343 32895
rect 30285 32855 30343 32861
rect 27982 32824 27988 32836
rect 26436 32796 26740 32824
rect 27943 32796 27988 32824
rect 27982 32784 27988 32796
rect 28040 32784 28046 32836
rect 28169 32827 28227 32833
rect 28169 32793 28181 32827
rect 28215 32824 28227 32827
rect 28718 32824 28724 32836
rect 28215 32796 28724 32824
rect 28215 32793 28227 32796
rect 28169 32787 28227 32793
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 20916 32728 22293 32756
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 23566 32756 23572 32768
rect 23527 32728 23572 32756
rect 22281 32719 22339 32725
rect 23566 32716 23572 32728
rect 23624 32716 23630 32768
rect 25774 32716 25780 32768
rect 25832 32756 25838 32768
rect 26605 32759 26663 32765
rect 26605 32756 26617 32759
rect 25832 32728 26617 32756
rect 25832 32716 25838 32728
rect 26605 32725 26617 32728
rect 26651 32725 26663 32759
rect 26605 32719 26663 32725
rect 27706 32716 27712 32768
rect 27764 32756 27770 32768
rect 28184 32756 28212 32787
rect 28718 32784 28724 32796
rect 28776 32784 28782 32836
rect 30300 32824 30328 32855
rect 30926 32852 30932 32904
rect 30984 32892 30990 32904
rect 31205 32895 31263 32901
rect 31205 32892 31217 32895
rect 30984 32864 31217 32892
rect 30984 32852 30990 32864
rect 31205 32861 31217 32864
rect 31251 32861 31263 32895
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 31205 32855 31263 32861
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 31481 32827 31539 32833
rect 30300 32796 31064 32824
rect 31036 32768 31064 32796
rect 31481 32793 31493 32827
rect 31527 32824 31539 32827
rect 31570 32824 31576 32836
rect 31527 32796 31576 32824
rect 31527 32793 31539 32796
rect 31481 32787 31539 32793
rect 31570 32784 31576 32796
rect 31628 32784 31634 32836
rect 31938 32784 31944 32836
rect 31996 32784 32002 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 47670 32824 47676 32836
rect 46523 32796 47676 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 47670 32784 47676 32796
rect 47728 32784 47734 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 27764 32728 28212 32756
rect 27764 32716 27770 32728
rect 31018 32716 31024 32768
rect 31076 32756 31082 32768
rect 32953 32759 33011 32765
rect 32953 32756 32965 32759
rect 31076 32728 32965 32756
rect 31076 32716 31082 32728
rect 32953 32725 32965 32728
rect 32999 32725 33011 32759
rect 32953 32719 33011 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 16666 32512 16672 32564
rect 16724 32552 16730 32564
rect 17221 32555 17279 32561
rect 17221 32552 17233 32555
rect 16724 32524 17233 32552
rect 16724 32512 16730 32524
rect 17221 32521 17233 32524
rect 17267 32521 17279 32555
rect 17221 32515 17279 32521
rect 18598 32512 18604 32564
rect 18656 32552 18662 32564
rect 19245 32555 19303 32561
rect 19245 32552 19257 32555
rect 18656 32524 19257 32552
rect 18656 32512 18662 32524
rect 19245 32521 19257 32524
rect 19291 32521 19303 32555
rect 19245 32515 19303 32521
rect 24854 32512 24860 32564
rect 24912 32552 24918 32564
rect 25225 32555 25283 32561
rect 25225 32552 25237 32555
rect 24912 32524 25237 32552
rect 24912 32512 24918 32524
rect 25225 32521 25237 32524
rect 25271 32521 25283 32555
rect 27614 32552 27620 32564
rect 27575 32524 27620 32552
rect 25225 32515 25283 32521
rect 27614 32512 27620 32524
rect 27672 32512 27678 32564
rect 31570 32552 31576 32564
rect 31531 32524 31576 32552
rect 31570 32512 31576 32524
rect 31628 32512 31634 32564
rect 47670 32552 47676 32564
rect 47631 32524 47676 32552
rect 47670 32512 47676 32524
rect 47728 32512 47734 32564
rect 2038 32484 2044 32496
rect 1999 32456 2044 32484
rect 2038 32444 2044 32456
rect 2096 32444 2102 32496
rect 16025 32487 16083 32493
rect 16025 32453 16037 32487
rect 16071 32484 16083 32487
rect 16853 32487 16911 32493
rect 16853 32484 16865 32487
rect 16071 32456 16865 32484
rect 16071 32453 16083 32456
rect 16025 32447 16083 32453
rect 16853 32453 16865 32456
rect 16899 32453 16911 32487
rect 16853 32447 16911 32453
rect 16945 32487 17003 32493
rect 16945 32453 16957 32487
rect 16991 32484 17003 32487
rect 16991 32456 17264 32484
rect 16991 32453 17003 32456
rect 16945 32447 17003 32453
rect 15289 32419 15347 32425
rect 15289 32385 15301 32419
rect 15335 32385 15347 32419
rect 15930 32416 15936 32428
rect 15891 32388 15936 32416
rect 15289 32379 15347 32385
rect 1762 32308 1768 32360
rect 1820 32348 1826 32360
rect 1857 32351 1915 32357
rect 1857 32348 1869 32351
rect 1820 32320 1869 32348
rect 1820 32308 1826 32320
rect 1857 32317 1869 32320
rect 1903 32317 1915 32351
rect 3234 32348 3240 32360
rect 3195 32320 3240 32348
rect 1857 32311 1915 32317
rect 3234 32308 3240 32320
rect 3292 32308 3298 32360
rect 15304 32348 15332 32379
rect 15930 32376 15936 32388
rect 15988 32376 15994 32428
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32416 16175 32419
rect 16163 32388 16620 32416
rect 16163 32385 16175 32388
rect 16117 32379 16175 32385
rect 15304 32320 16160 32348
rect 16132 32292 16160 32320
rect 14366 32240 14372 32292
rect 14424 32280 14430 32292
rect 14424 32252 15792 32280
rect 14424 32240 14430 32252
rect 15381 32215 15439 32221
rect 15381 32181 15393 32215
rect 15427 32212 15439 32215
rect 15654 32212 15660 32224
rect 15427 32184 15660 32212
rect 15427 32181 15439 32184
rect 15381 32175 15439 32181
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 15764 32212 15792 32252
rect 16114 32240 16120 32292
rect 16172 32240 16178 32292
rect 16592 32280 16620 32388
rect 16666 32376 16672 32428
rect 16724 32416 16730 32428
rect 17037 32419 17095 32425
rect 16724 32388 16769 32416
rect 16724 32376 16730 32388
rect 17037 32385 17049 32419
rect 17083 32385 17095 32419
rect 17037 32379 17095 32385
rect 16850 32280 16856 32292
rect 16592 32252 16856 32280
rect 16850 32240 16856 32252
rect 16908 32240 16914 32292
rect 17052 32212 17080 32379
rect 17236 32348 17264 32456
rect 17402 32444 17408 32496
rect 17460 32484 17466 32496
rect 23750 32484 23756 32496
rect 17460 32456 23756 32484
rect 17460 32444 17466 32456
rect 23750 32444 23756 32456
rect 23808 32444 23814 32496
rect 25066 32487 25124 32493
rect 25066 32453 25078 32487
rect 25112 32484 25124 32487
rect 25866 32484 25872 32496
rect 25112 32456 25872 32484
rect 25112 32453 25124 32456
rect 25066 32447 25124 32453
rect 25866 32444 25872 32456
rect 25924 32444 25930 32496
rect 26142 32444 26148 32496
rect 26200 32484 26206 32496
rect 27249 32487 27307 32493
rect 26200 32456 27200 32484
rect 26200 32444 26206 32456
rect 17310 32376 17316 32428
rect 17368 32416 17374 32428
rect 17773 32419 17831 32425
rect 17773 32416 17785 32419
rect 17368 32388 17785 32416
rect 17368 32376 17374 32388
rect 17773 32385 17785 32388
rect 17819 32385 17831 32419
rect 18046 32416 18052 32428
rect 18007 32388 18052 32416
rect 17773 32379 17831 32385
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 18230 32416 18236 32428
rect 18191 32388 18236 32416
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 18877 32419 18935 32425
rect 18877 32385 18889 32419
rect 18923 32385 18935 32419
rect 19058 32416 19064 32428
rect 19019 32388 19064 32416
rect 18877 32379 18935 32385
rect 18892 32348 18920 32379
rect 19058 32376 19064 32388
rect 19116 32416 19122 32428
rect 19116 32388 19472 32416
rect 19116 32376 19122 32388
rect 19334 32348 19340 32360
rect 17236 32320 18736 32348
rect 18892 32320 19340 32348
rect 18598 32280 18604 32292
rect 18248 32252 18604 32280
rect 18248 32221 18276 32252
rect 18598 32240 18604 32252
rect 18656 32240 18662 32292
rect 15764 32184 17080 32212
rect 18233 32215 18291 32221
rect 18233 32181 18245 32215
rect 18279 32181 18291 32215
rect 18414 32212 18420 32224
rect 18375 32184 18420 32212
rect 18233 32175 18291 32181
rect 18414 32172 18420 32184
rect 18472 32172 18478 32224
rect 18708 32212 18736 32320
rect 19334 32308 19340 32320
rect 19392 32308 19398 32360
rect 19444 32348 19472 32388
rect 19518 32376 19524 32428
rect 19576 32416 19582 32428
rect 20165 32419 20223 32425
rect 20165 32416 20177 32419
rect 19576 32388 20177 32416
rect 19576 32376 19582 32388
rect 20165 32385 20177 32388
rect 20211 32416 20223 32419
rect 23566 32416 23572 32428
rect 20211 32388 23572 32416
rect 20211 32385 20223 32388
rect 20165 32379 20223 32385
rect 23566 32376 23572 32388
rect 23624 32376 23630 32428
rect 24305 32419 24363 32425
rect 24305 32385 24317 32419
rect 24351 32416 24363 32419
rect 24351 32388 24716 32416
rect 24351 32385 24363 32388
rect 24305 32379 24363 32385
rect 20254 32348 20260 32360
rect 19444 32320 20260 32348
rect 20254 32308 20260 32320
rect 20312 32348 20318 32360
rect 20441 32351 20499 32357
rect 20441 32348 20453 32351
rect 20312 32320 20453 32348
rect 20312 32308 20318 32320
rect 20441 32317 20453 32320
rect 20487 32317 20499 32351
rect 20441 32311 20499 32317
rect 23474 32308 23480 32360
rect 23532 32348 23538 32360
rect 24320 32348 24348 32379
rect 23532 32320 24348 32348
rect 24581 32351 24639 32357
rect 23532 32308 23538 32320
rect 24581 32317 24593 32351
rect 24627 32317 24639 32351
rect 24688 32348 24716 32388
rect 24762 32376 24768 32428
rect 24820 32416 24826 32428
rect 24949 32419 25007 32425
rect 24949 32416 24961 32419
rect 24820 32388 24961 32416
rect 24820 32376 24826 32388
rect 24949 32385 24961 32388
rect 24995 32385 25007 32419
rect 25774 32416 25780 32428
rect 25735 32388 25780 32416
rect 24949 32379 25007 32385
rect 25774 32376 25780 32388
rect 25832 32376 25838 32428
rect 26970 32416 26976 32428
rect 26931 32388 26976 32416
rect 26970 32376 26976 32388
rect 27028 32376 27034 32428
rect 27066 32419 27124 32425
rect 27066 32385 27078 32419
rect 27112 32385 27124 32419
rect 27172 32416 27200 32456
rect 27249 32453 27261 32487
rect 27295 32484 27307 32487
rect 28258 32484 28264 32496
rect 27295 32456 28264 32484
rect 27295 32453 27307 32456
rect 27249 32447 27307 32453
rect 28258 32444 28264 32456
rect 28316 32444 28322 32496
rect 30558 32444 30564 32496
rect 30616 32484 30622 32496
rect 47486 32484 47492 32496
rect 30616 32456 31340 32484
rect 30616 32444 30622 32456
rect 31312 32428 31340 32456
rect 35866 32456 47492 32484
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 27172 32388 27353 32416
rect 27066 32379 27124 32385
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27479 32419 27537 32425
rect 27479 32385 27491 32419
rect 27525 32416 27537 32419
rect 27614 32416 27620 32428
rect 27525 32388 27620 32416
rect 27525 32385 27537 32388
rect 27479 32379 27537 32385
rect 24857 32351 24915 32357
rect 24857 32348 24869 32351
rect 24688 32320 24869 32348
rect 24581 32311 24639 32317
rect 24857 32317 24869 32320
rect 24903 32348 24915 32351
rect 26237 32351 26295 32357
rect 24903 32320 26096 32348
rect 24903 32317 24915 32320
rect 24857 32311 24915 32317
rect 24596 32280 24624 32311
rect 25038 32280 25044 32292
rect 24596 32252 25044 32280
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 26068 32280 26096 32320
rect 26237 32317 26249 32351
rect 26283 32348 26295 32351
rect 27080 32348 27108 32379
rect 27614 32376 27620 32388
rect 27672 32376 27678 32428
rect 28626 32416 28632 32428
rect 28587 32388 28632 32416
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 28813 32419 28871 32425
rect 28813 32385 28825 32419
rect 28859 32416 28871 32419
rect 29086 32416 29092 32428
rect 28859 32388 29092 32416
rect 28859 32385 28871 32388
rect 28813 32379 28871 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 30834 32376 30840 32428
rect 30892 32416 30898 32428
rect 30929 32419 30987 32425
rect 30929 32416 30941 32419
rect 30892 32388 30941 32416
rect 30892 32376 30898 32388
rect 30929 32385 30941 32388
rect 30975 32385 30987 32419
rect 30929 32379 30987 32385
rect 31018 32376 31024 32428
rect 31076 32416 31082 32428
rect 31205 32419 31263 32425
rect 31076 32388 31121 32416
rect 31076 32376 31082 32388
rect 31205 32385 31217 32419
rect 31251 32385 31263 32419
rect 31205 32379 31263 32385
rect 26283 32320 27108 32348
rect 26283 32317 26295 32320
rect 26237 32311 26295 32317
rect 30466 32308 30472 32360
rect 30524 32348 30530 32360
rect 31220 32348 31248 32379
rect 31294 32376 31300 32428
rect 31352 32416 31358 32428
rect 31435 32419 31493 32425
rect 31352 32388 31397 32416
rect 31352 32376 31358 32388
rect 31435 32385 31447 32419
rect 31481 32416 31493 32419
rect 35866 32416 35894 32456
rect 47486 32444 47492 32456
rect 47544 32444 47550 32496
rect 31481 32388 35894 32416
rect 31481 32385 31493 32388
rect 31435 32379 31493 32385
rect 46290 32376 46296 32428
rect 46348 32416 46354 32428
rect 47029 32419 47087 32425
rect 47029 32416 47041 32419
rect 46348 32388 47041 32416
rect 46348 32376 46354 32388
rect 47029 32385 47041 32388
rect 47075 32385 47087 32419
rect 47029 32379 47087 32385
rect 47581 32419 47639 32425
rect 47581 32385 47593 32419
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 44174 32348 44180 32360
rect 30524 32320 31248 32348
rect 35866 32320 44180 32348
rect 30524 32308 30530 32320
rect 35866 32280 35894 32320
rect 44174 32308 44180 32320
rect 44232 32308 44238 32360
rect 46658 32308 46664 32360
rect 46716 32348 46722 32360
rect 47596 32348 47624 32379
rect 46716 32320 47624 32348
rect 46716 32308 46722 32320
rect 26068 32252 35894 32280
rect 20162 32212 20168 32224
rect 18708 32184 20168 32212
rect 20162 32172 20168 32184
rect 20220 32172 20226 32224
rect 25866 32212 25872 32224
rect 25827 32184 25872 32212
rect 25866 32172 25872 32184
rect 25924 32172 25930 32224
rect 28534 32172 28540 32224
rect 28592 32212 28598 32224
rect 28721 32215 28779 32221
rect 28721 32212 28733 32215
rect 28592 32184 28733 32212
rect 28592 32172 28598 32184
rect 28721 32181 28733 32184
rect 28767 32181 28779 32215
rect 28721 32175 28779 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1394 32008 1400 32020
rect 1355 31980 1400 32008
rect 1394 31968 1400 31980
rect 1452 31968 1458 32020
rect 17221 32011 17279 32017
rect 17221 31977 17233 32011
rect 17267 32008 17279 32011
rect 17770 32008 17776 32020
rect 17267 31980 17776 32008
rect 17267 31977 17279 31980
rect 17221 31971 17279 31977
rect 17770 31968 17776 31980
rect 17828 31968 17834 32020
rect 18417 32011 18475 32017
rect 18417 32008 18429 32011
rect 17880 31980 18429 32008
rect 16669 31943 16727 31949
rect 16669 31909 16681 31943
rect 16715 31940 16727 31943
rect 16850 31940 16856 31952
rect 16715 31912 16856 31940
rect 16715 31909 16727 31912
rect 16669 31903 16727 31909
rect 16850 31900 16856 31912
rect 16908 31900 16914 31952
rect 14734 31832 14740 31884
rect 14792 31872 14798 31884
rect 14921 31875 14979 31881
rect 14921 31872 14933 31875
rect 14792 31844 14933 31872
rect 14792 31832 14798 31844
rect 14921 31841 14933 31844
rect 14967 31841 14979 31875
rect 15194 31872 15200 31884
rect 15155 31844 15200 31872
rect 14921 31835 14979 31841
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 15930 31832 15936 31884
rect 15988 31872 15994 31884
rect 17880 31872 17908 31980
rect 18417 31977 18429 31980
rect 18463 31977 18475 32011
rect 18417 31971 18475 31977
rect 18509 32011 18567 32017
rect 18509 31977 18521 32011
rect 18555 32008 18567 32011
rect 19334 32008 19340 32020
rect 18555 31980 19340 32008
rect 18555 31977 18567 31980
rect 18509 31971 18567 31977
rect 17954 31900 17960 31952
rect 18012 31940 18018 31952
rect 18432 31940 18460 31971
rect 19334 31968 19340 31980
rect 19392 32008 19398 32020
rect 19521 32011 19579 32017
rect 19521 32008 19533 32011
rect 19392 31980 19533 32008
rect 19392 31968 19398 31980
rect 19521 31977 19533 31980
rect 19567 32008 19579 32011
rect 20346 32008 20352 32020
rect 19567 31980 20352 32008
rect 19567 31977 19579 31980
rect 19521 31971 19579 31977
rect 20346 31968 20352 31980
rect 20404 31968 20410 32020
rect 20714 31968 20720 32020
rect 20772 32008 20778 32020
rect 21269 32011 21327 32017
rect 21269 32008 21281 32011
rect 20772 31980 21281 32008
rect 20772 31968 20778 31980
rect 21269 31977 21281 31980
rect 21315 31977 21327 32011
rect 21269 31971 21327 31977
rect 21726 31968 21732 32020
rect 21784 32008 21790 32020
rect 28626 32008 28632 32020
rect 21784 31980 23704 32008
rect 28587 31980 28632 32008
rect 21784 31968 21790 31980
rect 18690 31940 18696 31952
rect 18012 31912 18057 31940
rect 18432 31912 18696 31940
rect 18012 31900 18018 31912
rect 18690 31900 18696 31912
rect 18748 31940 18754 31952
rect 18748 31912 19380 31940
rect 18748 31900 18754 31912
rect 19352 31881 19380 31912
rect 19978 31900 19984 31952
rect 20036 31940 20042 31952
rect 20254 31940 20260 31952
rect 20036 31912 20260 31940
rect 20036 31900 20042 31912
rect 20254 31900 20260 31912
rect 20312 31900 20318 31952
rect 20990 31900 20996 31952
rect 21048 31940 21054 31952
rect 22005 31943 22063 31949
rect 22005 31940 22017 31943
rect 21048 31912 22017 31940
rect 21048 31900 21054 31912
rect 22005 31909 22017 31912
rect 22051 31909 22063 31943
rect 23676 31940 23704 31980
rect 28626 31968 28632 31980
rect 28684 31968 28690 32020
rect 30834 32008 30840 32020
rect 30795 31980 30840 32008
rect 30834 31968 30840 31980
rect 30892 31968 30898 32020
rect 23676 31912 27476 31940
rect 22005 31903 22063 31909
rect 15988 31844 17172 31872
rect 15988 31832 15994 31844
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 2038 31764 2044 31816
rect 2096 31804 2102 31816
rect 2317 31807 2375 31813
rect 2317 31804 2329 31807
rect 2096 31776 2329 31804
rect 2096 31764 2102 31776
rect 2317 31773 2329 31776
rect 2363 31773 2375 31807
rect 2317 31767 2375 31773
rect 2777 31807 2835 31813
rect 2777 31773 2789 31807
rect 2823 31804 2835 31807
rect 2958 31804 2964 31816
rect 2823 31776 2964 31804
rect 2823 31773 2835 31776
rect 2777 31767 2835 31773
rect 2958 31764 2964 31776
rect 3016 31764 3022 31816
rect 15654 31696 15660 31748
rect 15712 31696 15718 31748
rect 17144 31736 17172 31844
rect 17236 31844 17908 31872
rect 18325 31875 18383 31881
rect 17236 31813 17264 31844
rect 18325 31841 18337 31875
rect 18371 31872 18383 31875
rect 19337 31875 19395 31881
rect 18371 31844 19288 31872
rect 18371 31841 18383 31844
rect 18325 31835 18383 31841
rect 17221 31807 17279 31813
rect 17221 31773 17233 31807
rect 17267 31773 17279 31807
rect 17405 31807 17463 31813
rect 17405 31804 17417 31807
rect 17221 31767 17279 31773
rect 17328 31776 17417 31804
rect 17328 31736 17356 31776
rect 17405 31773 17417 31776
rect 17451 31804 17463 31807
rect 17451 31776 17908 31804
rect 17451 31773 17463 31776
rect 17405 31767 17463 31773
rect 17144 31708 17356 31736
rect 17880 31736 17908 31776
rect 18046 31764 18052 31816
rect 18104 31804 18110 31816
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 18104 31776 18245 31804
rect 18104 31764 18110 31776
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31804 18751 31807
rect 19058 31804 19064 31816
rect 18739 31776 19064 31804
rect 18739 31773 18751 31776
rect 18693 31767 18751 31773
rect 19058 31764 19064 31776
rect 19116 31764 19122 31816
rect 19260 31813 19288 31844
rect 19337 31841 19349 31875
rect 19383 31841 19395 31875
rect 19337 31835 19395 31841
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 21726 31872 21732 31884
rect 20956 31844 21732 31872
rect 20956 31832 20962 31844
rect 21726 31832 21732 31844
rect 21784 31832 21790 31884
rect 23385 31875 23443 31881
rect 23385 31872 23397 31875
rect 22066 31844 23397 31872
rect 19245 31807 19303 31813
rect 19245 31773 19257 31807
rect 19291 31804 19303 31807
rect 19518 31804 19524 31816
rect 19291 31776 19380 31804
rect 19479 31776 19524 31804
rect 19291 31773 19303 31776
rect 19245 31767 19303 31773
rect 19352 31748 19380 31776
rect 19518 31764 19524 31776
rect 19576 31764 19582 31816
rect 20622 31804 20628 31816
rect 20583 31776 20628 31804
rect 20622 31764 20628 31776
rect 20680 31764 20686 31816
rect 20806 31813 20812 31816
rect 20773 31807 20812 31813
rect 20773 31773 20785 31807
rect 20773 31767 20812 31773
rect 20806 31764 20812 31767
rect 20864 31764 20870 31816
rect 21082 31764 21088 31816
rect 21140 31813 21146 31816
rect 21140 31804 21148 31813
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21140 31776 21185 31804
rect 21284 31776 21833 31804
rect 21140 31767 21148 31776
rect 21140 31764 21146 31767
rect 18322 31736 18328 31748
rect 17880 31708 18328 31736
rect 18322 31696 18328 31708
rect 18380 31696 18386 31748
rect 19334 31696 19340 31748
rect 19392 31696 19398 31748
rect 20898 31736 20904 31748
rect 20859 31708 20904 31736
rect 20898 31696 20904 31708
rect 20956 31696 20962 31748
rect 20990 31696 20996 31748
rect 21048 31736 21054 31748
rect 21048 31708 21093 31736
rect 21048 31696 21054 31708
rect 2866 31668 2872 31680
rect 2827 31640 2872 31668
rect 2866 31628 2872 31640
rect 2924 31628 2930 31680
rect 11698 31628 11704 31680
rect 11756 31668 11762 31680
rect 16574 31668 16580 31680
rect 11756 31640 16580 31668
rect 11756 31628 11762 31640
rect 16574 31628 16580 31640
rect 16632 31628 16638 31680
rect 19705 31671 19763 31677
rect 19705 31637 19717 31671
rect 19751 31668 19763 31671
rect 19978 31668 19984 31680
rect 19751 31640 19984 31668
rect 19751 31637 19763 31640
rect 19705 31631 19763 31637
rect 19978 31628 19984 31640
rect 20036 31628 20042 31680
rect 20162 31628 20168 31680
rect 20220 31668 20226 31680
rect 21284 31668 21312 31776
rect 21821 31773 21833 31776
rect 21867 31804 21879 31807
rect 22066 31804 22094 31844
rect 23385 31841 23397 31844
rect 23431 31872 23443 31875
rect 23842 31872 23848 31884
rect 23431 31844 23848 31872
rect 23431 31841 23443 31844
rect 23385 31835 23443 31841
rect 23842 31832 23848 31844
rect 23900 31832 23906 31884
rect 27448 31872 27476 31912
rect 27522 31900 27528 31952
rect 27580 31940 27586 31952
rect 30926 31940 30932 31952
rect 27580 31912 30932 31940
rect 27580 31900 27586 31912
rect 30926 31900 30932 31912
rect 30984 31900 30990 31952
rect 27614 31872 27620 31884
rect 27448 31844 27620 31872
rect 27614 31832 27620 31844
rect 27672 31872 27678 31884
rect 30466 31872 30472 31884
rect 27672 31844 30472 31872
rect 27672 31832 27678 31844
rect 30466 31832 30472 31844
rect 30524 31832 30530 31884
rect 47302 31872 47308 31884
rect 47263 31844 47308 31872
rect 47302 31832 47308 31844
rect 47360 31832 47366 31884
rect 47486 31832 47492 31884
rect 47544 31872 47550 31884
rect 47581 31875 47639 31881
rect 47581 31872 47593 31875
rect 47544 31844 47593 31872
rect 47544 31832 47550 31844
rect 47581 31841 47593 31844
rect 47627 31841 47639 31875
rect 47581 31835 47639 31841
rect 21867 31776 22094 31804
rect 21867 31773 21879 31776
rect 21821 31767 21879 31773
rect 22554 31764 22560 31816
rect 22612 31804 22618 31816
rect 23201 31807 23259 31813
rect 23201 31804 23213 31807
rect 22612 31776 23213 31804
rect 22612 31764 22618 31776
rect 23201 31773 23213 31776
rect 23247 31773 23259 31807
rect 23201 31767 23259 31773
rect 24762 31764 24768 31816
rect 24820 31804 24826 31816
rect 24857 31807 24915 31813
rect 24857 31804 24869 31807
rect 24820 31776 24869 31804
rect 24820 31764 24826 31776
rect 24857 31773 24869 31776
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 25225 31807 25283 31813
rect 25225 31773 25237 31807
rect 25271 31804 25283 31807
rect 25314 31804 25320 31816
rect 25271 31776 25320 31804
rect 25271 31773 25283 31776
rect 25225 31767 25283 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 27154 31804 27160 31816
rect 27115 31776 27160 31804
rect 27154 31764 27160 31776
rect 27212 31764 27218 31816
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28442 31804 28448 31816
rect 28224 31776 28448 31804
rect 28224 31764 28230 31776
rect 28442 31764 28448 31776
rect 28500 31804 28506 31816
rect 28537 31807 28595 31813
rect 28537 31804 28549 31807
rect 28500 31776 28549 31804
rect 28500 31764 28506 31776
rect 28537 31773 28549 31776
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 28721 31807 28779 31813
rect 28721 31773 28733 31807
rect 28767 31804 28779 31807
rect 28994 31804 29000 31816
rect 28767 31776 29000 31804
rect 28767 31773 28779 31776
rect 28721 31767 28779 31773
rect 28994 31764 29000 31776
rect 29052 31764 29058 31816
rect 30650 31764 30656 31816
rect 30708 31804 30714 31816
rect 30837 31807 30895 31813
rect 30837 31804 30849 31807
rect 30708 31776 30849 31804
rect 30708 31764 30714 31776
rect 30837 31773 30849 31776
rect 30883 31773 30895 31807
rect 30837 31767 30895 31773
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 31076 31776 31121 31804
rect 31076 31764 31082 31776
rect 23750 31696 23756 31748
rect 23808 31736 23814 31748
rect 27706 31736 27712 31748
rect 23808 31708 27712 31736
rect 23808 31696 23814 31708
rect 27706 31696 27712 31708
rect 27764 31736 27770 31748
rect 27893 31739 27951 31745
rect 27893 31736 27905 31739
rect 27764 31708 27905 31736
rect 27764 31696 27770 31708
rect 27893 31705 27905 31708
rect 27939 31705 27951 31739
rect 27893 31699 27951 31705
rect 28077 31739 28135 31745
rect 28077 31705 28089 31739
rect 28123 31736 28135 31739
rect 28258 31736 28264 31748
rect 28123 31708 28264 31736
rect 28123 31705 28135 31708
rect 28077 31699 28135 31705
rect 28258 31696 28264 31708
rect 28316 31696 28322 31748
rect 20220 31640 21312 31668
rect 20220 31628 20226 31640
rect 26234 31628 26240 31680
rect 26292 31668 26298 31680
rect 27249 31671 27307 31677
rect 27249 31668 27261 31671
rect 26292 31640 27261 31668
rect 26292 31628 26298 31640
rect 27249 31637 27261 31640
rect 27295 31668 27307 31671
rect 27522 31668 27528 31680
rect 27295 31640 27528 31668
rect 27295 31637 27307 31640
rect 27249 31631 27307 31637
rect 27522 31628 27528 31640
rect 27580 31628 27586 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 16942 31424 16948 31476
rect 17000 31464 17006 31476
rect 17865 31467 17923 31473
rect 17865 31464 17877 31467
rect 17000 31436 17877 31464
rect 17000 31424 17006 31436
rect 17865 31433 17877 31436
rect 17911 31433 17923 31467
rect 22278 31464 22284 31476
rect 22239 31436 22284 31464
rect 17865 31427 17923 31433
rect 22278 31424 22284 31436
rect 22336 31424 22342 31476
rect 23198 31424 23204 31476
rect 23256 31464 23262 31476
rect 23256 31436 26464 31464
rect 23256 31424 23262 31436
rect 2225 31399 2283 31405
rect 2225 31365 2237 31399
rect 2271 31396 2283 31399
rect 2866 31396 2872 31408
rect 2271 31368 2872 31396
rect 2271 31365 2283 31368
rect 2225 31359 2283 31365
rect 2866 31356 2872 31368
rect 2924 31356 2930 31408
rect 16574 31356 16580 31408
rect 16632 31396 16638 31408
rect 22189 31399 22247 31405
rect 16632 31368 20760 31396
rect 16632 31356 16638 31368
rect 2038 31328 2044 31340
rect 1999 31300 2044 31328
rect 2038 31288 2044 31300
rect 2096 31288 2102 31340
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31297 18107 31331
rect 18230 31328 18236 31340
rect 18191 31300 18236 31328
rect 18049 31291 18107 31297
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 2832 31232 2877 31260
rect 2832 31220 2838 31232
rect 18064 31192 18092 31291
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 18322 31288 18328 31340
rect 18380 31328 18386 31340
rect 20346 31328 20352 31340
rect 18380 31300 18425 31328
rect 20307 31300 20352 31328
rect 18380 31288 18386 31300
rect 20346 31288 20352 31300
rect 20404 31288 20410 31340
rect 20530 31328 20536 31340
rect 20491 31300 20536 31328
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 20732 31337 20760 31368
rect 22189 31365 22201 31399
rect 22235 31396 22247 31399
rect 26326 31396 26332 31408
rect 22235 31368 26332 31396
rect 22235 31365 22247 31368
rect 22189 31359 22247 31365
rect 26326 31356 26332 31368
rect 26384 31356 26390 31408
rect 26436 31396 26464 31436
rect 28166 31424 28172 31476
rect 28224 31424 28230 31476
rect 28184 31396 28212 31424
rect 26436 31368 28212 31396
rect 20625 31331 20683 31337
rect 20625 31297 20637 31331
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20717 31331 20775 31337
rect 20717 31297 20729 31331
rect 20763 31297 20775 31331
rect 22830 31328 22836 31340
rect 22791 31300 22836 31328
rect 20717 31291 20775 31297
rect 20162 31220 20168 31272
rect 20220 31260 20226 31272
rect 20640 31260 20668 31291
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23106 31328 23112 31340
rect 23063 31300 23112 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23106 31288 23112 31300
rect 23164 31288 23170 31340
rect 23198 31288 23204 31340
rect 23256 31328 23262 31340
rect 23937 31331 23995 31337
rect 23256 31300 23301 31328
rect 23256 31288 23262 31300
rect 23937 31297 23949 31331
rect 23983 31328 23995 31331
rect 24762 31328 24768 31340
rect 23983 31300 24768 31328
rect 23983 31297 23995 31300
rect 23937 31291 23995 31297
rect 24762 31288 24768 31300
rect 24820 31288 24826 31340
rect 25130 31328 25136 31340
rect 25091 31300 25136 31328
rect 25130 31288 25136 31300
rect 25188 31288 25194 31340
rect 26436 31337 26464 31368
rect 28442 31356 28448 31408
rect 28500 31356 28506 31408
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31297 26295 31331
rect 26237 31291 26295 31297
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31297 26479 31331
rect 27522 31328 27528 31340
rect 27483 31300 27528 31328
rect 26421 31291 26479 31297
rect 20220 31232 20668 31260
rect 23661 31263 23719 31269
rect 20220 31220 20226 31232
rect 23661 31229 23673 31263
rect 23707 31229 23719 31263
rect 23661 31223 23719 31229
rect 20530 31192 20536 31204
rect 18064 31164 20536 31192
rect 20530 31152 20536 31164
rect 20588 31152 20594 31204
rect 23566 31192 23572 31204
rect 20640 31164 23572 31192
rect 14274 31084 14280 31136
rect 14332 31124 14338 31136
rect 19978 31124 19984 31136
rect 14332 31096 19984 31124
rect 14332 31084 14338 31096
rect 19978 31084 19984 31096
rect 20036 31124 20042 31136
rect 20640 31124 20668 31164
rect 23566 31152 23572 31164
rect 23624 31192 23630 31204
rect 23676 31192 23704 31223
rect 23624 31164 23704 31192
rect 26252 31192 26280 31291
rect 27522 31288 27528 31300
rect 27580 31288 27586 31340
rect 30558 31288 30564 31340
rect 30616 31328 30622 31340
rect 30837 31331 30895 31337
rect 30837 31328 30849 31331
rect 30616 31300 30849 31328
rect 30616 31288 30622 31300
rect 30837 31297 30849 31300
rect 30883 31297 30895 31331
rect 30837 31291 30895 31297
rect 31021 31331 31079 31337
rect 31021 31297 31033 31331
rect 31067 31297 31079 31331
rect 31021 31291 31079 31297
rect 27798 31260 27804 31272
rect 27759 31232 27804 31260
rect 27798 31220 27804 31232
rect 27856 31220 27862 31272
rect 31036 31260 31064 31291
rect 31110 31288 31116 31340
rect 31168 31328 31174 31340
rect 31168 31300 31213 31328
rect 31168 31288 31174 31300
rect 28828 31232 31064 31260
rect 26510 31192 26516 31204
rect 26252 31164 26516 31192
rect 23624 31152 23630 31164
rect 26510 31152 26516 31164
rect 26568 31152 26574 31204
rect 20898 31124 20904 31136
rect 20036 31096 20668 31124
rect 20859 31096 20904 31124
rect 20036 31084 20042 31096
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 24394 31084 24400 31136
rect 24452 31124 24458 31136
rect 25225 31127 25283 31133
rect 25225 31124 25237 31127
rect 24452 31096 25237 31124
rect 24452 31084 24458 31096
rect 25225 31093 25237 31096
rect 25271 31093 25283 31127
rect 25225 31087 25283 31093
rect 25682 31084 25688 31136
rect 25740 31124 25746 31136
rect 26237 31127 26295 31133
rect 26237 31124 26249 31127
rect 25740 31096 26249 31124
rect 25740 31084 25746 31096
rect 26237 31093 26249 31096
rect 26283 31093 26295 31127
rect 26237 31087 26295 31093
rect 27338 31084 27344 31136
rect 27396 31124 27402 31136
rect 28828 31124 28856 31232
rect 27396 31096 28856 31124
rect 27396 31084 27402 31096
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 29270 31124 29276 31136
rect 29052 31096 29276 31124
rect 29052 31084 29058 31096
rect 29270 31084 29276 31096
rect 29328 31084 29334 31136
rect 30653 31127 30711 31133
rect 30653 31093 30665 31127
rect 30699 31124 30711 31127
rect 31294 31124 31300 31136
rect 30699 31096 31300 31124
rect 30699 31093 30711 31096
rect 30653 31087 30711 31093
rect 31294 31084 31300 31096
rect 31352 31084 31358 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 19334 30880 19340 30932
rect 19392 30920 19398 30932
rect 19613 30923 19671 30929
rect 19613 30920 19625 30923
rect 19392 30892 19625 30920
rect 19392 30880 19398 30892
rect 19613 30889 19625 30892
rect 19659 30889 19671 30923
rect 19613 30883 19671 30889
rect 23569 30923 23627 30929
rect 23569 30889 23581 30923
rect 23615 30889 23627 30923
rect 23750 30920 23756 30932
rect 23711 30892 23756 30920
rect 23569 30883 23627 30889
rect 23584 30852 23612 30883
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 26053 30923 26111 30929
rect 26053 30889 26065 30923
rect 26099 30920 26111 30923
rect 26326 30920 26332 30932
rect 26099 30892 26332 30920
rect 26099 30889 26111 30892
rect 26053 30883 26111 30889
rect 26326 30880 26332 30892
rect 26384 30880 26390 30932
rect 26970 30880 26976 30932
rect 27028 30920 27034 30932
rect 27525 30923 27583 30929
rect 27525 30920 27537 30923
rect 27028 30892 27537 30920
rect 27028 30880 27034 30892
rect 27525 30889 27537 30892
rect 27571 30889 27583 30923
rect 27525 30883 27583 30889
rect 27798 30880 27804 30932
rect 27856 30920 27862 30932
rect 28997 30923 29055 30929
rect 28997 30920 29009 30923
rect 27856 30892 29009 30920
rect 27856 30880 27862 30892
rect 28997 30889 29009 30892
rect 29043 30889 29055 30923
rect 30558 30920 30564 30932
rect 30519 30892 30564 30920
rect 28997 30883 29055 30889
rect 30558 30880 30564 30892
rect 30616 30880 30622 30932
rect 24394 30852 24400 30864
rect 23584 30824 24400 30852
rect 17770 30784 17776 30796
rect 17696 30756 17776 30784
rect 16114 30716 16120 30728
rect 16075 30688 16120 30716
rect 16114 30676 16120 30688
rect 16172 30676 16178 30728
rect 17586 30716 17592 30728
rect 17547 30688 17592 30716
rect 17586 30676 17592 30688
rect 17644 30676 17650 30728
rect 17696 30725 17724 30756
rect 17770 30744 17776 30756
rect 17828 30744 17834 30796
rect 21177 30787 21235 30793
rect 21177 30753 21189 30787
rect 21223 30784 21235 30787
rect 23198 30784 23204 30796
rect 21223 30756 23204 30784
rect 21223 30753 21235 30756
rect 21177 30747 21235 30753
rect 23198 30744 23204 30756
rect 23256 30744 23262 30796
rect 17681 30719 17739 30725
rect 17681 30685 17693 30719
rect 17727 30685 17739 30719
rect 17681 30679 17739 30685
rect 18049 30719 18107 30725
rect 18049 30685 18061 30719
rect 18095 30716 18107 30719
rect 18138 30716 18144 30728
rect 18095 30688 18144 30716
rect 18095 30685 18107 30688
rect 18049 30679 18107 30685
rect 18138 30676 18144 30688
rect 18196 30716 18202 30728
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18196 30688 19257 30716
rect 18196 30676 18202 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 20346 30676 20352 30728
rect 20404 30716 20410 30728
rect 20714 30716 20720 30728
rect 20404 30688 20720 30716
rect 20404 30676 20410 30688
rect 20714 30676 20720 30688
rect 20772 30716 20778 30728
rect 21085 30719 21143 30725
rect 21085 30716 21097 30719
rect 20772 30688 21097 30716
rect 20772 30676 20778 30688
rect 21085 30685 21097 30688
rect 21131 30685 21143 30719
rect 21085 30679 21143 30685
rect 22649 30719 22707 30725
rect 22649 30685 22661 30719
rect 22695 30716 22707 30719
rect 23584 30716 23612 30824
rect 24394 30812 24400 30824
rect 24452 30812 24458 30864
rect 28166 30812 28172 30864
rect 28224 30852 28230 30864
rect 28224 30824 30604 30852
rect 28224 30812 28230 30824
rect 30466 30784 30472 30796
rect 28920 30756 30472 30784
rect 22695 30688 23612 30716
rect 22695 30685 22707 30688
rect 22649 30679 22707 30685
rect 26694 30676 26700 30728
rect 26752 30716 26758 30728
rect 27157 30719 27215 30725
rect 27157 30716 27169 30719
rect 26752 30688 27169 30716
rect 26752 30676 26758 30688
rect 27157 30685 27169 30688
rect 27203 30685 27215 30719
rect 27157 30679 27215 30685
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30685 27399 30719
rect 28350 30716 28356 30728
rect 28311 30688 28356 30716
rect 27341 30679 27399 30685
rect 17034 30608 17040 30660
rect 17092 30648 17098 30660
rect 17770 30648 17776 30660
rect 17092 30620 17776 30648
rect 17092 30608 17098 30620
rect 17770 30608 17776 30620
rect 17828 30608 17834 30660
rect 17911 30651 17969 30657
rect 17911 30617 17923 30651
rect 17957 30648 17969 30651
rect 18414 30648 18420 30660
rect 17957 30620 18420 30648
rect 17957 30617 17969 30620
rect 17911 30611 17969 30617
rect 18414 30608 18420 30620
rect 18472 30608 18478 30660
rect 19429 30651 19487 30657
rect 19429 30617 19441 30651
rect 19475 30617 19487 30651
rect 19429 30611 19487 30617
rect 16209 30583 16267 30589
rect 16209 30549 16221 30583
rect 16255 30580 16267 30583
rect 16574 30580 16580 30592
rect 16255 30552 16580 30580
rect 16255 30549 16267 30552
rect 16209 30543 16267 30549
rect 16574 30540 16580 30552
rect 16632 30540 16638 30592
rect 17402 30580 17408 30592
rect 17363 30552 17408 30580
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 17788 30580 17816 30608
rect 19444 30580 19472 30611
rect 20806 30608 20812 30660
rect 20864 30648 20870 30660
rect 23382 30648 23388 30660
rect 20864 30620 22876 30648
rect 23343 30620 23388 30648
rect 20864 30608 20870 30620
rect 17788 30552 19472 30580
rect 21174 30540 21180 30592
rect 21232 30580 21238 30592
rect 22848 30589 22876 30620
rect 23382 30608 23388 30620
rect 23440 30608 23446 30660
rect 23566 30648 23572 30660
rect 23527 30620 23572 30648
rect 23566 30608 23572 30620
rect 23624 30608 23630 30660
rect 24762 30648 24768 30660
rect 24723 30620 24768 30648
rect 24762 30608 24768 30620
rect 24820 30608 24826 30660
rect 26786 30608 26792 30660
rect 26844 30648 26850 30660
rect 27356 30648 27384 30679
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 28534 30725 28540 30728
rect 28501 30719 28540 30725
rect 28501 30685 28513 30719
rect 28501 30679 28540 30685
rect 28534 30676 28540 30679
rect 28592 30676 28598 30728
rect 28818 30719 28876 30725
rect 28818 30685 28830 30719
rect 28864 30716 28876 30719
rect 28920 30716 28948 30756
rect 30466 30744 30472 30756
rect 30524 30744 30530 30796
rect 30006 30716 30012 30728
rect 28864 30688 28948 30716
rect 29967 30688 30012 30716
rect 28864 30685 28876 30688
rect 28818 30679 28876 30685
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 30377 30719 30435 30725
rect 30377 30685 30389 30719
rect 30423 30716 30435 30719
rect 30576 30716 30604 30824
rect 30926 30744 30932 30796
rect 30984 30784 30990 30796
rect 31021 30787 31079 30793
rect 31021 30784 31033 30787
rect 30984 30756 31033 30784
rect 30984 30744 30990 30756
rect 31021 30753 31033 30756
rect 31067 30753 31079 30787
rect 31294 30784 31300 30796
rect 31255 30756 31300 30784
rect 31021 30747 31079 30753
rect 31294 30744 31300 30756
rect 31352 30744 31358 30796
rect 30423 30688 30604 30716
rect 30423 30685 30435 30688
rect 30377 30679 30435 30685
rect 26844 30620 27384 30648
rect 26844 30608 26850 30620
rect 28258 30608 28264 30660
rect 28316 30648 28322 30660
rect 28629 30651 28687 30657
rect 28629 30648 28641 30651
rect 28316 30620 28641 30648
rect 28316 30608 28322 30620
rect 28629 30617 28641 30620
rect 28675 30617 28687 30651
rect 28629 30611 28687 30617
rect 28721 30651 28779 30657
rect 28721 30617 28733 30651
rect 28767 30648 28779 30651
rect 29270 30648 29276 30660
rect 28767 30620 29276 30648
rect 28767 30617 28779 30620
rect 28721 30611 28779 30617
rect 21453 30583 21511 30589
rect 21453 30580 21465 30583
rect 21232 30552 21465 30580
rect 21232 30540 21238 30552
rect 21453 30549 21465 30552
rect 21499 30549 21511 30583
rect 21453 30543 21511 30549
rect 22833 30583 22891 30589
rect 22833 30549 22845 30583
rect 22879 30580 22891 30583
rect 27246 30580 27252 30592
rect 22879 30552 27252 30580
rect 22879 30549 22891 30552
rect 22833 30543 22891 30549
rect 27246 30540 27252 30552
rect 27304 30540 27310 30592
rect 28644 30580 28672 30611
rect 29270 30608 29276 30620
rect 29328 30608 29334 30660
rect 30193 30651 30251 30657
rect 30193 30648 30205 30651
rect 29380 30620 30205 30648
rect 29380 30580 29408 30620
rect 30193 30617 30205 30620
rect 30239 30617 30251 30651
rect 30193 30611 30251 30617
rect 30285 30651 30343 30657
rect 30285 30617 30297 30651
rect 30331 30648 30343 30651
rect 30331 30620 31340 30648
rect 30331 30617 30343 30620
rect 30285 30611 30343 30617
rect 31312 30592 31340 30620
rect 32306 30608 32312 30660
rect 32364 30608 32370 30660
rect 28644 30552 29408 30580
rect 31294 30540 31300 30592
rect 31352 30580 31358 30592
rect 32769 30583 32827 30589
rect 32769 30580 32781 30583
rect 31352 30552 32781 30580
rect 31352 30540 31358 30552
rect 32769 30549 32781 30552
rect 32815 30549 32827 30583
rect 32769 30543 32827 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 17405 30379 17463 30385
rect 17405 30345 17417 30379
rect 17451 30376 17463 30379
rect 17586 30376 17592 30388
rect 17451 30348 17592 30376
rect 17451 30345 17463 30348
rect 17405 30339 17463 30345
rect 17586 30336 17592 30348
rect 17644 30336 17650 30388
rect 17770 30336 17776 30388
rect 17828 30376 17834 30388
rect 17828 30348 18552 30376
rect 17828 30336 17834 30348
rect 18414 30308 18420 30320
rect 18248 30280 18420 30308
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30240 15991 30243
rect 16114 30240 16120 30252
rect 15979 30212 16120 30240
rect 15979 30209 15991 30212
rect 15933 30203 15991 30209
rect 16114 30200 16120 30212
rect 16172 30200 16178 30252
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 16816 30212 16957 30240
rect 16816 30200 16822 30212
rect 16945 30209 16957 30212
rect 16991 30240 17003 30243
rect 18138 30240 18144 30252
rect 16991 30212 18144 30240
rect 16991 30209 17003 30212
rect 16945 30203 17003 30209
rect 18138 30200 18144 30212
rect 18196 30200 18202 30252
rect 18248 30249 18276 30280
rect 18414 30268 18420 30280
rect 18472 30268 18478 30320
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18322 30200 18328 30252
rect 18380 30240 18386 30252
rect 18524 30249 18552 30348
rect 20530 30336 20536 30388
rect 20588 30376 20594 30388
rect 24578 30376 24584 30388
rect 20588 30348 24584 30376
rect 20588 30336 20594 30348
rect 24578 30336 24584 30348
rect 24636 30376 24642 30388
rect 28166 30376 28172 30388
rect 24636 30348 28172 30376
rect 24636 30336 24642 30348
rect 28166 30336 28172 30348
rect 28224 30336 28230 30388
rect 28350 30336 28356 30388
rect 28408 30376 28414 30388
rect 28537 30379 28595 30385
rect 28537 30376 28549 30379
rect 28408 30348 28549 30376
rect 28408 30336 28414 30348
rect 28537 30345 28549 30348
rect 28583 30345 28595 30379
rect 28537 30339 28595 30345
rect 30006 30336 30012 30388
rect 30064 30376 30070 30388
rect 31021 30379 31079 30385
rect 31021 30376 31033 30379
rect 30064 30348 31033 30376
rect 30064 30336 30070 30348
rect 31021 30345 31033 30348
rect 31067 30345 31079 30379
rect 31021 30339 31079 30345
rect 20073 30311 20131 30317
rect 20073 30277 20085 30311
rect 20119 30308 20131 30311
rect 22278 30308 22284 30320
rect 20119 30280 22284 30308
rect 20119 30277 20131 30280
rect 20073 30271 20131 30277
rect 22278 30268 22284 30280
rect 22336 30268 22342 30320
rect 23014 30268 23020 30320
rect 23072 30308 23078 30320
rect 23109 30311 23167 30317
rect 23109 30308 23121 30311
rect 23072 30280 23121 30308
rect 23072 30268 23078 30280
rect 23109 30277 23121 30280
rect 23155 30277 23167 30311
rect 23109 30271 23167 30277
rect 23569 30311 23627 30317
rect 23569 30277 23581 30311
rect 23615 30308 23627 30311
rect 29365 30311 29423 30317
rect 29365 30308 29377 30311
rect 23615 30280 24716 30308
rect 23615 30277 23627 30280
rect 23569 30271 23627 30277
rect 24688 30252 24716 30280
rect 25873 30280 29377 30308
rect 18509 30243 18567 30249
rect 18380 30212 18425 30240
rect 18380 30200 18386 30212
rect 18509 30209 18521 30243
rect 18555 30209 18567 30243
rect 18509 30203 18567 30209
rect 18969 30243 19027 30249
rect 18969 30209 18981 30243
rect 19015 30209 19027 30243
rect 20898 30240 20904 30252
rect 20859 30212 20904 30240
rect 18969 30203 19027 30209
rect 17770 30132 17776 30184
rect 17828 30172 17834 30184
rect 18984 30172 19012 30203
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 21085 30243 21143 30249
rect 21085 30209 21097 30243
rect 21131 30209 21143 30243
rect 21085 30203 21143 30209
rect 20806 30172 20812 30184
rect 17828 30144 20812 30172
rect 17828 30132 17834 30144
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 17310 30104 17316 30116
rect 17271 30076 17316 30104
rect 17310 30064 17316 30076
rect 17368 30064 17374 30116
rect 21100 30104 21128 30203
rect 21174 30200 21180 30252
rect 21232 30240 21238 30252
rect 23293 30243 23351 30249
rect 21232 30212 21277 30240
rect 21232 30200 21238 30212
rect 23293 30209 23305 30243
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 23477 30243 23535 30249
rect 23477 30209 23489 30243
rect 23523 30240 23535 30243
rect 23658 30240 23664 30252
rect 23523 30212 23664 30240
rect 23523 30209 23535 30212
rect 23477 30203 23535 30209
rect 23308 30172 23336 30203
rect 23658 30200 23664 30212
rect 23716 30240 23722 30252
rect 24029 30243 24087 30249
rect 24029 30240 24041 30243
rect 23716 30212 24041 30240
rect 23716 30200 23722 30212
rect 24029 30209 24041 30212
rect 24075 30209 24087 30243
rect 24394 30240 24400 30252
rect 24355 30212 24400 30240
rect 24029 30203 24087 30209
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 24670 30240 24676 30252
rect 24631 30212 24676 30240
rect 24670 30200 24676 30212
rect 24728 30200 24734 30252
rect 25222 30200 25228 30252
rect 25280 30240 25286 30252
rect 25593 30243 25651 30249
rect 25593 30240 25605 30243
rect 25280 30212 25605 30240
rect 25280 30200 25286 30212
rect 25593 30209 25605 30212
rect 25639 30209 25651 30243
rect 25774 30240 25780 30252
rect 25735 30212 25780 30240
rect 25593 30203 25651 30209
rect 25774 30200 25780 30212
rect 25832 30200 25838 30252
rect 25873 30249 25901 30280
rect 29365 30277 29377 30280
rect 29411 30277 29423 30311
rect 32306 30308 32312 30320
rect 32267 30280 32312 30308
rect 29365 30271 29423 30277
rect 32306 30268 32312 30280
rect 32364 30268 32370 30320
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 27246 30200 27252 30252
rect 27304 30240 27310 30252
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 27304 30212 27353 30240
rect 27304 30200 27310 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 27893 30243 27951 30249
rect 27893 30209 27905 30243
rect 27939 30240 27951 30243
rect 28353 30243 28411 30249
rect 28353 30240 28365 30243
rect 27939 30212 28365 30240
rect 27939 30209 27951 30212
rect 27893 30203 27951 30209
rect 28353 30209 28365 30212
rect 28399 30240 28411 30243
rect 28902 30240 28908 30252
rect 28399 30212 28908 30240
rect 28399 30209 28411 30212
rect 28353 30203 28411 30209
rect 28902 30200 28908 30212
rect 28960 30200 28966 30252
rect 29549 30243 29607 30249
rect 29549 30209 29561 30243
rect 29595 30209 29607 30243
rect 29549 30203 29607 30209
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 30653 30243 30711 30249
rect 30653 30209 30665 30243
rect 30699 30240 30711 30243
rect 31294 30240 31300 30252
rect 30699 30212 31300 30240
rect 30699 30209 30711 30212
rect 30653 30203 30711 30209
rect 23566 30172 23572 30184
rect 23308 30144 23572 30172
rect 23566 30132 23572 30144
rect 23624 30132 23630 30184
rect 24489 30175 24547 30181
rect 24489 30141 24501 30175
rect 24535 30172 24547 30175
rect 24535 30144 25636 30172
rect 24535 30141 24547 30144
rect 24489 30135 24547 30141
rect 21174 30104 21180 30116
rect 21100 30076 21180 30104
rect 21174 30064 21180 30076
rect 21232 30104 21238 30116
rect 25608 30104 25636 30144
rect 25682 30132 25688 30184
rect 25740 30172 25746 30184
rect 25740 30144 25785 30172
rect 25740 30132 25746 30144
rect 27430 30132 27436 30184
rect 27488 30172 27494 30184
rect 28169 30175 28227 30181
rect 28169 30172 28181 30175
rect 27488 30144 28181 30172
rect 27488 30132 27494 30144
rect 28169 30141 28181 30144
rect 28215 30141 28227 30175
rect 28169 30135 28227 30141
rect 28810 30132 28816 30184
rect 28868 30172 28874 30184
rect 29564 30172 29592 30203
rect 28868 30144 29592 30172
rect 28868 30132 28874 30144
rect 26970 30104 26976 30116
rect 21232 30076 25544 30104
rect 25608 30076 26976 30104
rect 21232 30064 21238 30076
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16025 30039 16083 30045
rect 16025 30036 16037 30039
rect 15988 30008 16037 30036
rect 15988 29996 15994 30008
rect 16025 30005 16037 30008
rect 16071 30005 16083 30039
rect 17862 30036 17868 30048
rect 17823 30008 17868 30036
rect 16025 29999 16083 30005
rect 17862 29996 17868 30008
rect 17920 29996 17926 30048
rect 18322 29996 18328 30048
rect 18380 30036 18386 30048
rect 19150 30036 19156 30048
rect 18380 30008 19156 30036
rect 18380 29996 18386 30008
rect 19150 29996 19156 30008
rect 19208 29996 19214 30048
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 20165 30039 20223 30045
rect 20165 30036 20177 30039
rect 19392 30008 20177 30036
rect 19392 29996 19398 30008
rect 20165 30005 20177 30008
rect 20211 30005 20223 30039
rect 20165 29999 20223 30005
rect 20254 29996 20260 30048
rect 20312 30036 20318 30048
rect 20717 30039 20775 30045
rect 20717 30036 20729 30039
rect 20312 30008 20729 30036
rect 20312 29996 20318 30008
rect 20717 30005 20729 30008
rect 20763 30005 20775 30039
rect 20717 29999 20775 30005
rect 20990 29996 20996 30048
rect 21048 30036 21054 30048
rect 25222 30036 25228 30048
rect 21048 30008 25228 30036
rect 21048 29996 21054 30008
rect 25222 29996 25228 30008
rect 25280 29996 25286 30048
rect 25406 30036 25412 30048
rect 25367 30008 25412 30036
rect 25406 29996 25412 30008
rect 25464 29996 25470 30048
rect 25516 30036 25544 30076
rect 26970 30064 26976 30076
rect 27028 30064 27034 30116
rect 27525 30107 27583 30113
rect 27525 30073 27537 30107
rect 27571 30104 27583 30107
rect 28828 30104 28856 30132
rect 27571 30076 28856 30104
rect 29089 30107 29147 30113
rect 27571 30073 27583 30076
rect 27525 30067 27583 30073
rect 29089 30073 29101 30107
rect 29135 30104 29147 30107
rect 29748 30104 29776 30203
rect 31294 30200 31300 30212
rect 31352 30200 31358 30252
rect 32217 30243 32275 30249
rect 32217 30209 32229 30243
rect 32263 30240 32275 30243
rect 33318 30240 33324 30252
rect 32263 30212 33324 30240
rect 32263 30209 32275 30212
rect 32217 30203 32275 30209
rect 33318 30200 33324 30212
rect 33376 30200 33382 30252
rect 30745 30175 30803 30181
rect 30745 30141 30757 30175
rect 30791 30172 30803 30175
rect 30834 30172 30840 30184
rect 30791 30144 30840 30172
rect 30791 30141 30803 30144
rect 30745 30135 30803 30141
rect 30834 30132 30840 30144
rect 30892 30132 30898 30184
rect 47946 30104 47952 30116
rect 29135 30076 47952 30104
rect 29135 30073 29147 30076
rect 29089 30067 29147 30073
rect 47946 30064 47952 30076
rect 48004 30064 48010 30116
rect 28258 30036 28264 30048
rect 25516 30008 28264 30036
rect 28258 29996 28264 30008
rect 28316 29996 28322 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 16758 29832 16764 29844
rect 16719 29804 16764 29832
rect 16758 29792 16764 29804
rect 16816 29792 16822 29844
rect 21637 29835 21695 29841
rect 21637 29801 21649 29835
rect 21683 29832 21695 29835
rect 22186 29832 22192 29844
rect 21683 29804 22192 29832
rect 21683 29801 21695 29804
rect 21637 29795 21695 29801
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 25574 29835 25632 29841
rect 25574 29832 25586 29835
rect 25464 29804 25586 29832
rect 25464 29792 25470 29804
rect 25574 29801 25586 29804
rect 25620 29801 25632 29835
rect 25574 29795 25632 29801
rect 28353 29835 28411 29841
rect 28353 29801 28365 29835
rect 28399 29832 28411 29835
rect 28442 29832 28448 29844
rect 28399 29804 28448 29832
rect 28399 29801 28411 29804
rect 28353 29795 28411 29801
rect 28442 29792 28448 29804
rect 28500 29792 28506 29844
rect 29638 29792 29644 29844
rect 29696 29832 29702 29844
rect 31846 29832 31852 29844
rect 29696 29804 31852 29832
rect 29696 29792 29702 29804
rect 31846 29792 31852 29804
rect 31904 29832 31910 29844
rect 32217 29835 32275 29841
rect 32217 29832 32229 29835
rect 31904 29804 32229 29832
rect 31904 29792 31910 29804
rect 32217 29801 32229 29804
rect 32263 29801 32275 29835
rect 32217 29795 32275 29801
rect 21542 29724 21548 29776
rect 21600 29764 21606 29776
rect 23477 29767 23535 29773
rect 21600 29736 23336 29764
rect 21600 29724 21606 29736
rect 15013 29699 15071 29705
rect 15013 29665 15025 29699
rect 15059 29696 15071 29699
rect 16022 29696 16028 29708
rect 15059 29668 16028 29696
rect 15059 29665 15071 29668
rect 15013 29659 15071 29665
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 17402 29656 17408 29708
rect 17460 29696 17466 29708
rect 17681 29699 17739 29705
rect 17681 29696 17693 29699
rect 17460 29668 17693 29696
rect 17460 29656 17466 29668
rect 17681 29665 17693 29668
rect 17727 29665 17739 29699
rect 17681 29659 17739 29665
rect 17770 29656 17776 29708
rect 17828 29696 17834 29708
rect 17828 29668 17873 29696
rect 17828 29656 17834 29668
rect 20714 29656 20720 29708
rect 20772 29696 20778 29708
rect 22002 29696 22008 29708
rect 20772 29668 22008 29696
rect 20772 29656 20778 29668
rect 22002 29656 22008 29668
rect 22060 29696 22066 29708
rect 22741 29699 22799 29705
rect 22741 29696 22753 29699
rect 22060 29668 22753 29696
rect 22060 29656 22066 29668
rect 22741 29665 22753 29668
rect 22787 29665 22799 29699
rect 22741 29659 22799 29665
rect 17862 29588 17868 29640
rect 17920 29628 17926 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 17920 29600 19441 29628
rect 17920 29588 17926 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29628 19763 29631
rect 19978 29628 19984 29640
rect 19751 29600 19984 29628
rect 19751 29597 19763 29600
rect 19705 29591 19763 29597
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 21269 29631 21327 29637
rect 21269 29597 21281 29631
rect 21315 29597 21327 29631
rect 21269 29591 21327 29597
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29628 21695 29631
rect 22281 29631 22339 29637
rect 22281 29628 22293 29631
rect 21683 29600 22293 29628
rect 21683 29597 21695 29600
rect 21637 29591 21695 29597
rect 22281 29597 22293 29600
rect 22327 29597 22339 29631
rect 22462 29628 22468 29640
rect 22423 29600 22468 29628
rect 22281 29591 22339 29597
rect 15286 29560 15292 29572
rect 15247 29532 15292 29560
rect 15286 29520 15292 29532
rect 15344 29520 15350 29572
rect 15930 29520 15936 29572
rect 15988 29520 15994 29572
rect 17310 29520 17316 29572
rect 17368 29560 17374 29572
rect 19613 29563 19671 29569
rect 17368 29532 19380 29560
rect 17368 29520 17374 29532
rect 17218 29492 17224 29504
rect 17179 29464 17224 29492
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 17589 29495 17647 29501
rect 17589 29492 17601 29495
rect 17552 29464 17601 29492
rect 17552 29452 17558 29464
rect 17589 29461 17601 29464
rect 17635 29461 17647 29495
rect 17589 29455 17647 29461
rect 17678 29452 17684 29504
rect 17736 29492 17742 29504
rect 19245 29495 19303 29501
rect 19245 29492 19257 29495
rect 17736 29464 19257 29492
rect 17736 29452 17742 29464
rect 19245 29461 19257 29464
rect 19291 29461 19303 29495
rect 19352 29492 19380 29532
rect 19613 29529 19625 29563
rect 19659 29560 19671 29563
rect 20990 29560 20996 29572
rect 19659 29532 20996 29560
rect 19659 29529 19671 29532
rect 19613 29523 19671 29529
rect 20990 29520 20996 29532
rect 21048 29520 21054 29572
rect 21284 29560 21312 29591
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22649 29631 22707 29637
rect 22649 29597 22661 29631
rect 22695 29628 22707 29631
rect 23198 29628 23204 29640
rect 22695 29600 23204 29628
rect 22695 29597 22707 29600
rect 22649 29591 22707 29597
rect 23198 29588 23204 29600
rect 23256 29588 23262 29640
rect 23308 29637 23336 29736
rect 23477 29733 23489 29767
rect 23523 29764 23535 29767
rect 23658 29764 23664 29776
rect 23523 29736 23664 29764
rect 23523 29733 23535 29736
rect 23477 29727 23535 29733
rect 23658 29724 23664 29736
rect 23716 29724 23722 29776
rect 24397 29767 24455 29773
rect 24397 29733 24409 29767
rect 24443 29764 24455 29767
rect 24854 29764 24860 29776
rect 24443 29736 24860 29764
rect 24443 29733 24455 29736
rect 24397 29727 24455 29733
rect 24854 29724 24860 29736
rect 24912 29724 24918 29776
rect 26694 29724 26700 29776
rect 26752 29764 26758 29776
rect 27430 29764 27436 29776
rect 26752 29736 27436 29764
rect 26752 29724 26758 29736
rect 27430 29724 27436 29736
rect 27488 29764 27494 29776
rect 27801 29767 27859 29773
rect 27801 29764 27813 29767
rect 27488 29736 27813 29764
rect 27488 29724 27494 29736
rect 27801 29733 27813 29736
rect 27847 29733 27859 29767
rect 30558 29764 30564 29776
rect 27801 29727 27859 29733
rect 29564 29736 30564 29764
rect 25317 29699 25375 29705
rect 25317 29665 25329 29699
rect 25363 29696 25375 29699
rect 26234 29696 26240 29708
rect 25363 29668 26240 29696
rect 25363 29665 25375 29668
rect 25317 29659 25375 29665
rect 26234 29656 26240 29668
rect 26292 29656 26298 29708
rect 26970 29656 26976 29708
rect 27028 29696 27034 29708
rect 29564 29696 29592 29736
rect 30558 29724 30564 29736
rect 30616 29764 30622 29776
rect 30616 29736 31754 29764
rect 30616 29724 30622 29736
rect 27028 29668 29592 29696
rect 27028 29656 27034 29668
rect 23293 29631 23351 29637
rect 23293 29597 23305 29631
rect 23339 29628 23351 29631
rect 23474 29628 23480 29640
rect 23339 29600 23480 29628
rect 23339 29597 23351 29600
rect 23293 29591 23351 29597
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 24670 29628 24676 29640
rect 24631 29600 24676 29628
rect 24670 29588 24676 29600
rect 24728 29588 24734 29640
rect 27062 29588 27068 29640
rect 27120 29628 27126 29640
rect 29564 29637 29592 29668
rect 30834 29656 30840 29708
rect 30892 29696 30898 29708
rect 31481 29699 31539 29705
rect 31481 29696 31493 29699
rect 30892 29668 31493 29696
rect 30892 29656 30898 29668
rect 31481 29665 31493 29668
rect 31527 29665 31539 29699
rect 31481 29659 31539 29665
rect 28261 29631 28319 29637
rect 28261 29628 28273 29631
rect 27120 29600 28273 29628
rect 27120 29588 27126 29600
rect 28261 29597 28273 29600
rect 28307 29597 28319 29631
rect 28261 29591 28319 29597
rect 29549 29631 29607 29637
rect 29549 29597 29561 29631
rect 29595 29597 29607 29631
rect 29549 29591 29607 29597
rect 30285 29631 30343 29637
rect 30285 29597 30297 29631
rect 30331 29628 30343 29631
rect 31110 29628 31116 29640
rect 30331 29600 31116 29628
rect 30331 29597 30343 29600
rect 30285 29591 30343 29597
rect 31110 29588 31116 29600
rect 31168 29588 31174 29640
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29597 31355 29631
rect 31297 29591 31355 29597
rect 22094 29560 22100 29572
rect 21284 29532 22100 29560
rect 22094 29520 22100 29532
rect 22152 29560 22158 29572
rect 23382 29560 23388 29572
rect 22152 29532 23388 29560
rect 22152 29520 22158 29532
rect 23382 29520 23388 29532
rect 23440 29520 23446 29572
rect 23566 29520 23572 29572
rect 23624 29560 23630 29572
rect 24397 29563 24455 29569
rect 24397 29560 24409 29563
rect 23624 29532 24409 29560
rect 23624 29520 23630 29532
rect 24397 29529 24409 29532
rect 24443 29560 24455 29563
rect 25130 29560 25136 29572
rect 24443 29532 25136 29560
rect 24443 29529 24455 29532
rect 24397 29523 24455 29529
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 26970 29560 26976 29572
rect 26818 29532 26976 29560
rect 26970 29520 26976 29532
rect 27028 29520 27034 29572
rect 27614 29560 27620 29572
rect 27527 29532 27620 29560
rect 27614 29520 27620 29532
rect 27672 29560 27678 29572
rect 29822 29560 29828 29572
rect 27672 29532 29828 29560
rect 27672 29520 27678 29532
rect 29822 29520 29828 29532
rect 29880 29520 29886 29572
rect 30469 29563 30527 29569
rect 30469 29529 30481 29563
rect 30515 29560 30527 29563
rect 30834 29560 30840 29572
rect 30515 29532 30840 29560
rect 30515 29529 30527 29532
rect 30469 29523 30527 29529
rect 30834 29520 30840 29532
rect 30892 29520 30898 29572
rect 31312 29560 31340 29591
rect 31386 29588 31392 29640
rect 31444 29628 31450 29640
rect 31573 29631 31631 29637
rect 31573 29628 31585 29631
rect 31444 29600 31585 29628
rect 31444 29588 31450 29600
rect 31573 29597 31585 29600
rect 31619 29597 31631 29631
rect 31726 29628 31754 29736
rect 45370 29656 45376 29708
rect 45428 29696 45434 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 45428 29668 47593 29696
rect 45428 29656 45434 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 32125 29631 32183 29637
rect 32125 29628 32137 29631
rect 31726 29600 32137 29628
rect 31573 29591 31631 29597
rect 32125 29597 32137 29600
rect 32171 29597 32183 29631
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 32125 29591 32183 29597
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 31312 29532 31616 29560
rect 31588 29504 31616 29532
rect 21542 29492 21548 29504
rect 19352 29464 21548 29492
rect 19245 29455 19303 29461
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 21818 29492 21824 29504
rect 21779 29464 21824 29492
rect 21818 29452 21824 29464
rect 21876 29452 21882 29504
rect 23658 29452 23664 29504
rect 23716 29492 23722 29504
rect 24581 29495 24639 29501
rect 24581 29492 24593 29495
rect 23716 29464 24593 29492
rect 23716 29452 23722 29464
rect 24581 29461 24593 29464
rect 24627 29461 24639 29495
rect 24581 29455 24639 29461
rect 25222 29452 25228 29504
rect 25280 29492 25286 29504
rect 27065 29495 27123 29501
rect 27065 29492 27077 29495
rect 25280 29464 27077 29492
rect 25280 29452 25286 29464
rect 27065 29461 27077 29464
rect 27111 29461 27123 29495
rect 27065 29455 27123 29461
rect 29178 29452 29184 29504
rect 29236 29492 29242 29504
rect 29733 29495 29791 29501
rect 29733 29492 29745 29495
rect 29236 29464 29745 29492
rect 29236 29452 29242 29464
rect 29733 29461 29745 29464
rect 29779 29492 29791 29495
rect 30282 29492 30288 29504
rect 29779 29464 30288 29492
rect 29779 29461 29791 29464
rect 29733 29455 29791 29461
rect 30282 29452 30288 29464
rect 30340 29452 30346 29504
rect 30650 29492 30656 29504
rect 30611 29464 30656 29492
rect 30650 29452 30656 29464
rect 30708 29452 30714 29504
rect 31113 29495 31171 29501
rect 31113 29461 31125 29495
rect 31159 29492 31171 29495
rect 31202 29492 31208 29504
rect 31159 29464 31208 29492
rect 31159 29461 31171 29464
rect 31113 29455 31171 29461
rect 31202 29452 31208 29464
rect 31260 29452 31266 29504
rect 31570 29452 31576 29504
rect 31628 29452 31634 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 2406 29248 2412 29300
rect 2464 29288 2470 29300
rect 20533 29291 20591 29297
rect 2464 29260 20484 29288
rect 2464 29248 2470 29260
rect 17218 29220 17224 29232
rect 15948 29192 17224 29220
rect 15948 29161 15976 29192
rect 17218 29180 17224 29192
rect 17276 29180 17282 29232
rect 19334 29220 19340 29232
rect 18800 29192 19340 29220
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29121 15991 29155
rect 15933 29115 15991 29121
rect 16022 29112 16028 29164
rect 16080 29152 16086 29164
rect 18800 29161 18828 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20070 29180 20076 29232
rect 20128 29180 20134 29232
rect 20456 29220 20484 29260
rect 20533 29257 20545 29291
rect 20579 29288 20591 29291
rect 20714 29288 20720 29300
rect 20579 29260 20720 29288
rect 20579 29257 20591 29260
rect 20533 29251 20591 29257
rect 20714 29248 20720 29260
rect 20772 29248 20778 29300
rect 22186 29288 22192 29300
rect 21928 29260 22192 29288
rect 21928 29220 21956 29260
rect 22186 29248 22192 29260
rect 22244 29248 22250 29300
rect 23382 29288 23388 29300
rect 23343 29260 23388 29288
rect 23382 29248 23388 29260
rect 23440 29248 23446 29300
rect 23474 29248 23480 29300
rect 23532 29288 23538 29300
rect 25038 29288 25044 29300
rect 23532 29260 25044 29288
rect 23532 29248 23538 29260
rect 25038 29248 25044 29260
rect 25096 29288 25102 29300
rect 26142 29288 26148 29300
rect 25096 29260 26148 29288
rect 25096 29248 25102 29260
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 27154 29288 27160 29300
rect 27115 29260 27160 29288
rect 27154 29248 27160 29260
rect 27212 29248 27218 29300
rect 31481 29291 31539 29297
rect 31481 29257 31493 29291
rect 31527 29257 31539 29291
rect 31481 29251 31539 29257
rect 20456 29192 21956 29220
rect 26326 29180 26332 29232
rect 26384 29220 26390 29232
rect 27065 29223 27123 29229
rect 27065 29220 27077 29223
rect 26384 29192 27077 29220
rect 26384 29180 26390 29192
rect 27065 29189 27077 29192
rect 27111 29189 27123 29223
rect 29825 29223 29883 29229
rect 29825 29220 29837 29223
rect 27065 29183 27123 29189
rect 28000 29192 29837 29220
rect 18785 29155 18843 29161
rect 18785 29152 18797 29155
rect 16080 29124 18797 29152
rect 16080 29112 16086 29124
rect 18785 29121 18797 29124
rect 18831 29121 18843 29155
rect 21818 29152 21824 29164
rect 21779 29124 21824 29152
rect 18785 29115 18843 29121
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 22278 29162 22284 29164
rect 21993 29153 22051 29159
rect 21993 29119 22005 29153
rect 22039 29119 22051 29153
rect 21993 29113 22051 29119
rect 22112 29134 22284 29162
rect 19061 29087 19119 29093
rect 19061 29053 19073 29087
rect 19107 29084 19119 29087
rect 20254 29084 20260 29096
rect 19107 29056 20260 29084
rect 19107 29053 19119 29056
rect 19061 29047 19119 29053
rect 20254 29044 20260 29056
rect 20312 29044 20318 29096
rect 21542 29044 21548 29096
rect 21600 29084 21606 29096
rect 22008 29084 22036 29113
rect 22112 29093 22140 29134
rect 22278 29112 22284 29134
rect 22336 29112 22342 29164
rect 22373 29155 22431 29161
rect 22373 29121 22385 29155
rect 22419 29152 22431 29155
rect 23014 29152 23020 29164
rect 22419 29124 22876 29152
rect 22975 29124 23020 29152
rect 22419 29121 22431 29124
rect 22373 29115 22431 29121
rect 21600 29056 22036 29084
rect 22097 29087 22155 29093
rect 21600 29044 21606 29056
rect 22097 29053 22109 29087
rect 22143 29053 22155 29087
rect 22097 29047 22155 29053
rect 22186 29044 22192 29096
rect 22244 29084 22250 29096
rect 22244 29056 22289 29084
rect 22244 29044 22250 29056
rect 15286 28976 15292 29028
rect 15344 29016 15350 29028
rect 15749 29019 15807 29025
rect 15749 29016 15761 29019
rect 15344 28988 15761 29016
rect 15344 28976 15350 28988
rect 15749 28985 15761 28988
rect 15795 28985 15807 29019
rect 15749 28979 15807 28985
rect 21082 28976 21088 29028
rect 21140 29016 21146 29028
rect 22557 29019 22615 29025
rect 22557 29016 22569 29019
rect 21140 28988 22569 29016
rect 21140 28976 21146 28988
rect 22557 28985 22569 28988
rect 22603 28985 22615 29019
rect 22848 29016 22876 29124
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 23198 29112 23204 29164
rect 23256 29152 23262 29164
rect 24673 29155 24731 29161
rect 23256 29124 23349 29152
rect 23256 29112 23262 29124
rect 24673 29121 24685 29155
rect 24719 29152 24731 29155
rect 24854 29152 24860 29164
rect 24719 29124 24860 29152
rect 24719 29121 24731 29124
rect 24673 29115 24731 29121
rect 24854 29112 24860 29124
rect 24912 29112 24918 29164
rect 25590 29112 25596 29164
rect 25648 29152 25654 29164
rect 28000 29152 28028 29192
rect 29825 29189 29837 29192
rect 29871 29220 29883 29223
rect 30650 29220 30656 29232
rect 29871 29192 30656 29220
rect 29871 29189 29883 29192
rect 29825 29183 29883 29189
rect 30650 29180 30656 29192
rect 30708 29180 30714 29232
rect 31496 29220 31524 29251
rect 31570 29248 31576 29300
rect 31628 29288 31634 29300
rect 32306 29288 32312 29300
rect 31628 29260 32312 29288
rect 31628 29248 31634 29260
rect 32306 29248 32312 29260
rect 32364 29288 32370 29300
rect 34333 29291 34391 29297
rect 34333 29288 34345 29291
rect 32364 29260 34345 29288
rect 32364 29248 32370 29260
rect 34333 29257 34345 29260
rect 34379 29257 34391 29291
rect 34333 29251 34391 29257
rect 31496 29192 31754 29220
rect 25648 29124 28028 29152
rect 28077 29155 28135 29161
rect 25648 29112 25654 29124
rect 28077 29121 28089 29155
rect 28123 29152 28135 29155
rect 28810 29152 28816 29164
rect 28123 29124 28816 29152
rect 28123 29121 28135 29124
rect 28077 29115 28135 29121
rect 28810 29112 28816 29124
rect 28868 29112 28874 29164
rect 30742 29112 30748 29164
rect 30800 29152 30806 29164
rect 30929 29155 30987 29161
rect 30929 29152 30941 29155
rect 30800 29124 30941 29152
rect 30800 29112 30806 29124
rect 30929 29121 30941 29124
rect 30975 29121 30987 29155
rect 31202 29152 31208 29164
rect 31163 29124 31208 29152
rect 30929 29115 30987 29121
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 23216 29084 23244 29112
rect 23216 29056 29592 29084
rect 23474 29016 23480 29028
rect 22848 28988 23480 29016
rect 22557 28979 22615 28985
rect 23474 28976 23480 28988
rect 23532 28976 23538 29028
rect 24578 28976 24584 29028
rect 24636 29016 24642 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 24636 28988 24869 29016
rect 24636 28976 24642 28988
rect 24857 28985 24869 28988
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 25130 28976 25136 29028
rect 25188 29016 25194 29028
rect 27614 29016 27620 29028
rect 25188 28988 27620 29016
rect 25188 28976 25194 28988
rect 27614 28976 27620 28988
rect 27672 28976 27678 29028
rect 28258 29016 28264 29028
rect 28219 28988 28264 29016
rect 28258 28976 28264 28988
rect 28316 28976 28322 29028
rect 29564 28960 29592 29056
rect 31726 29016 31754 29192
rect 33410 29180 33416 29232
rect 33468 29180 33474 29232
rect 32582 29084 32588 29096
rect 32543 29056 32588 29084
rect 32582 29044 32588 29056
rect 32640 29044 32646 29096
rect 32858 29084 32864 29096
rect 32819 29056 32864 29084
rect 32858 29044 32864 29056
rect 32916 29044 32922 29096
rect 32030 29016 32036 29028
rect 31404 28988 31616 29016
rect 31726 28988 32036 29016
rect 19150 28908 19156 28960
rect 19208 28948 19214 28960
rect 26878 28948 26884 28960
rect 19208 28920 26884 28948
rect 19208 28908 19214 28920
rect 26878 28908 26884 28920
rect 26936 28908 26942 28960
rect 29546 28908 29552 28960
rect 29604 28948 29610 28960
rect 29917 28951 29975 28957
rect 29917 28948 29929 28951
rect 29604 28920 29929 28948
rect 29604 28908 29610 28920
rect 29917 28917 29929 28920
rect 29963 28917 29975 28951
rect 29917 28911 29975 28917
rect 30006 28908 30012 28960
rect 30064 28948 30070 28960
rect 30742 28948 30748 28960
rect 30064 28920 30748 28948
rect 30064 28908 30070 28920
rect 30742 28908 30748 28920
rect 30800 28908 30806 28960
rect 31297 28951 31355 28957
rect 31297 28917 31309 28951
rect 31343 28948 31355 28951
rect 31404 28948 31432 28988
rect 31343 28920 31432 28948
rect 31588 28948 31616 28988
rect 32030 28976 32036 28988
rect 32088 28976 32094 29028
rect 31846 28948 31852 28960
rect 31588 28920 31852 28948
rect 31343 28917 31355 28920
rect 31297 28911 31355 28917
rect 31846 28908 31852 28920
rect 31904 28908 31910 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 15552 28747 15610 28753
rect 15552 28713 15564 28747
rect 15598 28744 15610 28747
rect 17678 28744 17684 28756
rect 15598 28716 17684 28744
rect 15598 28713 15610 28716
rect 15552 28707 15610 28713
rect 17678 28704 17684 28716
rect 17736 28704 17742 28756
rect 22278 28704 22284 28756
rect 22336 28744 22342 28756
rect 25314 28744 25320 28756
rect 22336 28716 25320 28744
rect 22336 28704 22342 28716
rect 25314 28704 25320 28716
rect 25372 28704 25378 28756
rect 26970 28704 26976 28756
rect 27028 28744 27034 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 27028 28716 27077 28744
rect 27028 28704 27034 28716
rect 27065 28713 27077 28716
rect 27111 28713 27123 28747
rect 27065 28707 27123 28713
rect 29638 28704 29644 28756
rect 29696 28744 29702 28756
rect 30653 28747 30711 28753
rect 30653 28744 30665 28747
rect 29696 28716 30665 28744
rect 29696 28704 29702 28716
rect 30653 28713 30665 28716
rect 30699 28713 30711 28747
rect 31110 28744 31116 28756
rect 31071 28716 31116 28744
rect 30653 28707 30711 28713
rect 31110 28704 31116 28716
rect 31168 28704 31174 28756
rect 32769 28747 32827 28753
rect 32769 28713 32781 28747
rect 32815 28744 32827 28747
rect 32858 28744 32864 28756
rect 32815 28716 32864 28744
rect 32815 28713 32827 28716
rect 32769 28707 32827 28713
rect 32858 28704 32864 28716
rect 32916 28704 32922 28756
rect 33410 28744 33416 28756
rect 33371 28716 33416 28744
rect 33410 28704 33416 28716
rect 33468 28704 33474 28756
rect 44082 28744 44088 28756
rect 35866 28716 44088 28744
rect 17034 28676 17040 28688
rect 16995 28648 17040 28676
rect 17034 28636 17040 28648
rect 17092 28636 17098 28688
rect 35866 28676 35894 28716
rect 44082 28704 44088 28716
rect 44140 28704 44146 28756
rect 25148 28648 35894 28676
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28608 15347 28611
rect 16022 28608 16028 28620
rect 15335 28580 16028 28608
rect 15335 28577 15347 28580
rect 15289 28571 15347 28577
rect 16022 28568 16028 28580
rect 16080 28568 16086 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 21082 28608 21088 28620
rect 20119 28580 21088 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 21082 28568 21088 28580
rect 21140 28568 21146 28620
rect 21545 28611 21603 28617
rect 21545 28577 21557 28611
rect 21591 28608 21603 28611
rect 22462 28608 22468 28620
rect 21591 28580 22468 28608
rect 21591 28577 21603 28580
rect 21545 28571 21603 28577
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 22204 28549 22232 28580
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 22738 28568 22744 28620
rect 22796 28608 22802 28620
rect 23658 28608 23664 28620
rect 22796 28580 23664 28608
rect 22796 28568 22802 28580
rect 23658 28568 23664 28580
rect 23716 28608 23722 28620
rect 23716 28580 23796 28608
rect 23716 28568 23722 28580
rect 19797 28543 19855 28549
rect 19797 28540 19809 28543
rect 19392 28512 19809 28540
rect 19392 28500 19398 28512
rect 19797 28509 19809 28512
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28540 22247 28543
rect 23566 28540 23572 28552
rect 22235 28512 22269 28540
rect 23527 28512 23572 28540
rect 22235 28509 22247 28512
rect 22189 28503 22247 28509
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 23768 28549 23796 28580
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 24578 28500 24584 28552
rect 24636 28540 24642 28552
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 24636 28512 24777 28540
rect 24636 28500 24642 28512
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 24854 28500 24860 28552
rect 24912 28540 24918 28552
rect 25148 28549 25176 28648
rect 26694 28608 26700 28620
rect 25332 28580 26700 28608
rect 24949 28543 25007 28549
rect 24949 28540 24961 28543
rect 24912 28512 24961 28540
rect 24912 28500 24918 28512
rect 24949 28509 24961 28512
rect 24995 28509 25007 28543
rect 24949 28503 25007 28509
rect 25133 28543 25191 28549
rect 25133 28509 25145 28543
rect 25179 28509 25191 28543
rect 25133 28503 25191 28509
rect 16574 28432 16580 28484
rect 16632 28432 16638 28484
rect 20806 28432 20812 28484
rect 20864 28432 20870 28484
rect 22002 28472 22008 28484
rect 21963 28444 22008 28472
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 25041 28475 25099 28481
rect 25041 28472 25053 28475
rect 22612 28444 25053 28472
rect 22612 28432 22618 28444
rect 25041 28441 25053 28444
rect 25087 28472 25099 28475
rect 25332 28472 25360 28580
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 30837 28611 30895 28617
rect 30837 28577 30849 28611
rect 30883 28608 30895 28611
rect 31386 28608 31392 28620
rect 30883 28580 31392 28608
rect 30883 28577 30895 28580
rect 30837 28571 30895 28577
rect 31386 28568 31392 28580
rect 31444 28608 31450 28620
rect 32306 28608 32312 28620
rect 31444 28580 32312 28608
rect 31444 28568 31450 28580
rect 32306 28568 32312 28580
rect 32364 28568 32370 28620
rect 32401 28611 32459 28617
rect 32401 28577 32413 28611
rect 32447 28608 32459 28611
rect 43990 28608 43996 28620
rect 32447 28580 43996 28608
rect 32447 28577 32459 28580
rect 32401 28571 32459 28577
rect 43990 28568 43996 28580
rect 44048 28568 44054 28620
rect 25406 28500 25412 28552
rect 25464 28540 25470 28552
rect 25961 28543 26019 28549
rect 25961 28540 25973 28543
rect 25464 28512 25973 28540
rect 25464 28500 25470 28512
rect 25961 28509 25973 28512
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27062 28540 27068 28552
rect 27019 28512 27068 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27062 28500 27068 28512
rect 27120 28500 27126 28552
rect 27154 28500 27160 28552
rect 27212 28540 27218 28552
rect 27801 28543 27859 28549
rect 27801 28540 27813 28543
rect 27212 28512 27813 28540
rect 27212 28500 27218 28512
rect 27801 28509 27813 28512
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 27982 28500 27988 28552
rect 28040 28540 28046 28552
rect 28537 28543 28595 28549
rect 28537 28540 28549 28543
rect 28040 28512 28549 28540
rect 28040 28500 28046 28512
rect 28537 28509 28549 28512
rect 28583 28540 28595 28543
rect 28718 28540 28724 28552
rect 28583 28512 28724 28540
rect 28583 28509 28595 28512
rect 28537 28503 28595 28509
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 29086 28500 29092 28552
rect 29144 28540 29150 28552
rect 29638 28540 29644 28552
rect 29144 28512 29644 28540
rect 29144 28500 29150 28512
rect 29638 28500 29644 28512
rect 29696 28500 29702 28552
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 30006 28540 30012 28552
rect 29779 28512 30012 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 30006 28500 30012 28512
rect 30064 28500 30070 28552
rect 30098 28500 30104 28552
rect 30156 28540 30162 28552
rect 30929 28543 30987 28549
rect 30929 28540 30941 28543
rect 30156 28538 30696 28540
rect 30852 28538 30941 28540
rect 30156 28512 30941 28538
rect 30156 28500 30162 28512
rect 30668 28510 30880 28512
rect 30929 28509 30941 28512
rect 30975 28509 30987 28543
rect 32030 28540 32036 28552
rect 31991 28512 32036 28540
rect 30929 28503 30987 28509
rect 32030 28500 32036 28512
rect 32088 28500 32094 28552
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 25087 28444 25360 28472
rect 25777 28475 25835 28481
rect 25087 28441 25099 28444
rect 25041 28435 25099 28441
rect 25777 28441 25789 28475
rect 25823 28441 25835 28475
rect 25777 28435 25835 28441
rect 22373 28407 22431 28413
rect 22373 28373 22385 28407
rect 22419 28404 22431 28407
rect 23014 28404 23020 28416
rect 22419 28376 23020 28404
rect 22419 28373 22431 28376
rect 22373 28367 22431 28373
rect 23014 28364 23020 28376
rect 23072 28404 23078 28416
rect 23198 28404 23204 28416
rect 23072 28376 23204 28404
rect 23072 28364 23078 28376
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23753 28407 23811 28413
rect 23753 28373 23765 28407
rect 23799 28404 23811 28407
rect 25130 28404 25136 28416
rect 23799 28376 25136 28404
rect 23799 28373 23811 28376
rect 23753 28367 23811 28373
rect 25130 28364 25136 28376
rect 25188 28364 25194 28416
rect 25317 28407 25375 28413
rect 25317 28373 25329 28407
rect 25363 28404 25375 28407
rect 25792 28404 25820 28435
rect 26050 28432 26056 28484
rect 26108 28472 26114 28484
rect 30653 28475 30711 28481
rect 26108 28444 30052 28472
rect 26108 28432 26114 28444
rect 25363 28376 25820 28404
rect 26145 28407 26203 28413
rect 25363 28373 25375 28376
rect 25317 28367 25375 28373
rect 26145 28373 26157 28407
rect 26191 28404 26203 28407
rect 26326 28404 26332 28416
rect 26191 28376 26332 28404
rect 26191 28373 26203 28376
rect 26145 28367 26203 28373
rect 26326 28364 26332 28376
rect 26384 28364 26390 28416
rect 27890 28404 27896 28416
rect 27851 28376 27896 28404
rect 27890 28364 27896 28376
rect 27948 28364 27954 28416
rect 28736 28413 28764 28444
rect 28721 28407 28779 28413
rect 28721 28373 28733 28407
rect 28767 28373 28779 28407
rect 29914 28404 29920 28416
rect 29875 28376 29920 28404
rect 28721 28367 28779 28373
rect 29914 28364 29920 28376
rect 29972 28364 29978 28416
rect 30024 28404 30052 28444
rect 30653 28441 30665 28475
rect 30699 28472 30711 28475
rect 31202 28472 31208 28484
rect 30699 28444 31208 28472
rect 30699 28441 30711 28444
rect 30653 28435 30711 28441
rect 31202 28432 31208 28444
rect 31260 28432 31266 28484
rect 32232 28404 32260 28503
rect 32490 28500 32496 28552
rect 32548 28540 32554 28552
rect 32585 28543 32643 28549
rect 32585 28540 32597 28543
rect 32548 28512 32597 28540
rect 32548 28500 32554 28512
rect 32585 28509 32597 28512
rect 32631 28509 32643 28543
rect 33318 28540 33324 28552
rect 33279 28512 33324 28540
rect 32585 28503 32643 28509
rect 33318 28500 33324 28512
rect 33376 28500 33382 28552
rect 32306 28404 32312 28416
rect 30024 28376 32312 28404
rect 32306 28364 32312 28376
rect 32364 28364 32370 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 19981 28203 20039 28209
rect 19981 28169 19993 28203
rect 20027 28200 20039 28203
rect 20070 28200 20076 28212
rect 20027 28172 20076 28200
rect 20027 28169 20039 28172
rect 19981 28163 20039 28169
rect 20070 28160 20076 28172
rect 20128 28160 20134 28212
rect 20806 28200 20812 28212
rect 20767 28172 20812 28200
rect 20806 28160 20812 28172
rect 20864 28160 20870 28212
rect 24489 28203 24547 28209
rect 24489 28200 24501 28203
rect 23216 28172 24501 28200
rect 23216 28166 23244 28172
rect 8404 28104 12434 28132
rect 8404 28073 8432 28104
rect 8389 28067 8447 28073
rect 8389 28033 8401 28067
rect 8435 28033 8447 28067
rect 12406 28064 12434 28104
rect 13446 28092 13452 28144
rect 13504 28132 13510 28144
rect 13725 28135 13783 28141
rect 13504 28104 13676 28132
rect 13504 28092 13510 28104
rect 13538 28064 13544 28076
rect 12406 28036 13544 28064
rect 8389 28027 8447 28033
rect 13538 28024 13544 28036
rect 13596 28024 13602 28076
rect 13648 28064 13676 28104
rect 13725 28101 13737 28135
rect 13771 28132 13783 28135
rect 14182 28132 14188 28144
rect 13771 28104 14188 28132
rect 13771 28101 13783 28104
rect 13725 28095 13783 28101
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 18046 28132 18052 28144
rect 14516 28104 18052 28132
rect 14516 28092 14522 28104
rect 18046 28092 18052 28104
rect 18104 28092 18110 28144
rect 22278 28132 22284 28144
rect 22239 28104 22284 28132
rect 22278 28092 22284 28104
rect 22336 28092 22342 28144
rect 22373 28135 22431 28141
rect 22373 28101 22385 28135
rect 22419 28132 22431 28135
rect 22738 28132 22744 28144
rect 22419 28104 22744 28132
rect 22419 28101 22431 28104
rect 22373 28095 22431 28101
rect 22738 28092 22744 28104
rect 22796 28092 22802 28144
rect 23124 28141 23244 28166
rect 24489 28169 24501 28172
rect 24535 28169 24547 28203
rect 24489 28163 24547 28169
rect 24949 28203 25007 28209
rect 24949 28169 24961 28203
rect 24995 28200 25007 28203
rect 25774 28200 25780 28212
rect 24995 28172 25780 28200
rect 24995 28169 25007 28172
rect 24949 28163 25007 28169
rect 25774 28160 25780 28172
rect 25832 28160 25838 28212
rect 28629 28203 28687 28209
rect 28629 28169 28641 28203
rect 28675 28169 28687 28203
rect 28629 28163 28687 28169
rect 29641 28203 29699 28209
rect 29641 28169 29653 28203
rect 29687 28200 29699 28203
rect 30190 28200 30196 28212
rect 29687 28172 30196 28200
rect 29687 28169 29699 28172
rect 29641 28163 29699 28169
rect 23109 28138 23244 28141
rect 23109 28135 23167 28138
rect 23109 28101 23121 28135
rect 23155 28101 23167 28135
rect 23109 28095 23167 28101
rect 24029 28135 24087 28141
rect 24029 28101 24041 28135
rect 24075 28132 24087 28135
rect 24578 28132 24584 28144
rect 24075 28104 24584 28132
rect 24075 28101 24087 28104
rect 24029 28095 24087 28101
rect 24578 28092 24584 28104
rect 24636 28092 24642 28144
rect 25130 28092 25136 28144
rect 25188 28132 25194 28144
rect 26510 28132 26516 28144
rect 25188 28104 26516 28132
rect 25188 28092 25194 28104
rect 13817 28067 13875 28073
rect 13817 28064 13829 28067
rect 13648 28036 13829 28064
rect 13817 28033 13829 28036
rect 13863 28033 13875 28067
rect 14274 28064 14280 28076
rect 14235 28036 14280 28064
rect 13817 28027 13875 28033
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 15013 28067 15071 28073
rect 15013 28033 15025 28067
rect 15059 28033 15071 28067
rect 15013 28027 15071 28033
rect 15197 28067 15255 28073
rect 15197 28033 15209 28067
rect 15243 28064 15255 28067
rect 17954 28064 17960 28076
rect 15243 28036 17960 28064
rect 15243 28033 15255 28036
rect 15197 28027 15255 28033
rect 8570 27996 8576 28008
rect 8531 27968 8576 27996
rect 8570 27956 8576 27968
rect 8628 27956 8634 28008
rect 8849 27999 8907 28005
rect 8849 27965 8861 27999
rect 8895 27965 8907 27999
rect 15028 27996 15056 28027
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 19886 28064 19892 28076
rect 19847 28036 19892 28064
rect 19886 28024 19892 28036
rect 19944 28064 19950 28076
rect 20717 28067 20775 28073
rect 20717 28064 20729 28067
rect 19944 28036 20729 28064
rect 19944 28024 19950 28036
rect 20717 28033 20729 28036
rect 20763 28033 20775 28067
rect 20717 28027 20775 28033
rect 20806 28024 20812 28076
rect 20864 28064 20870 28076
rect 22186 28064 22192 28076
rect 20864 28036 22192 28064
rect 20864 28024 20870 28036
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22554 28064 22560 28076
rect 22515 28036 22560 28064
rect 22554 28024 22560 28036
rect 22612 28024 22618 28076
rect 22649 28067 22707 28073
rect 22649 28033 22661 28067
rect 22695 28064 22707 28067
rect 22922 28064 22928 28076
rect 22695 28036 22928 28064
rect 22695 28033 22707 28036
rect 22649 28027 22707 28033
rect 22922 28024 22928 28036
rect 22980 28064 22986 28076
rect 23385 28067 23443 28073
rect 23385 28064 23397 28067
rect 22980 28036 23397 28064
rect 22980 28024 22986 28036
rect 23385 28033 23397 28036
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28064 24363 28067
rect 25222 28064 25228 28076
rect 24351 28036 25228 28064
rect 24351 28033 24363 28036
rect 24305 28027 24363 28033
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25424 28073 25452 28104
rect 26510 28092 26516 28104
rect 26568 28092 26574 28144
rect 28644 28132 28672 28163
rect 30190 28160 30196 28172
rect 30248 28160 30254 28212
rect 30300 28144 30604 28161
rect 28644 28104 29960 28132
rect 25409 28067 25467 28073
rect 25409 28033 25421 28067
rect 25455 28033 25467 28067
rect 25685 28067 25743 28073
rect 25685 28064 25697 28067
rect 25409 28027 25467 28033
rect 25516 28036 25697 28064
rect 23198 27996 23204 28008
rect 8849 27959 8907 27965
rect 13556 27968 15056 27996
rect 23159 27968 23204 27996
rect 3970 27888 3976 27940
rect 4028 27928 4034 27940
rect 8864 27928 8892 27959
rect 13556 27937 13584 27968
rect 23198 27956 23204 27968
rect 23256 27956 23262 28008
rect 24213 27999 24271 28005
rect 24213 27965 24225 27999
rect 24259 27996 24271 27999
rect 24486 27996 24492 28008
rect 24259 27968 24492 27996
rect 24259 27965 24271 27968
rect 24213 27959 24271 27965
rect 24486 27956 24492 27968
rect 24544 27956 24550 28008
rect 4028 27900 8892 27928
rect 13541 27931 13599 27937
rect 4028 27888 4034 27900
rect 13541 27897 13553 27931
rect 13587 27897 13599 27931
rect 13541 27891 13599 27897
rect 14461 27931 14519 27937
rect 14461 27897 14473 27931
rect 14507 27928 14519 27931
rect 14550 27928 14556 27940
rect 14507 27900 14556 27928
rect 14507 27897 14519 27900
rect 14461 27891 14519 27897
rect 14550 27888 14556 27900
rect 14608 27928 14614 27940
rect 15102 27928 15108 27940
rect 14608 27900 15108 27928
rect 14608 27888 14614 27900
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 22830 27888 22836 27940
rect 22888 27928 22894 27940
rect 23569 27931 23627 27937
rect 23569 27928 23581 27931
rect 22888 27900 23581 27928
rect 22888 27888 22894 27900
rect 23569 27897 23581 27900
rect 23615 27897 23627 27931
rect 24670 27928 24676 27940
rect 23569 27891 23627 27897
rect 24320 27900 24676 27928
rect 15010 27860 15016 27872
rect 14971 27832 15016 27860
rect 15010 27820 15016 27832
rect 15068 27820 15074 27872
rect 20714 27820 20720 27872
rect 20772 27860 20778 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 20772 27832 22017 27860
rect 20772 27820 20778 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 22554 27820 22560 27872
rect 22612 27860 22618 27872
rect 24320 27869 24348 27900
rect 24670 27888 24676 27900
rect 24728 27928 24734 27940
rect 25516 27928 25544 28036
rect 25685 28033 25697 28036
rect 25731 28033 25743 28067
rect 26326 28064 26332 28076
rect 26287 28036 26332 28064
rect 25685 28027 25743 28033
rect 26326 28024 26332 28036
rect 26384 28024 26390 28076
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 28350 28064 28356 28076
rect 27764 28036 28356 28064
rect 27764 28024 27770 28036
rect 28350 28024 28356 28036
rect 28408 28064 28414 28076
rect 28570 28067 28628 28073
rect 28570 28064 28582 28067
rect 28408 28036 28582 28064
rect 28408 28024 28414 28036
rect 28570 28033 28582 28036
rect 28616 28033 28628 28067
rect 29086 28064 29092 28076
rect 29047 28036 29092 28064
rect 28570 28027 28628 28033
rect 29086 28024 29092 28036
rect 29144 28024 29150 28076
rect 29546 28064 29552 28076
rect 29507 28036 29552 28064
rect 29546 28024 29552 28036
rect 29604 28024 29610 28076
rect 29932 28064 29960 28104
rect 30282 28092 30288 28144
rect 30340 28133 30604 28144
rect 30340 28092 30346 28133
rect 30576 28132 30604 28133
rect 30926 28132 30932 28144
rect 30576 28104 30696 28132
rect 30374 28064 30380 28076
rect 29932 28036 30380 28064
rect 30374 28024 30380 28036
rect 30432 28024 30438 28076
rect 30668 28073 30696 28104
rect 30852 28104 30932 28132
rect 30755 28089 30813 28095
rect 30469 28067 30527 28073
rect 30469 28033 30481 28067
rect 30515 28033 30527 28067
rect 30469 28027 30527 28033
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30755 28055 30767 28089
rect 30801 28086 30813 28089
rect 30852 28086 30880 28104
rect 30926 28092 30932 28104
rect 30984 28092 30990 28144
rect 36449 28135 36507 28141
rect 36449 28101 36461 28135
rect 36495 28132 36507 28135
rect 37461 28135 37519 28141
rect 37461 28132 37473 28135
rect 36495 28104 37473 28132
rect 36495 28101 36507 28104
rect 36449 28095 36507 28101
rect 37461 28101 37473 28104
rect 37507 28101 37519 28135
rect 37461 28095 37519 28101
rect 30801 28058 30880 28086
rect 31205 28067 31263 28073
rect 31205 28064 31217 28067
rect 30801 28055 30813 28058
rect 30755 28049 30813 28055
rect 30653 28027 30711 28033
rect 30944 28036 31217 28064
rect 28718 27956 28724 28008
rect 28776 27996 28782 28008
rect 28997 27999 29055 28005
rect 28997 27996 29009 27999
rect 28776 27968 29009 27996
rect 28776 27956 28782 27968
rect 28997 27965 29009 27968
rect 29043 27965 29055 27999
rect 28997 27959 29055 27965
rect 30190 27956 30196 28008
rect 30248 27996 30254 28008
rect 30484 27996 30512 28027
rect 30944 28008 30972 28036
rect 31205 28033 31217 28036
rect 31251 28033 31263 28067
rect 31386 28064 31392 28076
rect 31347 28036 31392 28064
rect 31205 28027 31263 28033
rect 31386 28024 31392 28036
rect 31444 28024 31450 28076
rect 32766 28064 32772 28076
rect 32727 28036 32772 28064
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 36354 28064 36360 28076
rect 36315 28036 36360 28064
rect 36354 28024 36360 28036
rect 36412 28024 36418 28076
rect 30248 27968 30512 27996
rect 30248 27956 30254 27968
rect 30926 27956 30932 28008
rect 30984 27956 30990 28008
rect 37274 27996 37280 28008
rect 37235 27968 37280 27996
rect 37274 27956 37280 27968
rect 37332 27956 37338 28008
rect 39117 27999 39175 28005
rect 39117 27965 39129 27999
rect 39163 27996 39175 27999
rect 46842 27996 46848 28008
rect 39163 27968 46848 27996
rect 39163 27965 39175 27968
rect 39117 27959 39175 27965
rect 46842 27956 46848 27968
rect 46900 27956 46906 28008
rect 24728 27900 25544 27928
rect 24728 27888 24734 27900
rect 26878 27888 26884 27940
rect 26936 27928 26942 27940
rect 32490 27928 32496 27940
rect 26936 27900 32496 27928
rect 26936 27888 26942 27900
rect 32490 27888 32496 27900
rect 32548 27928 32554 27940
rect 32674 27928 32680 27940
rect 32548 27900 32680 27928
rect 32548 27888 32554 27900
rect 32674 27888 32680 27900
rect 32732 27888 32738 27940
rect 23109 27863 23167 27869
rect 23109 27860 23121 27863
rect 22612 27832 23121 27860
rect 22612 27820 22618 27832
rect 23109 27829 23121 27832
rect 23155 27829 23167 27863
rect 23109 27823 23167 27829
rect 24305 27863 24363 27869
rect 24305 27829 24317 27863
rect 24351 27829 24363 27863
rect 24305 27823 24363 27829
rect 25038 27820 25044 27872
rect 25096 27860 25102 27872
rect 25317 27863 25375 27869
rect 25317 27860 25329 27863
rect 25096 27832 25329 27860
rect 25096 27820 25102 27832
rect 25317 27829 25329 27832
rect 25363 27829 25375 27863
rect 25317 27823 25375 27829
rect 25501 27863 25559 27869
rect 25501 27829 25513 27863
rect 25547 27860 25559 27863
rect 25590 27860 25596 27872
rect 25547 27832 25596 27860
rect 25547 27829 25559 27832
rect 25501 27823 25559 27829
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 26142 27860 26148 27872
rect 26103 27832 26148 27860
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 28166 27820 28172 27872
rect 28224 27860 28230 27872
rect 28445 27863 28503 27869
rect 28445 27860 28457 27863
rect 28224 27832 28457 27860
rect 28224 27820 28230 27832
rect 28445 27829 28457 27832
rect 28491 27829 28503 27863
rect 28445 27823 28503 27829
rect 30193 27863 30251 27869
rect 30193 27829 30205 27863
rect 30239 27860 30251 27863
rect 30926 27860 30932 27872
rect 30239 27832 30932 27860
rect 30239 27829 30251 27832
rect 30193 27823 30251 27829
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 31202 27860 31208 27872
rect 31163 27832 31208 27860
rect 31202 27820 31208 27832
rect 31260 27820 31266 27872
rect 31294 27820 31300 27872
rect 31352 27860 31358 27872
rect 31573 27863 31631 27869
rect 31573 27860 31585 27863
rect 31352 27832 31585 27860
rect 31352 27820 31358 27832
rect 31573 27829 31585 27832
rect 31619 27829 31631 27863
rect 31573 27823 31631 27829
rect 32861 27863 32919 27869
rect 32861 27829 32873 27863
rect 32907 27860 32919 27863
rect 33134 27860 33140 27872
rect 32907 27832 33140 27860
rect 32907 27829 32919 27832
rect 32861 27823 32919 27829
rect 33134 27820 33140 27832
rect 33192 27820 33198 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 8297 27659 8355 27665
rect 8297 27625 8309 27659
rect 8343 27656 8355 27659
rect 8570 27656 8576 27668
rect 8343 27628 8576 27656
rect 8343 27625 8355 27628
rect 8297 27619 8355 27625
rect 8570 27616 8576 27628
rect 8628 27616 8634 27668
rect 14908 27659 14966 27665
rect 14908 27625 14920 27659
rect 14954 27656 14966 27659
rect 15010 27656 15016 27668
rect 14954 27628 15016 27656
rect 14954 27625 14966 27628
rect 14908 27619 14966 27625
rect 15010 27616 15016 27628
rect 15068 27616 15074 27668
rect 15102 27616 15108 27668
rect 15160 27656 15166 27668
rect 23566 27656 23572 27668
rect 15160 27628 23572 27656
rect 15160 27616 15166 27628
rect 23566 27616 23572 27628
rect 23624 27616 23630 27668
rect 25672 27659 25730 27665
rect 25672 27625 25684 27659
rect 25718 27656 25730 27659
rect 26142 27656 26148 27668
rect 25718 27628 26148 27656
rect 25718 27625 25730 27628
rect 25672 27619 25730 27625
rect 26142 27616 26148 27628
rect 26200 27616 26206 27668
rect 30374 27656 30380 27668
rect 30335 27628 30380 27656
rect 30374 27616 30380 27628
rect 30432 27616 30438 27668
rect 37274 27656 37280 27668
rect 37235 27628 37280 27656
rect 37274 27616 37280 27628
rect 37332 27616 37338 27668
rect 20346 27588 20352 27600
rect 8220 27560 12434 27588
rect 8220 27464 8248 27560
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 9401 27523 9459 27529
rect 9401 27520 9413 27523
rect 8444 27492 9413 27520
rect 8444 27480 8450 27492
rect 9401 27489 9413 27492
rect 9447 27489 9459 27523
rect 9401 27483 9459 27489
rect 8202 27452 8208 27464
rect 8115 27424 8208 27452
rect 8202 27412 8208 27424
rect 8260 27412 8266 27464
rect 8941 27455 8999 27461
rect 8941 27421 8953 27455
rect 8987 27421 8999 27455
rect 12406 27452 12434 27560
rect 19536 27560 20352 27588
rect 14642 27452 14648 27464
rect 12406 27424 14504 27452
rect 14603 27424 14648 27452
rect 8941 27415 8999 27421
rect 8956 27316 8984 27415
rect 9122 27384 9128 27396
rect 9083 27356 9128 27384
rect 9122 27344 9128 27356
rect 9180 27344 9186 27396
rect 13354 27384 13360 27396
rect 13315 27356 13360 27384
rect 13354 27344 13360 27356
rect 13412 27344 13418 27396
rect 14476 27384 14504 27424
rect 14642 27412 14648 27424
rect 14700 27412 14706 27464
rect 16206 27412 16212 27464
rect 16264 27452 16270 27464
rect 19536 27461 19564 27560
rect 20346 27548 20352 27560
rect 20404 27548 20410 27600
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 22186 27588 22192 27600
rect 21775 27560 22192 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 22186 27548 22192 27560
rect 22244 27548 22250 27600
rect 24397 27591 24455 27597
rect 24397 27557 24409 27591
rect 24443 27588 24455 27591
rect 25406 27588 25412 27600
rect 24443 27560 25412 27588
rect 24443 27557 24455 27560
rect 24397 27551 24455 27557
rect 25406 27548 25412 27560
rect 25464 27548 25470 27600
rect 28258 27548 28264 27600
rect 28316 27588 28322 27600
rect 28316 27560 28488 27588
rect 28316 27548 28322 27560
rect 20714 27520 20720 27532
rect 19720 27492 20720 27520
rect 19720 27461 19748 27492
rect 20714 27480 20720 27492
rect 20772 27480 20778 27532
rect 23201 27523 23259 27529
rect 23201 27489 23213 27523
rect 23247 27520 23259 27523
rect 23474 27520 23480 27532
rect 23247 27492 23480 27520
rect 23247 27489 23259 27492
rect 23201 27483 23259 27489
rect 23474 27480 23480 27492
rect 23532 27520 23538 27532
rect 24578 27520 24584 27532
rect 23532 27492 24584 27520
rect 23532 27480 23538 27492
rect 24578 27480 24584 27492
rect 24636 27520 24642 27532
rect 27157 27523 27215 27529
rect 27157 27520 27169 27523
rect 24636 27492 27169 27520
rect 24636 27480 24642 27492
rect 27157 27489 27169 27492
rect 27203 27489 27215 27523
rect 27157 27483 27215 27489
rect 27706 27480 27712 27532
rect 27764 27520 27770 27532
rect 28353 27523 28411 27529
rect 28353 27520 28365 27523
rect 27764 27492 28365 27520
rect 27764 27480 27770 27492
rect 28353 27489 28365 27492
rect 28399 27489 28411 27523
rect 28353 27483 28411 27489
rect 16853 27455 16911 27461
rect 16853 27452 16865 27455
rect 16264 27424 16865 27452
rect 16264 27412 16270 27424
rect 16853 27421 16865 27424
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 20990 27452 20996 27464
rect 19935 27424 20392 27452
rect 20951 27424 20996 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 15194 27384 15200 27396
rect 14476 27356 15200 27384
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 16666 27384 16672 27396
rect 16146 27356 16672 27384
rect 16666 27344 16672 27356
rect 16724 27344 16730 27396
rect 17037 27387 17095 27393
rect 17037 27353 17049 27387
rect 17083 27384 17095 27387
rect 17126 27384 17132 27396
rect 17083 27356 17132 27384
rect 17083 27353 17095 27356
rect 17037 27347 17095 27353
rect 17126 27344 17132 27356
rect 17184 27344 17190 27396
rect 18690 27384 18696 27396
rect 18651 27356 18696 27384
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 19628 27384 19656 27415
rect 20070 27384 20076 27396
rect 19628 27356 20076 27384
rect 20070 27344 20076 27356
rect 20128 27344 20134 27396
rect 9674 27316 9680 27328
rect 8956 27288 9680 27316
rect 9674 27276 9680 27288
rect 9732 27276 9738 27328
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 13446 27316 13452 27328
rect 12768 27288 13452 27316
rect 12768 27276 12774 27288
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 13538 27276 13544 27328
rect 13596 27316 13602 27328
rect 13722 27316 13728 27328
rect 13596 27288 13728 27316
rect 13596 27276 13602 27288
rect 13722 27276 13728 27288
rect 13780 27316 13786 27328
rect 16393 27319 16451 27325
rect 16393 27316 16405 27319
rect 13780 27288 16405 27316
rect 13780 27276 13786 27288
rect 16393 27285 16405 27288
rect 16439 27285 16451 27319
rect 16393 27279 16451 27285
rect 18874 27276 18880 27328
rect 18932 27316 18938 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 18932 27288 19257 27316
rect 18932 27276 18938 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 20364 27316 20392 27424
rect 20990 27412 20996 27424
rect 21048 27412 21054 27464
rect 21729 27455 21787 27461
rect 21085 27433 21143 27439
rect 21085 27399 21097 27433
rect 21131 27418 21143 27433
rect 21729 27421 21741 27455
rect 21775 27421 21787 27455
rect 21910 27452 21916 27464
rect 21871 27424 21916 27452
rect 21131 27399 21220 27418
rect 21729 27415 21787 27421
rect 21085 27396 21220 27399
rect 20806 27384 20812 27396
rect 20767 27356 20812 27384
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 21085 27393 21180 27396
rect 21100 27390 21180 27393
rect 21174 27344 21180 27390
rect 21232 27344 21238 27396
rect 21744 27384 21772 27415
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22922 27452 22928 27464
rect 22883 27424 22928 27452
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 23072 27424 23117 27452
rect 23216 27424 24685 27452
rect 23072 27412 23078 27424
rect 22094 27384 22100 27396
rect 21744 27356 22100 27384
rect 22094 27344 22100 27356
rect 22152 27344 22158 27396
rect 23216 27393 23244 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 25314 27412 25320 27464
rect 25372 27452 25378 27464
rect 25409 27455 25467 27461
rect 25409 27452 25421 27455
rect 25372 27424 25421 27452
rect 25372 27412 25378 27424
rect 25409 27421 25421 27424
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 28077 27455 28135 27461
rect 28077 27421 28089 27455
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 23201 27387 23259 27393
rect 23201 27353 23213 27387
rect 23247 27353 23259 27387
rect 24394 27384 24400 27396
rect 24355 27356 24400 27384
rect 23201 27347 23259 27353
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 24581 27387 24639 27393
rect 24581 27353 24593 27387
rect 24627 27384 24639 27387
rect 25038 27384 25044 27396
rect 24627 27356 25044 27384
rect 24627 27353 24639 27356
rect 24581 27347 24639 27353
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 27062 27384 27068 27396
rect 26910 27356 27068 27384
rect 27062 27344 27068 27356
rect 27120 27344 27126 27396
rect 28092 27384 28120 27415
rect 28166 27412 28172 27464
rect 28224 27452 28230 27464
rect 28460 27461 28488 27560
rect 32122 27480 32128 27532
rect 32180 27520 32186 27532
rect 32217 27523 32275 27529
rect 32217 27520 32229 27523
rect 32180 27492 32229 27520
rect 32180 27480 32186 27492
rect 32217 27489 32229 27492
rect 32263 27520 32275 27523
rect 32582 27520 32588 27532
rect 32263 27492 32588 27520
rect 32263 27489 32275 27492
rect 32217 27483 32275 27489
rect 32582 27480 32588 27492
rect 32640 27480 32646 27532
rect 28445 27455 28503 27461
rect 28224 27424 28269 27452
rect 28224 27412 28230 27424
rect 28445 27421 28457 27455
rect 28491 27421 28503 27455
rect 28445 27415 28503 27421
rect 29638 27412 29644 27464
rect 29696 27452 29702 27464
rect 30193 27455 30251 27461
rect 30193 27452 30205 27455
rect 29696 27424 30205 27452
rect 29696 27412 29702 27424
rect 30193 27421 30205 27424
rect 30239 27421 30251 27455
rect 30193 27415 30251 27421
rect 29914 27384 29920 27396
rect 28092 27356 29920 27384
rect 29914 27344 29920 27356
rect 29972 27344 29978 27396
rect 30006 27344 30012 27396
rect 30064 27384 30070 27396
rect 31294 27384 31300 27396
rect 30064 27356 31300 27384
rect 30064 27344 30070 27356
rect 31294 27344 31300 27356
rect 31352 27344 31358 27396
rect 32490 27384 32496 27396
rect 32451 27356 32496 27384
rect 32490 27344 32496 27356
rect 32548 27344 32554 27396
rect 33134 27344 33140 27396
rect 33192 27344 33198 27396
rect 20901 27319 20959 27325
rect 20901 27316 20913 27319
rect 20364 27288 20913 27316
rect 19245 27279 19303 27285
rect 20901 27285 20913 27288
rect 20947 27285 20959 27319
rect 20901 27279 20959 27285
rect 27893 27319 27951 27325
rect 27893 27285 27905 27319
rect 27939 27316 27951 27319
rect 28166 27316 28172 27328
rect 27939 27288 28172 27316
rect 27939 27285 27951 27288
rect 27893 27279 27951 27285
rect 28166 27276 28172 27288
rect 28224 27276 28230 27328
rect 30190 27276 30196 27328
rect 30248 27316 30254 27328
rect 32398 27316 32404 27328
rect 30248 27288 32404 27316
rect 30248 27276 30254 27288
rect 32398 27276 32404 27288
rect 32456 27316 32462 27328
rect 33965 27319 34023 27325
rect 33965 27316 33977 27319
rect 32456 27288 33977 27316
rect 32456 27276 32462 27288
rect 33965 27285 33977 27288
rect 34011 27285 34023 27319
rect 33965 27279 34023 27285
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 8297 27115 8355 27121
rect 8297 27081 8309 27115
rect 8343 27112 8355 27115
rect 9122 27112 9128 27124
rect 8343 27084 9128 27112
rect 8343 27081 8355 27084
rect 8297 27075 8355 27081
rect 9122 27072 9128 27084
rect 9180 27072 9186 27124
rect 14182 27072 14188 27124
rect 14240 27112 14246 27124
rect 14277 27115 14335 27121
rect 14277 27112 14289 27115
rect 14240 27084 14289 27112
rect 14240 27072 14246 27084
rect 14277 27081 14289 27084
rect 14323 27081 14335 27115
rect 14458 27112 14464 27124
rect 14419 27084 14464 27112
rect 14277 27075 14335 27081
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 14642 27072 14648 27124
rect 14700 27112 14706 27124
rect 15933 27115 15991 27121
rect 15933 27112 15945 27115
rect 14700 27084 15945 27112
rect 14700 27072 14706 27084
rect 15933 27081 15945 27084
rect 15979 27081 15991 27115
rect 17126 27112 17132 27124
rect 17087 27084 17132 27112
rect 15933 27075 15991 27081
rect 17126 27072 17132 27084
rect 17184 27072 17190 27124
rect 18690 27072 18696 27124
rect 18748 27112 18754 27124
rect 46566 27112 46572 27124
rect 18748 27084 46572 27112
rect 18748 27072 18754 27084
rect 46566 27072 46572 27084
rect 46624 27072 46630 27124
rect 12434 27004 12440 27056
rect 12492 27004 12498 27056
rect 13722 27004 13728 27056
rect 13780 27044 13786 27056
rect 13909 27047 13967 27053
rect 13909 27044 13921 27047
rect 13780 27016 13921 27044
rect 13780 27004 13786 27016
rect 13909 27013 13921 27016
rect 13955 27013 13967 27047
rect 13909 27007 13967 27013
rect 14366 27004 14372 27056
rect 14424 27044 14430 27056
rect 14921 27047 14979 27053
rect 14921 27044 14933 27047
rect 14424 27016 14933 27044
rect 14424 27004 14430 27016
rect 14921 27013 14933 27016
rect 14967 27013 14979 27047
rect 15121 27047 15179 27053
rect 15121 27044 15133 27047
rect 14921 27007 14979 27013
rect 15028 27016 15133 27044
rect 8202 26976 8208 26988
rect 8163 26948 8208 26976
rect 8202 26936 8208 26948
rect 8260 26936 8266 26988
rect 9033 26979 9091 26985
rect 9033 26945 9045 26979
rect 9079 26976 9091 26979
rect 10226 26976 10232 26988
rect 9079 26948 10232 26976
rect 9079 26945 9091 26948
rect 9033 26939 9091 26945
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14185 26979 14243 26985
rect 14185 26945 14197 26979
rect 14231 26976 14243 26979
rect 14734 26976 14740 26988
rect 14231 26948 14740 26976
rect 14231 26945 14243 26948
rect 14185 26939 14243 26945
rect 11514 26908 11520 26920
rect 11475 26880 11520 26908
rect 11514 26868 11520 26880
rect 11572 26868 11578 26920
rect 11790 26908 11796 26920
rect 11751 26880 11796 26908
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 13722 26868 13728 26920
rect 13780 26908 13786 26920
rect 14108 26908 14136 26939
rect 14734 26936 14740 26948
rect 14792 26976 14798 26988
rect 15028 26976 15056 27016
rect 15121 27013 15133 27016
rect 15167 27013 15179 27047
rect 15121 27007 15179 27013
rect 15286 27004 15292 27056
rect 15344 27044 15350 27056
rect 18874 27044 18880 27056
rect 15344 27016 16988 27044
rect 18835 27016 18880 27044
rect 15344 27004 15350 27016
rect 16960 26988 16988 27016
rect 18874 27004 18880 27016
rect 18932 27004 18938 27056
rect 19886 27004 19892 27056
rect 19944 27004 19950 27056
rect 21910 27044 21916 27056
rect 21823 27016 21916 27044
rect 21910 27004 21916 27016
rect 21968 27044 21974 27056
rect 22281 27047 22339 27053
rect 22281 27044 22293 27047
rect 21968 27016 22293 27044
rect 21968 27004 21974 27016
rect 22281 27013 22293 27016
rect 22327 27013 22339 27047
rect 22281 27007 22339 27013
rect 22465 27047 22523 27053
rect 22465 27013 22477 27047
rect 22511 27044 22523 27047
rect 23014 27044 23020 27056
rect 22511 27016 23020 27044
rect 22511 27013 22523 27016
rect 22465 27007 22523 27013
rect 23014 27004 23020 27016
rect 23072 27004 23078 27056
rect 27062 27044 27068 27056
rect 27023 27016 27068 27044
rect 27062 27004 27068 27016
rect 27120 27004 27126 27056
rect 28166 27044 28172 27056
rect 28127 27016 28172 27044
rect 28166 27004 28172 27016
rect 28224 27004 28230 27056
rect 29638 27044 29644 27056
rect 29394 27016 29644 27044
rect 29638 27004 29644 27016
rect 29696 27004 29702 27056
rect 32490 27004 32496 27056
rect 32548 27044 32554 27056
rect 32861 27047 32919 27053
rect 32861 27044 32873 27047
rect 32548 27016 32873 27044
rect 32548 27004 32554 27016
rect 32861 27013 32873 27016
rect 32907 27013 32919 27047
rect 32861 27007 32919 27013
rect 14792 26948 15056 26976
rect 14792 26936 14798 26948
rect 15378 26936 15384 26988
rect 15436 26976 15442 26988
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15436 26948 15761 26976
rect 15436 26936 15442 26948
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 16942 26936 16948 26988
rect 17000 26976 17006 26988
rect 17037 26979 17095 26985
rect 17037 26976 17049 26979
rect 17000 26948 17049 26976
rect 17000 26936 17006 26948
rect 17037 26945 17049 26948
rect 17083 26945 17095 26979
rect 17037 26939 17095 26945
rect 13780 26880 14136 26908
rect 18601 26911 18659 26917
rect 13780 26868 13786 26880
rect 18601 26877 18613 26911
rect 18647 26877 18659 26911
rect 18601 26871 18659 26877
rect 13354 26800 13360 26852
rect 13412 26840 13418 26852
rect 15289 26843 15347 26849
rect 15289 26840 15301 26843
rect 13412 26812 15301 26840
rect 13412 26800 13418 26812
rect 15289 26809 15301 26812
rect 15335 26809 15347 26843
rect 15289 26803 15347 26809
rect 8849 26775 8907 26781
rect 8849 26741 8861 26775
rect 8895 26772 8907 26775
rect 8938 26772 8944 26784
rect 8895 26744 8944 26772
rect 8895 26741 8907 26744
rect 8849 26735 8907 26741
rect 8938 26732 8944 26744
rect 8996 26732 9002 26784
rect 13170 26732 13176 26784
rect 13228 26772 13234 26784
rect 13265 26775 13323 26781
rect 13265 26772 13277 26775
rect 13228 26744 13277 26772
rect 13228 26732 13234 26744
rect 13265 26741 13277 26744
rect 13311 26741 13323 26775
rect 13265 26735 13323 26741
rect 13722 26732 13728 26784
rect 13780 26772 13786 26784
rect 15105 26775 15163 26781
rect 15105 26772 15117 26775
rect 13780 26744 15117 26772
rect 13780 26732 13786 26744
rect 15105 26741 15117 26744
rect 15151 26741 15163 26775
rect 18616 26772 18644 26871
rect 21542 26868 21548 26920
rect 21600 26908 21606 26920
rect 21928 26908 21956 27004
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22152 26948 22937 26976
rect 22152 26936 22158 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26976 23259 26979
rect 23474 26976 23480 26988
rect 23247 26948 23480 26976
rect 23247 26945 23259 26948
rect 23201 26939 23259 26945
rect 23474 26936 23480 26948
rect 23532 26936 23538 26988
rect 26970 26976 26976 26988
rect 26931 26948 26976 26976
rect 26970 26936 26976 26948
rect 27028 26936 27034 26988
rect 30926 26936 30932 26988
rect 30984 26976 30990 26988
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 30984 26948 32137 26976
rect 30984 26936 30990 26948
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32306 26976 32312 26988
rect 32267 26948 32312 26976
rect 32125 26939 32183 26945
rect 32306 26936 32312 26948
rect 32364 26936 32370 26988
rect 32398 26936 32404 26988
rect 32456 26976 32462 26988
rect 32674 26976 32680 26988
rect 32456 26948 32501 26976
rect 32635 26948 32680 26976
rect 32456 26936 32462 26948
rect 32674 26936 32680 26948
rect 32732 26936 32738 26988
rect 22830 26908 22836 26920
rect 21600 26880 22836 26908
rect 21600 26868 21606 26880
rect 22830 26868 22836 26880
rect 22888 26908 22894 26920
rect 23017 26911 23075 26917
rect 23017 26908 23029 26911
rect 22888 26880 23029 26908
rect 22888 26868 22894 26880
rect 23017 26877 23029 26880
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 27890 26908 27896 26920
rect 25372 26880 27896 26908
rect 25372 26868 25378 26880
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 29641 26911 29699 26917
rect 29641 26877 29653 26911
rect 29687 26908 29699 26911
rect 29730 26908 29736 26920
rect 29687 26880 29736 26908
rect 29687 26877 29699 26880
rect 29641 26871 29699 26877
rect 29730 26868 29736 26880
rect 29788 26868 29794 26920
rect 32493 26911 32551 26917
rect 32493 26877 32505 26911
rect 32539 26908 32551 26911
rect 32582 26908 32588 26920
rect 32539 26880 32588 26908
rect 32539 26877 32551 26880
rect 32493 26871 32551 26877
rect 32582 26868 32588 26880
rect 32640 26868 32646 26920
rect 21634 26800 21640 26852
rect 21692 26840 21698 26852
rect 21818 26840 21824 26852
rect 21692 26812 21824 26840
rect 21692 26800 21698 26812
rect 21818 26800 21824 26812
rect 21876 26800 21882 26852
rect 23385 26843 23443 26849
rect 23385 26809 23397 26843
rect 23431 26840 23443 26843
rect 25038 26840 25044 26852
rect 23431 26812 25044 26840
rect 23431 26809 23443 26812
rect 23385 26803 23443 26809
rect 25038 26800 25044 26812
rect 25096 26800 25102 26852
rect 19334 26772 19340 26784
rect 18616 26744 19340 26772
rect 15105 26735 15163 26741
rect 19334 26732 19340 26744
rect 19392 26732 19398 26784
rect 20349 26775 20407 26781
rect 20349 26741 20361 26775
rect 20395 26772 20407 26775
rect 21174 26772 21180 26784
rect 20395 26744 21180 26772
rect 20395 26741 20407 26744
rect 20349 26735 20407 26741
rect 21174 26732 21180 26744
rect 21232 26772 21238 26784
rect 22922 26772 22928 26784
rect 21232 26744 22928 26772
rect 21232 26732 21238 26744
rect 22922 26732 22928 26744
rect 22980 26732 22986 26784
rect 24394 26732 24400 26784
rect 24452 26772 24458 26784
rect 30282 26772 30288 26784
rect 24452 26744 30288 26772
rect 24452 26732 24458 26744
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 2590 26528 2596 26580
rect 2648 26568 2654 26580
rect 11701 26571 11759 26577
rect 2648 26540 10272 26568
rect 2648 26528 2654 26540
rect 10244 26500 10272 26540
rect 11701 26537 11713 26571
rect 11747 26568 11759 26571
rect 11790 26568 11796 26580
rect 11747 26540 11796 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 11790 26528 11796 26540
rect 11848 26528 11854 26580
rect 27430 26568 27436 26580
rect 12406 26540 27436 26568
rect 12406 26500 12434 26540
rect 27430 26528 27436 26540
rect 27488 26528 27494 26580
rect 29638 26568 29644 26580
rect 27816 26540 28028 26568
rect 29599 26540 29644 26568
rect 10244 26472 12434 26500
rect 16117 26503 16175 26509
rect 16117 26469 16129 26503
rect 16163 26500 16175 26503
rect 16206 26500 16212 26512
rect 16163 26472 16212 26500
rect 16163 26469 16175 26472
rect 16117 26463 16175 26469
rect 8938 26432 8944 26444
rect 8899 26404 8944 26432
rect 8938 26392 8944 26404
rect 8996 26392 9002 26444
rect 11517 26435 11575 26441
rect 11517 26401 11529 26435
rect 11563 26432 11575 26435
rect 11606 26432 11612 26444
rect 11563 26404 11612 26432
rect 11563 26401 11575 26404
rect 11517 26395 11575 26401
rect 11606 26392 11612 26404
rect 11664 26392 11670 26444
rect 12713 26435 12771 26441
rect 12713 26401 12725 26435
rect 12759 26432 12771 26435
rect 13354 26432 13360 26444
rect 12759 26404 13360 26432
rect 12759 26401 12771 26404
rect 12713 26395 12771 26401
rect 13354 26392 13360 26404
rect 13412 26392 13418 26444
rect 14090 26392 14096 26444
rect 14148 26432 14154 26444
rect 16132 26432 16160 26463
rect 16206 26460 16212 26472
rect 16264 26460 16270 26512
rect 16666 26500 16672 26512
rect 16627 26472 16672 26500
rect 16666 26460 16672 26472
rect 16724 26460 16730 26512
rect 19886 26500 19892 26512
rect 19847 26472 19892 26500
rect 19886 26460 19892 26472
rect 19944 26460 19950 26512
rect 21450 26460 21456 26512
rect 21508 26500 21514 26512
rect 21729 26503 21787 26509
rect 21729 26500 21741 26503
rect 21508 26472 21741 26500
rect 21508 26460 21514 26472
rect 21729 26469 21741 26472
rect 21775 26469 21787 26503
rect 21729 26463 21787 26469
rect 21818 26460 21824 26512
rect 21876 26500 21882 26512
rect 27816 26500 27844 26540
rect 21876 26472 27844 26500
rect 27893 26503 27951 26509
rect 21876 26460 21882 26472
rect 27893 26469 27905 26503
rect 27939 26469 27951 26503
rect 28000 26500 28028 26540
rect 29638 26528 29644 26540
rect 29696 26528 29702 26580
rect 30377 26571 30435 26577
rect 30377 26537 30389 26571
rect 30423 26568 30435 26571
rect 30466 26568 30472 26580
rect 30423 26540 30472 26568
rect 30423 26537 30435 26540
rect 30377 26531 30435 26537
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 31110 26568 31116 26580
rect 31071 26540 31116 26568
rect 31110 26528 31116 26540
rect 31168 26528 31174 26580
rect 31128 26500 31156 26528
rect 32306 26500 32312 26512
rect 28000 26472 31156 26500
rect 31956 26472 32312 26500
rect 27893 26463 27951 26469
rect 14148 26404 16160 26432
rect 21177 26435 21235 26441
rect 14148 26392 14154 26404
rect 21177 26401 21189 26435
rect 21223 26432 21235 26435
rect 22554 26432 22560 26444
rect 21223 26404 22048 26432
rect 22515 26404 22560 26432
rect 21223 26401 21235 26404
rect 21177 26395 21235 26401
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26364 11483 26367
rect 12618 26364 12624 26376
rect 11471 26336 12624 26364
rect 11471 26333 11483 26336
rect 11425 26327 11483 26333
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 12986 26364 12992 26376
rect 12947 26336 12992 26364
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 14366 26364 14372 26376
rect 14327 26336 14372 26364
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 15746 26324 15752 26376
rect 15804 26324 15810 26376
rect 16574 26364 16580 26376
rect 16535 26336 16580 26364
rect 16574 26324 16580 26336
rect 16632 26324 16638 26376
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 19978 26364 19984 26376
rect 19843 26336 19984 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21542 26364 21548 26376
rect 21315 26336 21548 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 9214 26296 9220 26308
rect 9175 26268 9220 26296
rect 9214 26256 9220 26268
rect 9272 26256 9278 26308
rect 9950 26256 9956 26308
rect 10008 26256 10014 26308
rect 14642 26296 14648 26308
rect 14603 26268 14648 26296
rect 14642 26256 14648 26268
rect 14700 26256 14706 26308
rect 21100 26296 21128 26327
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 21729 26367 21787 26373
rect 21729 26333 21741 26367
rect 21775 26364 21787 26367
rect 21818 26364 21824 26376
rect 21775 26336 21824 26364
rect 21775 26333 21787 26336
rect 21729 26327 21787 26333
rect 21818 26324 21824 26336
rect 21876 26324 21882 26376
rect 22020 26373 22048 26404
rect 22554 26392 22560 26404
rect 22612 26392 22618 26444
rect 22830 26432 22836 26444
rect 22791 26404 22836 26432
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 24486 26392 24492 26444
rect 24544 26432 24550 26444
rect 24581 26435 24639 26441
rect 24581 26432 24593 26435
rect 24544 26404 24593 26432
rect 24544 26392 24550 26404
rect 24581 26401 24593 26404
rect 24627 26432 24639 26435
rect 27908 26432 27936 26463
rect 24627 26404 25636 26432
rect 24627 26401 24639 26404
rect 24581 26395 24639 26401
rect 25608 26376 25636 26404
rect 27172 26404 27936 26432
rect 22005 26367 22063 26373
rect 22005 26333 22017 26367
rect 22051 26333 22063 26367
rect 22005 26327 22063 26333
rect 24765 26367 24823 26373
rect 24765 26333 24777 26367
rect 24811 26364 24823 26367
rect 25038 26364 25044 26376
rect 24811 26336 25044 26364
rect 24811 26333 24823 26336
rect 24765 26327 24823 26333
rect 25038 26324 25044 26336
rect 25096 26364 25102 26376
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 25096 26336 25421 26364
rect 25096 26324 25102 26336
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 27062 26364 27068 26376
rect 25648 26336 27068 26364
rect 25648 26324 25654 26336
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 27172 26373 27200 26404
rect 28074 26392 28080 26444
rect 28132 26432 28138 26444
rect 28353 26435 28411 26441
rect 28353 26432 28365 26435
rect 28132 26404 28365 26432
rect 28132 26392 28138 26404
rect 28353 26401 28365 26404
rect 28399 26401 28411 26435
rect 28353 26395 28411 26401
rect 28537 26435 28595 26441
rect 28537 26401 28549 26435
rect 28583 26432 28595 26435
rect 29454 26432 29460 26444
rect 28583 26404 29460 26432
rect 28583 26401 28595 26404
rect 28537 26395 28595 26401
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27338 26364 27344 26376
rect 27299 26336 27344 26364
rect 27157 26327 27215 26333
rect 27338 26324 27344 26336
rect 27396 26324 27402 26376
rect 27430 26324 27436 26376
rect 27488 26364 27494 26376
rect 27488 26336 27533 26364
rect 27488 26324 27494 26336
rect 21913 26299 21971 26305
rect 21100 26268 21680 26296
rect 8478 26188 8484 26240
rect 8536 26228 8542 26240
rect 10689 26231 10747 26237
rect 10689 26228 10701 26231
rect 8536 26200 10701 26228
rect 8536 26188 8542 26200
rect 10689 26197 10701 26200
rect 10735 26228 10747 26231
rect 11790 26228 11796 26240
rect 10735 26200 11796 26228
rect 10735 26197 10747 26200
rect 10689 26191 10747 26197
rect 11790 26188 11796 26200
rect 11848 26188 11854 26240
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 14090 26228 14096 26240
rect 12584 26200 14096 26228
rect 12584 26188 12590 26200
rect 14090 26188 14096 26200
rect 14148 26188 14154 26240
rect 21652 26228 21680 26268
rect 21913 26265 21925 26299
rect 21959 26296 21971 26299
rect 23014 26296 23020 26308
rect 21959 26268 23020 26296
rect 21959 26265 21971 26268
rect 21913 26259 21971 26265
rect 23014 26256 23020 26268
rect 23072 26256 23078 26308
rect 26973 26299 27031 26305
rect 26973 26265 26985 26299
rect 27019 26296 27031 26299
rect 27246 26296 27252 26308
rect 27019 26268 27252 26296
rect 27019 26265 27031 26268
rect 26973 26259 27031 26265
rect 27246 26256 27252 26268
rect 27304 26256 27310 26308
rect 28258 26296 28264 26308
rect 28219 26268 28264 26296
rect 28258 26256 28264 26268
rect 28316 26256 28322 26308
rect 28368 26296 28396 26395
rect 29454 26392 29460 26404
rect 29512 26392 29518 26444
rect 29546 26364 29552 26376
rect 29507 26336 29552 26364
rect 29546 26324 29552 26336
rect 29604 26324 29610 26376
rect 30193 26367 30251 26373
rect 30193 26333 30205 26367
rect 30239 26333 30251 26367
rect 30193 26327 30251 26333
rect 30208 26296 30236 26327
rect 30558 26324 30564 26376
rect 30616 26364 30622 26376
rect 30929 26367 30987 26373
rect 30929 26364 30941 26367
rect 30616 26336 30941 26364
rect 30616 26324 30622 26336
rect 30929 26333 30941 26336
rect 30975 26333 30987 26367
rect 31754 26364 31760 26376
rect 31715 26336 31760 26364
rect 30929 26327 30987 26333
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 31956 26373 31984 26472
rect 32306 26460 32312 26472
rect 32364 26460 32370 26512
rect 32125 26435 32183 26441
rect 32125 26401 32137 26435
rect 32171 26432 32183 26435
rect 40402 26432 40408 26444
rect 32171 26404 40408 26432
rect 32171 26401 32183 26404
rect 32125 26395 32183 26401
rect 40402 26392 40408 26404
rect 40460 26392 40466 26444
rect 31941 26367 31999 26373
rect 31941 26333 31953 26367
rect 31987 26333 31999 26367
rect 32033 26367 32091 26373
rect 32033 26354 32045 26367
rect 32079 26354 32091 26367
rect 32309 26367 32367 26373
rect 31941 26327 31999 26333
rect 32030 26302 32036 26354
rect 32088 26302 32094 26354
rect 32309 26333 32321 26367
rect 32355 26364 32367 26367
rect 32674 26364 32680 26376
rect 32355 26336 32680 26364
rect 32355 26333 32367 26336
rect 32309 26327 32367 26333
rect 32674 26324 32680 26336
rect 32732 26324 32738 26376
rect 28368 26268 30236 26296
rect 22094 26228 22100 26240
rect 21652 26200 22100 26228
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 24949 26231 25007 26237
rect 24949 26197 24961 26231
rect 24995 26228 25007 26231
rect 25406 26228 25412 26240
rect 24995 26200 25412 26228
rect 24995 26197 25007 26200
rect 24949 26191 25007 26197
rect 25406 26188 25412 26200
rect 25464 26188 25470 26240
rect 25501 26231 25559 26237
rect 25501 26197 25513 26231
rect 25547 26228 25559 26231
rect 25958 26228 25964 26240
rect 25547 26200 25964 26228
rect 25547 26197 25559 26200
rect 25501 26191 25559 26197
rect 25958 26188 25964 26200
rect 26016 26188 26022 26240
rect 32490 26228 32496 26240
rect 32451 26200 32496 26228
rect 32490 26188 32496 26200
rect 32548 26188 32554 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 8849 26027 8907 26033
rect 8849 25993 8861 26027
rect 8895 26024 8907 26027
rect 9214 26024 9220 26036
rect 8895 25996 9220 26024
rect 8895 25993 8907 25996
rect 8849 25987 8907 25993
rect 9214 25984 9220 25996
rect 9272 25984 9278 26036
rect 9950 25984 9956 26036
rect 10008 26024 10014 26036
rect 10045 26027 10103 26033
rect 10045 26024 10057 26027
rect 10008 25996 10057 26024
rect 10008 25984 10014 25996
rect 10045 25993 10057 25996
rect 10091 25993 10103 26027
rect 11606 26024 11612 26036
rect 11567 25996 11612 26024
rect 10045 25987 10103 25993
rect 11606 25984 11612 25996
rect 11664 25984 11670 26036
rect 11790 25984 11796 26036
rect 11848 26024 11854 26036
rect 12805 26027 12863 26033
rect 12805 26024 12817 26027
rect 11848 25996 12817 26024
rect 11848 25984 11854 25996
rect 12805 25993 12817 25996
rect 12851 26024 12863 26027
rect 13725 26027 13783 26033
rect 13725 26024 13737 26027
rect 12851 25996 13737 26024
rect 12851 25993 12863 25996
rect 12805 25987 12863 25993
rect 13725 25993 13737 25996
rect 13771 25993 13783 26027
rect 13725 25987 13783 25993
rect 13814 25984 13820 26036
rect 13872 26024 13878 26036
rect 14001 26027 14059 26033
rect 13872 25996 13917 26024
rect 13872 25984 13878 25996
rect 14001 25993 14013 26027
rect 14047 26024 14059 26027
rect 14182 26024 14188 26036
rect 14047 25996 14188 26024
rect 14047 25993 14059 25996
rect 14001 25987 14059 25993
rect 14182 25984 14188 25996
rect 14240 26024 14246 26036
rect 14240 25996 14596 26024
rect 14240 25984 14246 25996
rect 11698 25956 11704 25968
rect 11611 25928 11704 25956
rect 11698 25916 11704 25928
rect 11756 25956 11762 25968
rect 12345 25959 12403 25965
rect 11756 25928 12020 25956
rect 11756 25916 11762 25928
rect 8478 25888 8484 25900
rect 8439 25860 8484 25888
rect 8478 25848 8484 25860
rect 8536 25848 8542 25900
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10042 25888 10048 25900
rect 9999 25860 10048 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 10652 25860 11529 25888
rect 10652 25848 10658 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11790 25848 11796 25900
rect 11848 25888 11854 25900
rect 11992 25888 12020 25928
rect 12345 25925 12357 25959
rect 12391 25956 12403 25959
rect 14568 25956 14596 25996
rect 14642 25984 14648 26036
rect 14700 26024 14706 26036
rect 14737 26027 14795 26033
rect 14737 26024 14749 26027
rect 14700 25996 14749 26024
rect 14700 25984 14706 25996
rect 14737 25993 14749 25996
rect 14783 25993 14795 26027
rect 14737 25987 14795 25993
rect 15746 25984 15752 26036
rect 15804 26024 15810 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15804 25996 15853 26024
rect 15804 25984 15810 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 15841 25987 15899 25993
rect 31389 26027 31447 26033
rect 31389 25993 31401 26027
rect 31435 26024 31447 26027
rect 31754 26024 31760 26036
rect 31435 25996 31760 26024
rect 31435 25993 31447 25996
rect 31389 25987 31447 25993
rect 31754 25984 31760 25996
rect 31812 25984 31818 26036
rect 14829 25959 14887 25965
rect 14829 25956 14841 25959
rect 12391 25928 14504 25956
rect 14568 25928 14841 25956
rect 12391 25925 12403 25928
rect 12345 25919 12403 25925
rect 12526 25888 12532 25900
rect 11848 25860 11893 25888
rect 11992 25860 12434 25888
rect 12487 25860 12532 25888
rect 11848 25848 11854 25860
rect 8570 25820 8576 25832
rect 8531 25792 8576 25820
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 12406 25684 12434 25860
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25888 12955 25891
rect 12943 25860 13124 25888
rect 12943 25857 12955 25860
rect 12897 25851 12955 25857
rect 12618 25780 12624 25832
rect 12676 25820 12682 25832
rect 12986 25820 12992 25832
rect 12676 25792 12769 25820
rect 12947 25792 12992 25820
rect 12676 25780 12682 25792
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 13096 25820 13124 25860
rect 13170 25848 13176 25900
rect 13228 25888 13234 25900
rect 14476 25897 14504 25928
rect 14829 25925 14841 25928
rect 14875 25925 14887 25959
rect 14829 25919 14887 25925
rect 21177 25959 21235 25965
rect 21177 25925 21189 25959
rect 21223 25956 21235 25959
rect 25590 25956 25596 25968
rect 21223 25928 22586 25956
rect 24964 25928 25596 25956
rect 21223 25925 21235 25928
rect 21177 25919 21235 25925
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 13228 25860 13645 25888
rect 13228 25848 13234 25860
rect 13633 25857 13645 25860
rect 13679 25888 13691 25891
rect 14461 25891 14519 25897
rect 13679 25860 13952 25888
rect 13679 25857 13691 25860
rect 13633 25851 13691 25857
rect 13814 25820 13820 25832
rect 13096 25792 13820 25820
rect 12636 25752 12664 25780
rect 13170 25752 13176 25764
rect 12636 25724 13176 25752
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 13280 25684 13308 25792
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 13924 25820 13952 25860
rect 14461 25857 14473 25891
rect 14507 25857 14519 25891
rect 14918 25888 14924 25900
rect 14879 25860 14924 25888
rect 14461 25851 14519 25857
rect 14918 25848 14924 25860
rect 14976 25848 14982 25900
rect 15654 25848 15660 25900
rect 15712 25888 15718 25900
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 15712 25860 15761 25888
rect 15712 25848 15718 25860
rect 15749 25857 15761 25860
rect 15795 25888 15807 25891
rect 16574 25888 16580 25900
rect 15795 25860 16580 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 21082 25888 21088 25900
rect 20036 25860 21088 25888
rect 20036 25848 20042 25860
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 24673 25891 24731 25897
rect 24673 25857 24685 25891
rect 24719 25857 24731 25891
rect 24854 25888 24860 25900
rect 24815 25860 24860 25888
rect 24673 25851 24731 25857
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 13924 25792 16681 25820
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16850 25820 16856 25832
rect 16811 25792 16856 25820
rect 16669 25783 16727 25789
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25820 18567 25823
rect 18874 25820 18880 25832
rect 18555 25792 18880 25820
rect 18555 25789 18567 25792
rect 18509 25783 18567 25789
rect 18874 25780 18880 25792
rect 18932 25780 18938 25832
rect 19334 25780 19340 25832
rect 19392 25820 19398 25832
rect 21821 25823 21879 25829
rect 21821 25820 21833 25823
rect 19392 25792 21833 25820
rect 19392 25780 19398 25792
rect 21821 25789 21833 25792
rect 21867 25789 21879 25823
rect 21821 25783 21879 25789
rect 22094 25780 22100 25832
rect 22152 25820 22158 25832
rect 22152 25792 22197 25820
rect 22152 25780 22158 25792
rect 22554 25780 22560 25832
rect 22612 25820 22618 25832
rect 23569 25823 23627 25829
rect 23569 25820 23581 25823
rect 22612 25792 23581 25820
rect 22612 25780 22618 25792
rect 23569 25789 23581 25792
rect 23615 25789 23627 25823
rect 23569 25783 23627 25789
rect 13449 25755 13507 25761
rect 13449 25721 13461 25755
rect 13495 25752 13507 25755
rect 14090 25752 14096 25764
rect 13495 25724 14096 25752
rect 13495 25721 13507 25724
rect 13449 25715 13507 25721
rect 14090 25712 14096 25724
rect 14148 25712 14154 25764
rect 24688 25752 24716 25851
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 24964 25897 24992 25928
rect 25590 25916 25596 25928
rect 25648 25916 25654 25968
rect 30558 25956 30564 25968
rect 26068 25928 30564 25956
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25857 25007 25891
rect 24949 25851 25007 25857
rect 25130 25848 25136 25900
rect 25188 25888 25194 25900
rect 25225 25891 25283 25897
rect 25225 25888 25237 25891
rect 25188 25860 25237 25888
rect 25188 25848 25194 25860
rect 25225 25857 25237 25860
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 25038 25780 25044 25832
rect 25096 25820 25102 25832
rect 25240 25820 25268 25851
rect 25406 25848 25412 25900
rect 25464 25888 25470 25900
rect 26068 25897 26096 25928
rect 30558 25916 30564 25928
rect 30616 25956 30622 25968
rect 32490 25956 32496 25968
rect 30616 25928 31156 25956
rect 32451 25928 32496 25956
rect 30616 25916 30622 25928
rect 25869 25891 25927 25897
rect 25869 25888 25881 25891
rect 25464 25860 25881 25888
rect 25464 25848 25470 25860
rect 25869 25857 25881 25860
rect 25915 25857 25927 25891
rect 25869 25851 25927 25857
rect 26053 25891 26111 25897
rect 26053 25857 26065 25891
rect 26099 25857 26111 25891
rect 26970 25888 26976 25900
rect 26931 25860 26976 25888
rect 26053 25851 26111 25857
rect 26970 25848 26976 25860
rect 27028 25848 27034 25900
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25888 28779 25891
rect 28810 25888 28816 25900
rect 28767 25860 28816 25888
rect 28767 25857 28779 25860
rect 28721 25851 28779 25857
rect 28810 25848 28816 25860
rect 28868 25848 28874 25900
rect 29822 25848 29828 25900
rect 29880 25888 29886 25900
rect 30101 25891 30159 25897
rect 30101 25888 30113 25891
rect 29880 25860 30113 25888
rect 29880 25848 29886 25860
rect 30101 25857 30113 25860
rect 30147 25857 30159 25891
rect 30834 25888 30840 25900
rect 30795 25860 30840 25888
rect 30101 25851 30159 25857
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 31128 25897 31156 25928
rect 32490 25916 32496 25928
rect 32548 25916 32554 25968
rect 33226 25916 33232 25968
rect 33284 25916 33290 25968
rect 31113 25891 31171 25897
rect 31113 25857 31125 25891
rect 31159 25857 31171 25891
rect 31113 25851 31171 25857
rect 25096 25792 25141 25820
rect 25240 25792 28948 25820
rect 25096 25780 25102 25792
rect 28920 25761 28948 25792
rect 32122 25780 32128 25832
rect 32180 25820 32186 25832
rect 32217 25823 32275 25829
rect 32217 25820 32229 25823
rect 32180 25792 32229 25820
rect 32180 25780 32186 25792
rect 32217 25789 32229 25792
rect 32263 25789 32275 25823
rect 32217 25783 32275 25789
rect 26237 25755 26295 25761
rect 26237 25752 26249 25755
rect 24688 25724 26249 25752
rect 26237 25721 26249 25724
rect 26283 25721 26295 25755
rect 26237 25715 26295 25721
rect 28905 25755 28963 25761
rect 28905 25721 28917 25755
rect 28951 25721 28963 25755
rect 28905 25715 28963 25721
rect 30285 25755 30343 25761
rect 30285 25721 30297 25755
rect 30331 25752 30343 25755
rect 31478 25752 31484 25764
rect 30331 25724 31484 25752
rect 30331 25721 30343 25724
rect 30285 25715 30343 25721
rect 12406 25656 13308 25684
rect 21082 25644 21088 25696
rect 21140 25684 21146 25696
rect 25222 25684 25228 25696
rect 21140 25656 25228 25684
rect 21140 25644 21146 25656
rect 25222 25644 25228 25656
rect 25280 25644 25286 25696
rect 25409 25687 25467 25693
rect 25409 25653 25421 25687
rect 25455 25684 25467 25687
rect 25590 25684 25596 25696
rect 25455 25656 25596 25684
rect 25455 25653 25467 25656
rect 25409 25647 25467 25653
rect 25590 25644 25596 25656
rect 25648 25644 25654 25696
rect 25958 25684 25964 25696
rect 25919 25656 25964 25684
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 27065 25687 27123 25693
rect 27065 25684 27077 25687
rect 26936 25656 27077 25684
rect 26936 25644 26942 25656
rect 27065 25653 27077 25656
rect 27111 25653 27123 25687
rect 27065 25647 27123 25653
rect 27338 25644 27344 25696
rect 27396 25684 27402 25696
rect 30300 25684 30328 25715
rect 31478 25712 31484 25724
rect 31536 25712 31542 25764
rect 27396 25656 30328 25684
rect 31205 25687 31263 25693
rect 27396 25644 27402 25656
rect 31205 25653 31217 25687
rect 31251 25684 31263 25687
rect 31386 25684 31392 25696
rect 31251 25656 31392 25684
rect 31251 25653 31263 25656
rect 31205 25647 31263 25653
rect 31386 25644 31392 25656
rect 31444 25644 31450 25696
rect 32030 25644 32036 25696
rect 32088 25684 32094 25696
rect 33965 25687 34023 25693
rect 33965 25684 33977 25687
rect 32088 25656 33977 25684
rect 32088 25644 32094 25656
rect 33965 25653 33977 25656
rect 34011 25653 34023 25687
rect 33965 25647 34023 25653
rect 46290 25644 46296 25696
rect 46348 25684 46354 25696
rect 47765 25687 47823 25693
rect 47765 25684 47777 25687
rect 46348 25656 47777 25684
rect 46348 25644 46354 25656
rect 47765 25653 47777 25656
rect 47811 25653 47823 25687
rect 47765 25647 47823 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 11514 25480 11520 25492
rect 11471 25452 11520 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 14366 25480 14372 25492
rect 12492 25452 12537 25480
rect 14327 25452 14372 25480
rect 12492 25440 12498 25452
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 16850 25480 16856 25492
rect 16811 25452 16856 25480
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 22094 25440 22100 25492
rect 22152 25480 22158 25492
rect 22152 25452 22197 25480
rect 22152 25440 22158 25452
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 27801 25483 27859 25489
rect 27801 25480 27813 25483
rect 25280 25452 27813 25480
rect 25280 25440 25286 25452
rect 27801 25449 27813 25452
rect 27847 25449 27859 25483
rect 27801 25443 27859 25449
rect 30653 25483 30711 25489
rect 30653 25449 30665 25483
rect 30699 25449 30711 25483
rect 30834 25480 30840 25492
rect 30795 25452 30840 25480
rect 30653 25443 30711 25449
rect 10594 25372 10600 25424
rect 10652 25412 10658 25424
rect 12526 25412 12532 25424
rect 10652 25384 12532 25412
rect 10652 25372 10658 25384
rect 12526 25372 12532 25384
rect 12584 25412 12590 25424
rect 12986 25412 12992 25424
rect 12584 25384 12992 25412
rect 12584 25372 12590 25384
rect 12986 25372 12992 25384
rect 13044 25372 13050 25424
rect 27062 25412 27068 25424
rect 27023 25384 27068 25412
rect 27062 25372 27068 25384
rect 27120 25372 27126 25424
rect 9493 25347 9551 25353
rect 9493 25313 9505 25347
rect 9539 25344 9551 25347
rect 9674 25344 9680 25356
rect 9539 25316 9680 25344
rect 9539 25313 9551 25316
rect 9493 25307 9551 25313
rect 9674 25304 9680 25316
rect 9732 25304 9738 25356
rect 11698 25344 11704 25356
rect 10796 25316 11704 25344
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 8628 25248 9229 25276
rect 8628 25236 8634 25248
rect 9217 25245 9229 25248
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 9401 25279 9459 25285
rect 9401 25245 9413 25279
rect 9447 25276 9459 25279
rect 9582 25276 9588 25288
rect 9447 25248 9588 25276
rect 9447 25245 9459 25248
rect 9401 25239 9459 25245
rect 1670 25208 1676 25220
rect 1631 25180 1676 25208
rect 1670 25168 1676 25180
rect 1728 25168 1734 25220
rect 9232 25208 9260 25239
rect 9582 25236 9588 25248
rect 9640 25236 9646 25288
rect 9953 25279 10011 25285
rect 9953 25245 9965 25279
rect 9999 25276 10011 25279
rect 10042 25276 10048 25288
rect 9999 25248 10048 25276
rect 9999 25245 10011 25248
rect 9953 25239 10011 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 10594 25276 10600 25288
rect 10555 25248 10600 25276
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10796 25285 10824 25316
rect 11698 25304 11704 25316
rect 11756 25304 11762 25356
rect 12710 25304 12716 25356
rect 12768 25344 12774 25356
rect 14918 25344 14924 25356
rect 12768 25316 14924 25344
rect 12768 25304 12774 25316
rect 14918 25304 14924 25316
rect 14976 25304 14982 25356
rect 16574 25304 16580 25356
rect 16632 25344 16638 25356
rect 16632 25316 19288 25344
rect 16632 25304 16638 25316
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25245 10839 25279
rect 11330 25276 11336 25288
rect 11243 25248 11336 25276
rect 10781 25239 10839 25245
rect 11330 25236 11336 25248
rect 11388 25276 11394 25288
rect 11440 25276 11560 25278
rect 12342 25276 12348 25288
rect 11388 25250 12204 25276
rect 11388 25248 11468 25250
rect 11532 25248 12204 25250
rect 12303 25248 12348 25276
rect 11388 25236 11394 25248
rect 10689 25211 10747 25217
rect 10689 25208 10701 25211
rect 9232 25180 10701 25208
rect 10689 25177 10701 25180
rect 10735 25177 10747 25211
rect 12176 25208 12204 25248
rect 12342 25236 12348 25248
rect 12400 25236 12406 25288
rect 14366 25276 14372 25288
rect 14279 25248 14372 25276
rect 14366 25236 14372 25248
rect 14424 25276 14430 25288
rect 15378 25276 15384 25288
rect 14424 25248 15384 25276
rect 14424 25236 14430 25248
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 16850 25276 16856 25288
rect 16807 25248 16856 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 17696 25285 17724 25316
rect 17681 25279 17739 25285
rect 17681 25245 17693 25279
rect 17727 25245 17739 25279
rect 17681 25239 17739 25245
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18322 25276 18328 25288
rect 18012 25248 18328 25276
rect 18012 25236 18018 25248
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 18506 25276 18512 25288
rect 18467 25248 18512 25276
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 19260 25285 19288 25316
rect 21174 25304 21180 25356
rect 21232 25344 21238 25356
rect 25590 25344 25596 25356
rect 21232 25316 21956 25344
rect 25551 25316 25596 25344
rect 21232 25304 21238 25316
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 21450 25276 21456 25288
rect 21411 25248 21456 25276
rect 19245 25239 19303 25245
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 21542 25236 21548 25288
rect 21600 25276 21606 25288
rect 21600 25248 21645 25276
rect 21600 25236 21606 25248
rect 21726 25236 21732 25288
rect 21784 25276 21790 25288
rect 21928 25285 21956 25316
rect 25590 25304 25596 25316
rect 25648 25304 25654 25356
rect 27816 25344 27844 25443
rect 30006 25372 30012 25424
rect 30064 25412 30070 25424
rect 30668 25412 30696 25443
rect 30834 25440 30840 25452
rect 30892 25440 30898 25492
rect 31386 25480 31392 25492
rect 31347 25452 31392 25480
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 31478 25440 31484 25492
rect 31536 25480 31542 25492
rect 32766 25480 32772 25492
rect 31536 25452 32772 25480
rect 31536 25440 31542 25452
rect 32766 25440 32772 25452
rect 32824 25440 32830 25492
rect 33226 25480 33232 25492
rect 33187 25452 33232 25480
rect 33226 25440 33232 25452
rect 33284 25440 33290 25492
rect 31846 25412 31852 25424
rect 30064 25384 31852 25412
rect 30064 25372 30070 25384
rect 31846 25372 31852 25384
rect 31904 25372 31910 25424
rect 31478 25344 31484 25356
rect 27816 25316 31484 25344
rect 31478 25304 31484 25316
rect 31536 25304 31542 25356
rect 32030 25344 32036 25356
rect 31588 25316 32036 25344
rect 21918 25279 21976 25285
rect 21784 25248 21829 25276
rect 21784 25236 21790 25248
rect 21918 25245 21930 25279
rect 21964 25245 21976 25279
rect 24670 25276 24676 25288
rect 24631 25248 24676 25276
rect 21918 25239 21976 25245
rect 24670 25236 24676 25248
rect 24728 25276 24734 25288
rect 25130 25276 25136 25288
rect 24728 25248 25136 25276
rect 24728 25236 24734 25248
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25314 25276 25320 25288
rect 25275 25248 25320 25276
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 29454 25236 29460 25288
rect 29512 25276 29518 25288
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29512 25248 29561 25276
rect 29512 25236 29518 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 14384 25208 14412 25236
rect 12176 25180 14412 25208
rect 10689 25171 10747 25177
rect 17862 25168 17868 25220
rect 17920 25208 17926 25220
rect 18417 25211 18475 25217
rect 18417 25208 18429 25211
rect 17920 25180 18429 25208
rect 17920 25168 17926 25180
rect 18417 25177 18429 25180
rect 18463 25177 18475 25211
rect 18417 25171 18475 25177
rect 21821 25211 21879 25217
rect 21821 25177 21833 25211
rect 21867 25208 21879 25211
rect 24854 25208 24860 25220
rect 21867 25180 24860 25208
rect 21867 25177 21879 25180
rect 21821 25171 21879 25177
rect 24854 25168 24860 25180
rect 24912 25168 24918 25220
rect 26878 25208 26884 25220
rect 26818 25180 26884 25208
rect 26878 25168 26884 25180
rect 26936 25168 26942 25220
rect 27614 25168 27620 25220
rect 27672 25208 27678 25220
rect 27709 25211 27767 25217
rect 27709 25208 27721 25211
rect 27672 25180 27721 25208
rect 27672 25168 27678 25180
rect 27709 25177 27721 25180
rect 27755 25177 27767 25211
rect 29564 25208 29592 25239
rect 29638 25236 29644 25288
rect 29696 25276 29702 25288
rect 31588 25285 31616 25316
rect 32030 25304 32036 25316
rect 32088 25304 32094 25356
rect 46290 25344 46296 25356
rect 46251 25316 46296 25344
rect 46290 25304 46296 25316
rect 46348 25304 46354 25356
rect 29733 25279 29791 25285
rect 29733 25276 29745 25279
rect 29696 25248 29745 25276
rect 29696 25236 29702 25248
rect 29733 25245 29745 25248
rect 29779 25276 29791 25279
rect 30561 25279 30619 25285
rect 30561 25276 30573 25279
rect 29779 25248 30573 25276
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 30561 25245 30573 25248
rect 30607 25245 30619 25279
rect 30561 25239 30619 25245
rect 30653 25279 30711 25285
rect 30653 25245 30665 25279
rect 30699 25276 30711 25279
rect 31573 25279 31631 25285
rect 31573 25276 31585 25279
rect 30699 25248 31585 25276
rect 30699 25245 30711 25248
rect 30653 25239 30711 25245
rect 31573 25245 31585 25248
rect 31619 25245 31631 25279
rect 31573 25239 31631 25245
rect 31757 25279 31815 25285
rect 31757 25245 31769 25279
rect 31803 25245 31815 25279
rect 31757 25239 31815 25245
rect 30282 25208 30288 25220
rect 29564 25180 30288 25208
rect 27709 25171 27767 25177
rect 30282 25168 30288 25180
rect 30340 25208 30346 25220
rect 30377 25211 30435 25217
rect 30377 25208 30389 25211
rect 30340 25180 30389 25208
rect 30340 25168 30346 25180
rect 30377 25177 30389 25180
rect 30423 25177 30435 25211
rect 30377 25171 30435 25177
rect 9033 25143 9091 25149
rect 9033 25109 9045 25143
rect 9079 25140 9091 25143
rect 9214 25140 9220 25152
rect 9079 25112 9220 25140
rect 9079 25109 9091 25112
rect 9033 25103 9091 25109
rect 9214 25100 9220 25112
rect 9272 25100 9278 25152
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 10045 25143 10103 25149
rect 10045 25140 10057 25143
rect 10008 25112 10057 25140
rect 10008 25100 10014 25112
rect 10045 25109 10057 25112
rect 10091 25109 10103 25143
rect 10045 25103 10103 25109
rect 17773 25143 17831 25149
rect 17773 25109 17785 25143
rect 17819 25140 17831 25143
rect 18046 25140 18052 25152
rect 17819 25112 18052 25140
rect 17819 25109 17831 25112
rect 17773 25103 17831 25109
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 19334 25140 19340 25152
rect 19295 25112 19340 25140
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 24394 25100 24400 25152
rect 24452 25140 24458 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 24452 25112 24777 25140
rect 24452 25100 24458 25112
rect 24765 25109 24777 25112
rect 24811 25109 24823 25143
rect 29914 25140 29920 25152
rect 29875 25112 29920 25140
rect 24765 25103 24823 25109
rect 29914 25100 29920 25112
rect 29972 25140 29978 25152
rect 31772 25140 31800 25239
rect 31846 25236 31852 25288
rect 31904 25276 31910 25288
rect 33134 25276 33140 25288
rect 31904 25248 31949 25276
rect 33095 25248 33140 25276
rect 31904 25236 31910 25248
rect 33134 25236 33140 25248
rect 33192 25236 33198 25288
rect 46477 25211 46535 25217
rect 46477 25177 46489 25211
rect 46523 25208 46535 25211
rect 47670 25208 47676 25220
rect 46523 25180 47676 25208
rect 46523 25177 46535 25180
rect 46477 25171 46535 25177
rect 47670 25168 47676 25180
rect 47728 25168 47734 25220
rect 48130 25208 48136 25220
rect 48091 25180 48136 25208
rect 48130 25168 48136 25180
rect 48188 25168 48194 25220
rect 29972 25112 31800 25140
rect 29972 25100 29978 25112
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 24026 24936 24032 24948
rect 23987 24908 24032 24936
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 25958 24936 25964 24948
rect 24228 24908 25964 24936
rect 8478 24868 8484 24880
rect 7760 24840 8484 24868
rect 7760 24809 7788 24840
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 14366 24868 14372 24880
rect 14327 24840 14372 24868
rect 14366 24828 14372 24840
rect 14424 24828 14430 24880
rect 18046 24828 18052 24880
rect 18104 24828 18110 24880
rect 19334 24828 19340 24880
rect 19392 24868 19398 24880
rect 19392 24840 19734 24868
rect 19392 24828 19398 24840
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24769 7803 24803
rect 10226 24800 10232 24812
rect 10139 24772 10232 24800
rect 7745 24763 7803 24769
rect 10226 24760 10232 24772
rect 10284 24800 10290 24812
rect 11330 24800 11336 24812
rect 10284 24772 11336 24800
rect 10284 24760 10290 24772
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 12621 24803 12679 24809
rect 12621 24800 12633 24803
rect 12584 24772 12633 24800
rect 12584 24760 12590 24772
rect 12621 24769 12633 24772
rect 12667 24769 12679 24803
rect 12802 24800 12808 24812
rect 12763 24772 12808 24800
rect 12621 24763 12679 24769
rect 12802 24760 12808 24772
rect 12860 24760 12866 24812
rect 14001 24803 14059 24809
rect 14001 24769 14013 24803
rect 14047 24800 14059 24803
rect 14090 24800 14096 24812
rect 14047 24772 14096 24800
rect 14047 24769 14059 24772
rect 14001 24763 14059 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 24228 24809 24256 24908
rect 25958 24896 25964 24908
rect 26016 24896 26022 24948
rect 26970 24896 26976 24948
rect 27028 24936 27034 24948
rect 27157 24939 27215 24945
rect 27157 24936 27169 24939
rect 27028 24908 27169 24936
rect 27028 24896 27034 24908
rect 27157 24905 27169 24908
rect 27203 24905 27215 24939
rect 27157 24899 27215 24905
rect 28445 24939 28503 24945
rect 28445 24905 28457 24939
rect 28491 24905 28503 24939
rect 28445 24899 28503 24905
rect 24394 24868 24400 24880
rect 24355 24840 24400 24868
rect 24394 24828 24400 24840
rect 24452 24828 24458 24880
rect 24515 24871 24573 24877
rect 24515 24837 24527 24871
rect 24561 24868 24573 24871
rect 24854 24868 24860 24880
rect 24561 24840 24860 24868
rect 24561 24837 24573 24840
rect 24515 24831 24573 24837
rect 24854 24828 24860 24840
rect 24912 24828 24918 24880
rect 25130 24828 25136 24880
rect 25188 24868 25194 24880
rect 25501 24871 25559 24877
rect 25501 24868 25513 24871
rect 25188 24840 25513 24868
rect 25188 24828 25194 24840
rect 25501 24837 25513 24840
rect 25547 24837 25559 24871
rect 26329 24871 26387 24877
rect 26329 24868 26341 24871
rect 25501 24831 25559 24837
rect 25976 24840 26341 24868
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22066 24772 22661 24800
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8202 24732 8208 24744
rect 7975 24704 8208 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24701 8355 24735
rect 16758 24732 16764 24744
rect 16719 24704 16764 24732
rect 8297 24695 8355 24701
rect 4798 24624 4804 24676
rect 4856 24664 4862 24676
rect 8312 24664 8340 24695
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 17037 24735 17095 24741
rect 17037 24701 17049 24735
rect 17083 24732 17095 24735
rect 17770 24732 17776 24744
rect 17083 24704 17776 24732
rect 17083 24701 17095 24704
rect 17037 24695 17095 24701
rect 17770 24692 17776 24704
rect 17828 24692 17834 24744
rect 18966 24732 18972 24744
rect 18927 24704 18972 24732
rect 18966 24692 18972 24704
rect 19024 24692 19030 24744
rect 19245 24735 19303 24741
rect 19245 24701 19257 24735
rect 19291 24732 19303 24735
rect 20622 24732 20628 24744
rect 19291 24704 20628 24732
rect 19291 24701 19303 24704
rect 19245 24695 19303 24701
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 22066 24664 22094 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 24302 24760 24308 24812
rect 24360 24800 24366 24812
rect 24360 24772 24405 24800
rect 24360 24760 24366 24772
rect 24670 24760 24676 24812
rect 24728 24800 24734 24812
rect 24728 24772 24773 24800
rect 24728 24760 24734 24772
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 25317 24803 25375 24809
rect 25317 24800 25329 24803
rect 25280 24772 25329 24800
rect 25280 24760 25286 24772
rect 25317 24769 25329 24772
rect 25363 24769 25375 24803
rect 25317 24763 25375 24769
rect 25593 24803 25651 24809
rect 25593 24769 25605 24803
rect 25639 24800 25651 24803
rect 25976 24800 26004 24840
rect 26329 24837 26341 24840
rect 26375 24837 26387 24871
rect 27338 24868 27344 24880
rect 26329 24831 26387 24837
rect 26436 24840 27344 24868
rect 25639 24772 26004 24800
rect 26053 24803 26111 24809
rect 25639 24769 25651 24772
rect 25593 24763 25651 24769
rect 26053 24769 26065 24803
rect 26099 24800 26111 24803
rect 26234 24800 26240 24812
rect 26099 24772 26240 24800
rect 26099 24769 26111 24772
rect 26053 24763 26111 24769
rect 26234 24760 26240 24772
rect 26292 24800 26298 24812
rect 26436 24800 26464 24840
rect 27338 24828 27344 24840
rect 27396 24828 27402 24880
rect 26292 24772 26464 24800
rect 26292 24760 26298 24772
rect 26694 24760 26700 24812
rect 26752 24800 26758 24812
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26752 24772 26985 24800
rect 26752 24760 26758 24772
rect 26973 24769 26985 24772
rect 27019 24800 27031 24803
rect 27614 24800 27620 24812
rect 27019 24772 27620 24800
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 27614 24760 27620 24772
rect 27672 24800 27678 24812
rect 28261 24803 28319 24809
rect 28261 24800 28273 24803
rect 27672 24772 28273 24800
rect 27672 24760 27678 24772
rect 28261 24769 28273 24772
rect 28307 24769 28319 24803
rect 28460 24800 28488 24899
rect 29546 24868 29552 24880
rect 29380 24840 29552 24868
rect 29380 24800 29408 24840
rect 29546 24828 29552 24840
rect 29604 24868 29610 24880
rect 29604 24840 30328 24868
rect 29604 24828 29610 24840
rect 29730 24800 29736 24812
rect 28460 24772 29408 24800
rect 29472 24772 29736 24800
rect 28261 24763 28319 24769
rect 25958 24692 25964 24744
rect 26016 24732 26022 24744
rect 26145 24735 26203 24741
rect 26145 24732 26157 24735
rect 26016 24704 26157 24732
rect 26016 24692 26022 24704
rect 26145 24701 26157 24704
rect 26191 24701 26203 24735
rect 26145 24695 26203 24701
rect 26329 24735 26387 24741
rect 26329 24701 26341 24735
rect 26375 24732 26387 24735
rect 28626 24732 28632 24744
rect 26375 24704 28632 24732
rect 26375 24701 26387 24704
rect 26329 24695 26387 24701
rect 28626 24692 28632 24704
rect 28684 24732 28690 24744
rect 29472 24732 29500 24772
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 29825 24803 29883 24809
rect 29825 24769 29837 24803
rect 29871 24800 29883 24803
rect 30006 24800 30012 24812
rect 29871 24772 30012 24800
rect 29871 24769 29883 24772
rect 29825 24763 29883 24769
rect 30006 24760 30012 24772
rect 30064 24760 30070 24812
rect 30098 24760 30104 24812
rect 30156 24800 30162 24812
rect 30300 24800 30328 24840
rect 30760 24840 30972 24868
rect 30760 24800 30788 24840
rect 30156 24772 30201 24800
rect 30300 24772 30788 24800
rect 30837 24803 30895 24809
rect 30156 24760 30162 24772
rect 30837 24769 30849 24803
rect 30883 24769 30895 24803
rect 30944 24800 30972 24840
rect 32217 24803 32275 24809
rect 32217 24800 32229 24803
rect 30944 24772 32229 24800
rect 30837 24763 30895 24769
rect 32217 24769 32229 24772
rect 32263 24800 32275 24803
rect 33134 24800 33140 24812
rect 32263 24772 33140 24800
rect 32263 24769 32275 24772
rect 32217 24763 32275 24769
rect 28684 24704 29500 24732
rect 29549 24735 29607 24741
rect 28684 24692 28690 24704
rect 29549 24701 29561 24735
rect 29595 24732 29607 24735
rect 30852 24732 30880 24763
rect 33134 24760 33140 24772
rect 33192 24760 33198 24812
rect 46750 24800 46756 24812
rect 35866 24772 46756 24800
rect 31110 24732 31116 24744
rect 29595 24724 29684 24732
rect 29840 24724 30880 24732
rect 29595 24704 30880 24724
rect 31071 24704 31116 24732
rect 29595 24701 29607 24704
rect 29549 24695 29607 24701
rect 29656 24696 29868 24704
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 4856 24636 8340 24664
rect 18064 24636 18644 24664
rect 4856 24624 4862 24636
rect 3694 24556 3700 24608
rect 3752 24596 3758 24608
rect 8570 24596 8576 24608
rect 3752 24568 8576 24596
rect 3752 24556 3758 24568
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 10045 24599 10103 24605
rect 10045 24596 10057 24599
rect 8996 24568 10057 24596
rect 8996 24556 9002 24568
rect 10045 24565 10057 24568
rect 10091 24565 10103 24599
rect 10045 24559 10103 24565
rect 12618 24556 12624 24608
rect 12676 24596 12682 24608
rect 12713 24599 12771 24605
rect 12713 24596 12725 24599
rect 12676 24568 12725 24596
rect 12676 24556 12682 24568
rect 12713 24565 12725 24568
rect 12759 24565 12771 24599
rect 12713 24559 12771 24565
rect 15194 24556 15200 24608
rect 15252 24596 15258 24608
rect 15838 24596 15844 24608
rect 15252 24568 15844 24596
rect 15252 24556 15258 24568
rect 15838 24556 15844 24568
rect 15896 24596 15902 24608
rect 18064 24596 18092 24636
rect 15896 24568 18092 24596
rect 15896 24556 15902 24568
rect 18138 24556 18144 24608
rect 18196 24596 18202 24608
rect 18506 24596 18512 24608
rect 18196 24568 18512 24596
rect 18196 24556 18202 24568
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 18616 24596 18644 24636
rect 20272 24636 22094 24664
rect 20272 24596 20300 24636
rect 24762 24624 24768 24676
rect 24820 24664 24826 24676
rect 35866 24664 35894 24772
rect 46750 24760 46756 24772
rect 46808 24760 46814 24812
rect 46845 24803 46903 24809
rect 46845 24769 46857 24803
rect 46891 24769 46903 24803
rect 46845 24763 46903 24769
rect 45922 24692 45928 24744
rect 45980 24732 45986 24744
rect 46106 24732 46112 24744
rect 45980 24704 46112 24732
rect 45980 24692 45986 24704
rect 46106 24692 46112 24704
rect 46164 24732 46170 24744
rect 46860 24732 46888 24763
rect 47486 24760 47492 24812
rect 47544 24800 47550 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47544 24772 47593 24800
rect 47544 24760 47550 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 47670 24760 47676 24812
rect 47728 24800 47734 24812
rect 47728 24772 47773 24800
rect 47728 24760 47734 24772
rect 46164 24704 46888 24732
rect 46164 24692 46170 24704
rect 24820 24636 35894 24664
rect 24820 24624 24826 24636
rect 18616 24568 20300 24596
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20717 24599 20775 24605
rect 20717 24596 20729 24599
rect 20588 24568 20729 24596
rect 20588 24556 20594 24568
rect 20717 24565 20729 24568
rect 20763 24565 20775 24599
rect 22830 24596 22836 24608
rect 22791 24568 22836 24596
rect 20717 24559 20775 24565
rect 22830 24556 22836 24568
rect 22888 24556 22894 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 25133 24599 25191 24605
rect 25133 24596 25145 24599
rect 24728 24568 25145 24596
rect 24728 24556 24734 24568
rect 25133 24565 25145 24568
rect 25179 24565 25191 24599
rect 25133 24559 25191 24565
rect 25222 24556 25228 24608
rect 25280 24596 25286 24608
rect 28258 24596 28264 24608
rect 25280 24568 28264 24596
rect 25280 24556 25286 24568
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 30006 24596 30012 24608
rect 29967 24568 30012 24596
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 30650 24596 30656 24608
rect 30611 24568 30656 24596
rect 30650 24556 30656 24568
rect 30708 24556 30714 24608
rect 31018 24596 31024 24608
rect 30979 24568 31024 24596
rect 31018 24556 31024 24568
rect 31076 24556 31082 24608
rect 32309 24599 32367 24605
rect 32309 24565 32321 24599
rect 32355 24596 32367 24599
rect 32398 24596 32404 24608
rect 32355 24568 32404 24596
rect 32355 24565 32367 24568
rect 32309 24559 32367 24565
rect 32398 24556 32404 24568
rect 32456 24556 32462 24608
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 46937 24599 46995 24605
rect 46937 24596 46949 24599
rect 46532 24568 46949 24596
rect 46532 24556 46538 24568
rect 46937 24565 46949 24568
rect 46983 24565 46995 24599
rect 46937 24559 46995 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 8202 24392 8208 24404
rect 8163 24364 8208 24392
rect 8202 24352 8208 24364
rect 8260 24352 8266 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 10689 24395 10747 24401
rect 10689 24392 10701 24395
rect 9732 24364 10701 24392
rect 9732 24352 9738 24364
rect 10689 24361 10701 24364
rect 10735 24392 10747 24395
rect 11698 24392 11704 24404
rect 10735 24364 11192 24392
rect 11659 24364 11704 24392
rect 10735 24361 10747 24364
rect 10689 24355 10747 24361
rect 11164 24333 11192 24364
rect 11698 24352 11704 24364
rect 11756 24352 11762 24404
rect 18966 24352 18972 24404
rect 19024 24392 19030 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 19024 24364 19257 24392
rect 19024 24352 19030 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 20622 24392 20628 24404
rect 20583 24364 20628 24392
rect 19245 24355 19303 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 25038 24392 25044 24404
rect 22066 24364 25044 24392
rect 11149 24327 11207 24333
rect 11149 24293 11161 24327
rect 11195 24293 11207 24327
rect 11149 24287 11207 24293
rect 14734 24284 14740 24336
rect 14792 24324 14798 24336
rect 22066 24324 22094 24364
rect 25038 24352 25044 24364
rect 25096 24352 25102 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 26145 24395 26203 24401
rect 26145 24392 26157 24395
rect 25188 24364 26157 24392
rect 25188 24352 25194 24364
rect 26145 24361 26157 24364
rect 26191 24361 26203 24395
rect 26145 24355 26203 24361
rect 28721 24395 28779 24401
rect 28721 24361 28733 24395
rect 28767 24392 28779 24395
rect 29454 24392 29460 24404
rect 28767 24364 29460 24392
rect 28767 24361 28779 24364
rect 28721 24355 28779 24361
rect 29454 24352 29460 24364
rect 29512 24352 29518 24404
rect 30190 24352 30196 24404
rect 30248 24352 30254 24404
rect 30561 24395 30619 24401
rect 30561 24361 30573 24395
rect 30607 24392 30619 24395
rect 31018 24392 31024 24404
rect 30607 24364 31024 24392
rect 30607 24361 30619 24364
rect 30561 24355 30619 24361
rect 31018 24352 31024 24364
rect 31076 24352 31082 24404
rect 31846 24352 31852 24404
rect 31904 24392 31910 24404
rect 32861 24395 32919 24401
rect 32861 24392 32873 24395
rect 31904 24364 32873 24392
rect 31904 24352 31910 24364
rect 32861 24361 32873 24364
rect 32907 24361 32919 24395
rect 40034 24392 40040 24404
rect 32861 24355 32919 24361
rect 35866 24364 40040 24392
rect 14792 24296 22094 24324
rect 14792 24284 14798 24296
rect 28810 24284 28816 24336
rect 28868 24324 28874 24336
rect 30208 24324 30236 24352
rect 30926 24324 30932 24336
rect 28868 24296 30932 24324
rect 28868 24284 28874 24296
rect 30926 24284 30932 24296
rect 30984 24284 30990 24336
rect 8938 24256 8944 24268
rect 8899 24228 8944 24256
rect 8938 24216 8944 24228
rect 8996 24216 9002 24268
rect 9214 24256 9220 24268
rect 9175 24228 9220 24256
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 12066 24256 12072 24268
rect 9640 24228 12072 24256
rect 9640 24216 9646 24228
rect 12066 24216 12072 24228
rect 12124 24216 12130 24268
rect 12618 24256 12624 24268
rect 12579 24228 12624 24256
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 14277 24259 14335 24265
rect 14277 24225 14289 24259
rect 14323 24256 14335 24259
rect 15194 24256 15200 24268
rect 14323 24228 15200 24256
rect 14323 24225 14335 24228
rect 14277 24219 14335 24225
rect 15194 24216 15200 24228
rect 15252 24216 15258 24268
rect 17402 24256 17408 24268
rect 17363 24228 17408 24256
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 17586 24216 17592 24268
rect 17644 24256 17650 24268
rect 20073 24259 20131 24265
rect 17644 24228 19380 24256
rect 17644 24216 17650 24228
rect 19352 24200 19380 24228
rect 20073 24225 20085 24259
rect 20119 24256 20131 24259
rect 24397 24259 24455 24265
rect 20119 24228 20668 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 11425 24191 11483 24197
rect 11425 24188 11437 24191
rect 10836 24160 11437 24188
rect 10836 24148 10842 24160
rect 11425 24157 11437 24160
rect 11471 24188 11483 24191
rect 11698 24188 11704 24200
rect 11471 24160 11704 24188
rect 11471 24157 11483 24160
rect 11425 24151 11483 24157
rect 11698 24148 11704 24160
rect 11756 24188 11762 24200
rect 12713 24191 12771 24197
rect 12713 24188 12725 24191
rect 11756 24160 12725 24188
rect 11756 24148 11762 24160
rect 12713 24157 12725 24160
rect 12759 24157 12771 24191
rect 12713 24151 12771 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 14826 24188 14832 24200
rect 14599 24160 14832 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 9950 24080 9956 24132
rect 10008 24080 10014 24132
rect 12728 24120 12756 24151
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 15565 24191 15623 24197
rect 15565 24188 15577 24191
rect 14976 24160 15577 24188
rect 14976 24148 14982 24160
rect 15565 24157 15577 24160
rect 15611 24157 15623 24191
rect 18138 24188 18144 24200
rect 18099 24160 18144 24188
rect 15565 24151 15623 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18322 24188 18328 24200
rect 18283 24160 18328 24188
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 19334 24188 19340 24200
rect 19295 24160 19340 24188
rect 19334 24148 19340 24160
rect 19392 24148 19398 24200
rect 19981 24191 20039 24197
rect 19981 24190 19993 24191
rect 19904 24162 19993 24190
rect 14936 24120 14964 24148
rect 15746 24120 15752 24132
rect 12728 24092 14964 24120
rect 15707 24092 15752 24120
rect 15746 24080 15752 24092
rect 15804 24080 15810 24132
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 18509 24123 18567 24129
rect 18509 24120 18521 24123
rect 18012 24092 18521 24120
rect 18012 24080 18018 24092
rect 18509 24089 18521 24092
rect 18555 24120 18567 24123
rect 19904 24120 19932 24162
rect 19981 24157 19993 24162
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24188 20223 24191
rect 20530 24188 20536 24200
rect 20211 24160 20536 24188
rect 20211 24157 20223 24160
rect 20165 24151 20223 24157
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 20640 24197 20668 24228
rect 24397 24225 24409 24259
rect 24443 24256 24455 24259
rect 25314 24256 25320 24268
rect 24443 24228 25320 24256
rect 24443 24225 24455 24228
rect 24397 24219 24455 24225
rect 25314 24216 25320 24228
rect 25372 24256 25378 24268
rect 27246 24256 27252 24268
rect 25372 24228 27016 24256
rect 27207 24228 27252 24256
rect 25372 24216 25378 24228
rect 26988 24200 27016 24228
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 29914 24216 29920 24268
rect 29972 24256 29978 24268
rect 30193 24259 30251 24265
rect 30193 24256 30205 24259
rect 29972 24228 30205 24256
rect 29972 24216 29978 24228
rect 30193 24225 30205 24228
rect 30239 24225 30251 24259
rect 31110 24256 31116 24268
rect 31023 24228 31116 24256
rect 30193 24219 30251 24225
rect 31110 24216 31116 24228
rect 31168 24256 31174 24268
rect 32122 24256 32128 24268
rect 31168 24228 32128 24256
rect 31168 24216 31174 24228
rect 32122 24216 32128 24228
rect 32180 24216 32186 24268
rect 20625 24191 20683 24197
rect 20625 24157 20637 24191
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 26970 24188 26976 24200
rect 26931 24160 26976 24188
rect 20809 24151 20867 24157
rect 18555 24092 19932 24120
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 11238 24012 11244 24064
rect 11296 24052 11302 24064
rect 11333 24055 11391 24061
rect 11333 24052 11345 24055
rect 11296 24024 11345 24052
rect 11296 24012 11302 24024
rect 11333 24021 11345 24024
rect 11379 24021 11391 24055
rect 11333 24015 11391 24021
rect 11517 24055 11575 24061
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 11790 24052 11796 24064
rect 11563 24024 11796 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 13446 24052 13452 24064
rect 13127 24024 13452 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 19058 24012 19064 24064
rect 19116 24052 19122 24064
rect 20824 24052 20852 24151
rect 26970 24148 26976 24160
rect 27028 24148 27034 24200
rect 30098 24148 30104 24200
rect 30156 24188 30162 24200
rect 30285 24191 30343 24197
rect 30285 24188 30297 24191
rect 30156 24160 30297 24188
rect 30156 24148 30162 24160
rect 30285 24157 30297 24160
rect 30331 24157 30343 24191
rect 35866 24188 35894 24364
rect 40034 24352 40040 24364
rect 40092 24352 40098 24404
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 46290 24188 46296 24200
rect 30285 24151 30343 24157
rect 32692 24160 35894 24188
rect 46251 24160 46296 24188
rect 24670 24120 24676 24132
rect 24631 24092 24676 24120
rect 24670 24080 24676 24092
rect 24728 24080 24734 24132
rect 26326 24120 26332 24132
rect 25898 24092 26332 24120
rect 26326 24080 26332 24092
rect 26384 24080 26390 24132
rect 27982 24080 27988 24132
rect 28040 24080 28046 24132
rect 28644 24092 28856 24120
rect 19116 24024 20852 24052
rect 19116 24012 19122 24024
rect 22830 24012 22836 24064
rect 22888 24052 22894 24064
rect 26694 24052 26700 24064
rect 22888 24024 26700 24052
rect 22888 24012 22894 24024
rect 26694 24012 26700 24024
rect 26752 24052 26758 24064
rect 27338 24052 27344 24064
rect 26752 24024 27344 24052
rect 26752 24012 26758 24024
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 27890 24012 27896 24064
rect 27948 24052 27954 24064
rect 28644 24052 28672 24092
rect 27948 24024 28672 24052
rect 28828 24052 28856 24092
rect 30650 24080 30656 24132
rect 30708 24120 30714 24132
rect 31389 24123 31447 24129
rect 31389 24120 31401 24123
rect 30708 24092 31401 24120
rect 30708 24080 30714 24092
rect 31389 24089 31401 24092
rect 31435 24089 31447 24123
rect 31389 24083 31447 24089
rect 32398 24080 32404 24132
rect 32456 24080 32462 24132
rect 32692 24052 32720 24160
rect 46290 24148 46296 24160
rect 46348 24148 46354 24200
rect 28828 24024 32720 24052
rect 27948 24012 27954 24024
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1949 23851 2007 23857
rect 1949 23817 1961 23851
rect 1995 23848 2007 23851
rect 14734 23848 14740 23860
rect 1995 23820 14740 23848
rect 1995 23817 2007 23820
rect 1949 23811 2007 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 14918 23848 14924 23860
rect 14879 23820 14924 23848
rect 14918 23808 14924 23820
rect 14976 23808 14982 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15749 23851 15807 23857
rect 15749 23848 15761 23851
rect 15712 23820 15761 23848
rect 15712 23808 15718 23820
rect 15749 23817 15761 23820
rect 15795 23817 15807 23851
rect 15749 23811 15807 23817
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17037 23851 17095 23857
rect 17037 23848 17049 23851
rect 16816 23820 17049 23848
rect 16816 23808 16822 23820
rect 17037 23817 17049 23820
rect 17083 23817 17095 23851
rect 17037 23811 17095 23817
rect 17770 23808 17776 23860
rect 17828 23848 17834 23860
rect 17865 23851 17923 23857
rect 17865 23848 17877 23851
rect 17828 23820 17877 23848
rect 17828 23808 17834 23820
rect 17865 23817 17877 23820
rect 17911 23817 17923 23851
rect 17865 23811 17923 23817
rect 18322 23808 18328 23860
rect 18380 23848 18386 23860
rect 18893 23851 18951 23857
rect 18893 23848 18905 23851
rect 18380 23820 18905 23848
rect 18380 23808 18386 23820
rect 18892 23817 18905 23820
rect 18939 23817 18951 23851
rect 19058 23848 19064 23860
rect 19019 23820 19064 23848
rect 18892 23811 18951 23817
rect 10612 23752 11652 23780
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23712 9551 23715
rect 9582 23712 9588 23724
rect 9539 23684 9588 23712
rect 9539 23681 9551 23684
rect 9493 23675 9551 23681
rect 9324 23576 9352 23675
rect 9582 23672 9588 23684
rect 9640 23672 9646 23724
rect 9950 23712 9956 23724
rect 9911 23684 9956 23712
rect 9950 23672 9956 23684
rect 10008 23672 10014 23724
rect 10612 23721 10640 23752
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23681 10655 23715
rect 10597 23675 10655 23681
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23712 10747 23715
rect 10965 23715 11023 23721
rect 10735 23684 10916 23712
rect 10735 23681 10747 23684
rect 10689 23675 10747 23681
rect 10778 23644 10784 23656
rect 10739 23616 10784 23644
rect 10778 23604 10784 23616
rect 10836 23604 10842 23656
rect 10888 23644 10916 23684
rect 10965 23681 10977 23715
rect 11011 23712 11023 23715
rect 11011 23684 11284 23712
rect 11011 23681 11023 23684
rect 10965 23675 11023 23681
rect 10888 23616 11100 23644
rect 10965 23579 11023 23585
rect 10965 23576 10977 23579
rect 9324 23548 10977 23576
rect 10965 23545 10977 23548
rect 11011 23545 11023 23579
rect 10965 23539 11023 23545
rect 9309 23511 9367 23517
rect 9309 23477 9321 23511
rect 9355 23508 9367 23511
rect 9766 23508 9772 23520
rect 9355 23480 9772 23508
rect 9355 23477 9367 23480
rect 9309 23471 9367 23477
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 10042 23508 10048 23520
rect 10003 23480 10048 23508
rect 10042 23468 10048 23480
rect 10100 23468 10106 23520
rect 11072 23508 11100 23616
rect 11256 23588 11284 23684
rect 11238 23536 11244 23588
rect 11296 23576 11302 23588
rect 11517 23579 11575 23585
rect 11517 23576 11529 23579
rect 11296 23548 11529 23576
rect 11296 23536 11302 23548
rect 11517 23545 11529 23548
rect 11563 23545 11575 23579
rect 11624 23576 11652 23752
rect 11698 23740 11704 23792
rect 11756 23780 11762 23792
rect 12526 23780 12532 23792
rect 11756 23752 11801 23780
rect 12268 23752 12532 23780
rect 11756 23740 11762 23752
rect 11790 23712 11796 23724
rect 11703 23684 11796 23712
rect 11790 23672 11796 23684
rect 11848 23672 11854 23724
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23712 11943 23715
rect 12268 23712 12296 23752
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 13446 23780 13452 23792
rect 13407 23752 13452 23780
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 13998 23740 14004 23792
rect 14056 23740 14062 23792
rect 18693 23783 18751 23789
rect 18693 23749 18705 23783
rect 18739 23749 18751 23783
rect 18892 23780 18920 23811
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 20806 23848 20812 23860
rect 19392 23820 20812 23848
rect 19392 23808 19398 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 26326 23848 26332 23860
rect 26287 23820 26332 23848
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 26970 23808 26976 23860
rect 27028 23848 27034 23860
rect 31110 23848 31116 23860
rect 27028 23820 31116 23848
rect 27028 23808 27034 23820
rect 24121 23783 24179 23789
rect 18892 23752 19748 23780
rect 18693 23743 18751 23749
rect 11931 23684 12296 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 15565 23715 15623 23721
rect 15565 23712 15577 23715
rect 14884 23684 15577 23712
rect 14884 23672 14890 23684
rect 15565 23681 15577 23684
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 16942 23672 16948 23724
rect 17000 23712 17006 23724
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 17000 23684 17049 23712
rect 17000 23672 17006 23684
rect 17037 23681 17049 23684
rect 17083 23712 17095 23715
rect 17586 23712 17592 23724
rect 17083 23684 17592 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17586 23672 17592 23684
rect 17644 23672 17650 23724
rect 17773 23715 17831 23721
rect 17773 23681 17785 23715
rect 17819 23712 17831 23715
rect 17862 23712 17868 23724
rect 17819 23684 17868 23712
rect 17819 23681 17831 23684
rect 17773 23675 17831 23681
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 18708 23712 18736 23743
rect 19334 23712 19340 23724
rect 18012 23684 18057 23712
rect 18708 23684 19340 23712
rect 18012 23672 18018 23684
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 19610 23712 19616 23724
rect 19571 23684 19616 23712
rect 19610 23672 19616 23684
rect 19668 23672 19674 23724
rect 19720 23721 19748 23752
rect 24121 23749 24133 23783
rect 24167 23780 24179 23783
rect 27890 23780 27896 23792
rect 24167 23752 27896 23780
rect 24167 23749 24179 23752
rect 24121 23743 24179 23749
rect 27890 23740 27896 23752
rect 27948 23740 27954 23792
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23681 20499 23715
rect 20441 23675 20499 23681
rect 11808 23644 11836 23672
rect 12618 23644 12624 23656
rect 11808 23616 12624 23644
rect 12618 23604 12624 23616
rect 12676 23644 12682 23656
rect 12802 23644 12808 23656
rect 12676 23616 12808 23644
rect 12676 23604 12682 23616
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 13170 23644 13176 23656
rect 13131 23616 13176 23644
rect 13170 23604 13176 23616
rect 13228 23604 13234 23656
rect 14090 23604 14096 23656
rect 14148 23644 14154 23656
rect 20456 23644 20484 23675
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 22281 23715 22339 23721
rect 22281 23712 22293 23715
rect 20588 23684 22293 23712
rect 20588 23672 20594 23684
rect 22281 23681 22293 23684
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 25038 23712 25044 23724
rect 24719 23684 25044 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25590 23712 25596 23724
rect 25503 23684 25596 23712
rect 25590 23672 25596 23684
rect 25648 23712 25654 23724
rect 26237 23715 26295 23721
rect 25648 23684 26188 23712
rect 25648 23672 25654 23684
rect 22462 23644 22468 23656
rect 14148 23616 20484 23644
rect 22423 23616 22468 23644
rect 14148 23604 14154 23616
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 11624 23548 12434 23576
rect 11517 23539 11575 23545
rect 11790 23508 11796 23520
rect 11072 23480 11796 23508
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12066 23508 12072 23520
rect 12027 23480 12072 23508
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 12406 23508 12434 23548
rect 16850 23536 16856 23588
rect 16908 23576 16914 23588
rect 24857 23579 24915 23585
rect 24857 23576 24869 23579
rect 16908 23548 24869 23576
rect 16908 23536 16914 23548
rect 24857 23545 24869 23548
rect 24903 23545 24915 23579
rect 24857 23539 24915 23545
rect 12710 23508 12716 23520
rect 12406 23480 12716 23508
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18877 23511 18935 23517
rect 18877 23508 18889 23511
rect 18196 23480 18889 23508
rect 18196 23468 18202 23480
rect 18877 23477 18889 23480
rect 18923 23477 18935 23511
rect 18877 23471 18935 23477
rect 19889 23511 19947 23517
rect 19889 23477 19901 23511
rect 19935 23508 19947 23511
rect 20346 23508 20352 23520
rect 19935 23480 20352 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 20625 23511 20683 23517
rect 20625 23477 20637 23511
rect 20671 23508 20683 23511
rect 20806 23508 20812 23520
rect 20671 23480 20812 23508
rect 20671 23477 20683 23480
rect 20625 23471 20683 23477
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25685 23511 25743 23517
rect 25685 23508 25697 23511
rect 25096 23480 25697 23508
rect 25096 23468 25102 23480
rect 25685 23477 25697 23480
rect 25731 23477 25743 23511
rect 26160 23508 26188 23684
rect 26237 23681 26249 23715
rect 26283 23712 26295 23715
rect 26878 23712 26884 23724
rect 26283 23684 26884 23712
rect 26283 23681 26295 23684
rect 26237 23675 26295 23681
rect 26878 23672 26884 23684
rect 26936 23672 26942 23724
rect 28184 23721 28212 23820
rect 31110 23808 31116 23820
rect 31168 23808 31174 23860
rect 47762 23848 47768 23860
rect 38626 23820 47768 23848
rect 28994 23740 29000 23792
rect 29052 23740 29058 23792
rect 29914 23740 29920 23792
rect 29972 23780 29978 23792
rect 29972 23752 31616 23780
rect 29972 23740 29978 23752
rect 28169 23715 28227 23721
rect 28169 23681 28181 23715
rect 28215 23681 28227 23715
rect 28169 23675 28227 23681
rect 29730 23672 29736 23724
rect 29788 23712 29794 23724
rect 30561 23715 30619 23721
rect 30561 23712 30573 23715
rect 29788 23684 30573 23712
rect 29788 23672 29794 23684
rect 30561 23681 30573 23684
rect 30607 23681 30619 23715
rect 30561 23675 30619 23681
rect 30650 23672 30656 23724
rect 30708 23712 30714 23724
rect 30926 23712 30932 23724
rect 30708 23684 30801 23712
rect 30887 23684 30932 23712
rect 30708 23672 30714 23684
rect 28445 23647 28503 23653
rect 28445 23613 28457 23647
rect 28491 23644 28503 23647
rect 29454 23644 29460 23656
rect 28491 23616 29460 23644
rect 28491 23613 28503 23616
rect 28445 23607 28503 23613
rect 29454 23604 29460 23616
rect 29512 23604 29518 23656
rect 29638 23604 29644 23656
rect 29696 23644 29702 23656
rect 29917 23647 29975 23653
rect 29917 23644 29929 23647
rect 29696 23616 29929 23644
rect 29696 23604 29702 23616
rect 29917 23613 29929 23616
rect 29963 23644 29975 23647
rect 30760 23644 30788 23684
rect 30926 23672 30932 23684
rect 30984 23672 30990 23724
rect 31386 23712 31392 23724
rect 31347 23684 31392 23712
rect 31386 23672 31392 23684
rect 31444 23672 31450 23724
rect 31588 23721 31616 23752
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23681 31631 23715
rect 31573 23675 31631 23681
rect 38626 23644 38654 23820
rect 47762 23808 47768 23820
rect 47820 23808 47826 23860
rect 46290 23672 46296 23724
rect 46348 23712 46354 23724
rect 47765 23715 47823 23721
rect 47765 23712 47777 23715
rect 46348 23684 47777 23712
rect 46348 23672 46354 23684
rect 47765 23681 47777 23684
rect 47811 23681 47823 23715
rect 47765 23675 47823 23681
rect 46198 23644 46204 23656
rect 29963 23616 30788 23644
rect 30852 23616 38654 23644
rect 46159 23616 46204 23644
rect 29963 23613 29975 23616
rect 29917 23607 29975 23613
rect 30852 23576 30880 23616
rect 46198 23604 46204 23616
rect 46256 23604 46262 23656
rect 46477 23647 46535 23653
rect 46477 23613 46489 23647
rect 46523 23613 46535 23647
rect 46477 23607 46535 23613
rect 45278 23576 45284 23588
rect 29932 23548 30880 23576
rect 30944 23548 45284 23576
rect 29932 23508 29960 23548
rect 26160 23480 29960 23508
rect 25685 23471 25743 23477
rect 30006 23468 30012 23520
rect 30064 23508 30070 23520
rect 30190 23508 30196 23520
rect 30064 23480 30196 23508
rect 30064 23468 30070 23480
rect 30190 23468 30196 23480
rect 30248 23468 30254 23520
rect 30374 23508 30380 23520
rect 30335 23480 30380 23508
rect 30374 23468 30380 23480
rect 30432 23468 30438 23520
rect 30837 23511 30895 23517
rect 30837 23477 30849 23511
rect 30883 23508 30895 23511
rect 30944 23508 30972 23548
rect 45278 23536 45284 23548
rect 45336 23536 45342 23588
rect 45462 23536 45468 23588
rect 45520 23576 45526 23588
rect 46492 23576 46520 23607
rect 45520 23548 46520 23576
rect 45520 23536 45526 23548
rect 31478 23508 31484 23520
rect 30883 23480 30972 23508
rect 31439 23480 31484 23508
rect 30883 23477 30895 23480
rect 30837 23471 30895 23477
rect 31478 23468 31484 23480
rect 31536 23468 31542 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 9950 23264 9956 23316
rect 10008 23304 10014 23316
rect 12342 23304 12348 23316
rect 10008 23276 12348 23304
rect 10008 23264 10014 23276
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 13081 23307 13139 23313
rect 13081 23273 13093 23307
rect 13127 23304 13139 23307
rect 13170 23304 13176 23316
rect 13127 23276 13176 23304
rect 13127 23273 13139 23276
rect 13081 23267 13139 23273
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 15746 23304 15752 23316
rect 15707 23276 15752 23304
rect 15746 23264 15752 23276
rect 15804 23264 15810 23316
rect 19610 23264 19616 23316
rect 19668 23304 19674 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 19668 23276 19809 23304
rect 19668 23264 19674 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 19797 23267 19855 23273
rect 22462 23264 22468 23316
rect 22520 23304 22526 23316
rect 23017 23307 23075 23313
rect 23017 23304 23029 23307
rect 22520 23276 23029 23304
rect 22520 23264 22526 23276
rect 23017 23273 23029 23276
rect 23063 23273 23075 23307
rect 27982 23304 27988 23316
rect 27943 23276 27988 23304
rect 23017 23267 23075 23273
rect 27982 23264 27988 23276
rect 28040 23264 28046 23316
rect 28629 23307 28687 23313
rect 28629 23273 28641 23307
rect 28675 23304 28687 23307
rect 28994 23304 29000 23316
rect 28675 23276 29000 23304
rect 28675 23273 28687 23276
rect 28629 23267 28687 23273
rect 28994 23264 29000 23276
rect 29052 23264 29058 23316
rect 29454 23264 29460 23316
rect 29512 23304 29518 23316
rect 29549 23307 29607 23313
rect 29549 23304 29561 23307
rect 29512 23276 29561 23304
rect 29512 23264 29518 23276
rect 29549 23273 29561 23276
rect 29595 23273 29607 23307
rect 29549 23267 29607 23273
rect 30561 23307 30619 23313
rect 30561 23273 30573 23307
rect 30607 23304 30619 23307
rect 31386 23304 31392 23316
rect 30607 23276 31392 23304
rect 30607 23273 30619 23276
rect 30561 23267 30619 23273
rect 31386 23264 31392 23276
rect 31444 23264 31450 23316
rect 15654 23196 15660 23248
rect 15712 23196 15718 23248
rect 29917 23239 29975 23245
rect 29917 23205 29929 23239
rect 29963 23236 29975 23239
rect 31478 23236 31484 23248
rect 29963 23208 31484 23236
rect 29963 23205 29975 23208
rect 29917 23199 29975 23205
rect 31478 23196 31484 23208
rect 31536 23196 31542 23248
rect 9766 23168 9772 23180
rect 9727 23140 9772 23168
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 15672 23168 15700 23196
rect 19245 23171 19303 23177
rect 15672 23140 17632 23168
rect 9490 23100 9496 23112
rect 9451 23072 9496 23100
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13078 23100 13084 23112
rect 13035 23072 13084 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23100 14151 23103
rect 14826 23100 14832 23112
rect 14139 23072 14832 23100
rect 14139 23069 14151 23072
rect 14093 23063 14151 23069
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15654 23100 15660 23112
rect 15615 23072 15660 23100
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 16942 23100 16948 23112
rect 16903 23072 16948 23100
rect 16942 23060 16948 23072
rect 17000 23060 17006 23112
rect 17604 23109 17632 23140
rect 19245 23137 19257 23171
rect 19291 23168 19303 23171
rect 19978 23168 19984 23180
rect 19291 23140 19984 23168
rect 19291 23137 19303 23140
rect 19245 23131 19303 23137
rect 19978 23128 19984 23140
rect 20036 23168 20042 23180
rect 20036 23140 22508 23168
rect 20036 23128 20042 23140
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 19392 23072 19533 23100
rect 19392 23060 19398 23072
rect 19521 23069 19533 23072
rect 19567 23100 19579 23103
rect 20530 23100 20536 23112
rect 19567 23072 20536 23100
rect 19567 23069 19579 23072
rect 19521 23063 19579 23069
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20714 23100 20720 23112
rect 20675 23072 20720 23100
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 22094 23060 22100 23112
rect 22152 23060 22158 23112
rect 10042 22992 10048 23044
rect 10100 23032 10106 23044
rect 10100 23004 10258 23032
rect 10100 22992 10106 23004
rect 18138 22992 18144 23044
rect 18196 23032 18202 23044
rect 19613 23035 19671 23041
rect 19613 23032 19625 23035
rect 18196 23004 19625 23032
rect 18196 22992 18202 23004
rect 19613 23001 19625 23004
rect 19659 23001 19671 23035
rect 20990 23032 20996 23044
rect 20951 23004 20996 23032
rect 19613 22995 19671 23001
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 22480 22976 22508 23140
rect 24210 23128 24216 23180
rect 24268 23168 24274 23180
rect 25317 23171 25375 23177
rect 25317 23168 25329 23171
rect 24268 23140 25329 23168
rect 24268 23128 24274 23140
rect 25317 23137 25329 23140
rect 25363 23168 25375 23171
rect 25406 23168 25412 23180
rect 25363 23140 25412 23168
rect 25363 23137 25375 23140
rect 25317 23131 25375 23137
rect 25406 23128 25412 23140
rect 25464 23168 25470 23180
rect 30374 23168 30380 23180
rect 25464 23140 29684 23168
rect 25464 23128 25470 23140
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23100 22983 23103
rect 23290 23100 23296 23112
rect 22971 23072 23296 23100
rect 22971 23069 22983 23072
rect 22925 23063 22983 23069
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 25038 23100 25044 23112
rect 24999 23072 25044 23100
rect 25038 23060 25044 23072
rect 25096 23100 25102 23112
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 25096 23072 26249 23100
rect 25096 23060 25102 23072
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 26237 23063 26295 23069
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23069 27123 23103
rect 27065 23063 27123 23069
rect 27893 23103 27951 23109
rect 27893 23069 27905 23103
rect 27939 23100 27951 23103
rect 28534 23100 28540 23112
rect 27939 23072 28540 23100
rect 27939 23069 27951 23072
rect 27893 23063 27951 23069
rect 26605 23035 26663 23041
rect 26605 23001 26617 23035
rect 26651 23032 26663 23035
rect 27080 23032 27108 23063
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 29546 23032 29552 23044
rect 26651 23004 29552 23032
rect 26651 23001 26663 23004
rect 26605 22995 26663 23001
rect 29546 22992 29552 23004
rect 29604 22992 29610 23044
rect 11238 22964 11244 22976
rect 11199 22936 11244 22964
rect 11238 22924 11244 22936
rect 11296 22924 11302 22976
rect 12342 22924 12348 22976
rect 12400 22964 12406 22976
rect 13906 22964 13912 22976
rect 12400 22936 13912 22964
rect 12400 22924 12406 22936
rect 13906 22924 13912 22936
rect 13964 22964 13970 22976
rect 14277 22967 14335 22973
rect 14277 22964 14289 22967
rect 13964 22936 14289 22964
rect 13964 22924 13970 22936
rect 14277 22933 14289 22936
rect 14323 22933 14335 22967
rect 14277 22927 14335 22933
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 16945 22967 17003 22973
rect 16945 22964 16957 22967
rect 16724 22936 16957 22964
rect 16724 22924 16730 22936
rect 16945 22933 16957 22936
rect 16991 22933 17003 22967
rect 17678 22964 17684 22976
rect 17639 22936 17684 22964
rect 16945 22927 17003 22933
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 19300 22936 19441 22964
rect 19300 22924 19306 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 22462 22964 22468 22976
rect 22423 22936 22468 22964
rect 19429 22927 19487 22933
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 27154 22964 27160 22976
rect 27115 22936 27160 22964
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 29656 22964 29684 23140
rect 29748 23140 30380 23168
rect 29748 23109 29776 23140
rect 30374 23128 30380 23140
rect 30432 23128 30438 23180
rect 45005 23171 45063 23177
rect 45005 23137 45017 23171
rect 45051 23168 45063 23171
rect 46750 23168 46756 23180
rect 45051 23140 46756 23168
rect 45051 23137 45063 23140
rect 45005 23131 45063 23137
rect 46750 23128 46756 23140
rect 46808 23128 46814 23180
rect 46842 23128 46848 23180
rect 46900 23168 46906 23180
rect 46900 23140 46945 23168
rect 46900 23128 46906 23140
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 30009 23103 30067 23109
rect 30009 23069 30021 23103
rect 30055 23069 30067 23103
rect 30009 23063 30067 23069
rect 30024 23032 30052 23063
rect 30282 23060 30288 23112
rect 30340 23100 30346 23112
rect 30469 23103 30527 23109
rect 30469 23100 30481 23103
rect 30340 23072 30481 23100
rect 30340 23060 30346 23072
rect 30469 23069 30481 23072
rect 30515 23069 30527 23103
rect 30650 23100 30656 23112
rect 30611 23072 30656 23100
rect 30469 23063 30527 23069
rect 30650 23060 30656 23072
rect 30708 23060 30714 23112
rect 42794 23060 42800 23112
rect 42852 23100 42858 23112
rect 45281 23103 45339 23109
rect 45281 23100 45293 23103
rect 42852 23072 45293 23100
rect 42852 23060 42858 23072
rect 45281 23069 45293 23072
rect 45327 23069 45339 23103
rect 45281 23063 45339 23069
rect 45554 23060 45560 23112
rect 45612 23100 45618 23112
rect 46293 23103 46351 23109
rect 46293 23100 46305 23103
rect 45612 23072 46305 23100
rect 45612 23060 45618 23072
rect 46293 23069 46305 23072
rect 46339 23069 46351 23103
rect 46293 23063 46351 23069
rect 31202 23032 31208 23044
rect 30024 23004 31208 23032
rect 31202 22992 31208 23004
rect 31260 22992 31266 23044
rect 46477 23035 46535 23041
rect 46477 23001 46489 23035
rect 46523 23032 46535 23035
rect 47670 23032 47676 23044
rect 46523 23004 47676 23032
rect 46523 23001 46535 23004
rect 46477 22995 46535 23001
rect 47670 22992 47676 23004
rect 47728 22992 47734 23044
rect 36354 22964 36360 22976
rect 29656 22936 36360 22964
rect 36354 22924 36360 22936
rect 36412 22924 36418 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9769 22763 9827 22769
rect 9769 22760 9781 22763
rect 9548 22732 9781 22760
rect 9548 22720 9554 22732
rect 9769 22729 9781 22732
rect 9815 22729 9827 22763
rect 13998 22760 14004 22772
rect 13959 22732 14004 22760
rect 9769 22723 9827 22729
rect 13998 22720 14004 22732
rect 14056 22720 14062 22772
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 19116 22732 20116 22760
rect 19116 22720 19122 22732
rect 17678 22652 17684 22704
rect 17736 22652 17742 22704
rect 19889 22695 19947 22701
rect 19889 22661 19901 22695
rect 19935 22692 19947 22695
rect 19978 22692 19984 22704
rect 19935 22664 19984 22692
rect 19935 22661 19947 22664
rect 19889 22655 19947 22661
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 20088 22692 20116 22732
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 20809 22763 20867 22769
rect 20809 22760 20821 22763
rect 20772 22732 20821 22760
rect 20772 22720 20778 22732
rect 20809 22729 20821 22732
rect 20855 22729 20867 22763
rect 20809 22723 20867 22729
rect 20990 22720 20996 22772
rect 21048 22760 21054 22772
rect 21913 22763 21971 22769
rect 21913 22760 21925 22763
rect 21048 22732 21925 22760
rect 21048 22720 21054 22732
rect 21913 22729 21925 22732
rect 21959 22729 21971 22763
rect 47670 22760 47676 22772
rect 21913 22723 21971 22729
rect 24872 22732 31754 22760
rect 47631 22732 47676 22760
rect 20088 22664 20208 22692
rect 9674 22624 9680 22636
rect 9635 22596 9680 22624
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 12618 22624 12624 22636
rect 12579 22596 12624 22624
rect 12618 22584 12624 22596
rect 12676 22584 12682 22636
rect 13906 22624 13912 22636
rect 13867 22596 13912 22624
rect 13906 22584 13912 22596
rect 13964 22584 13970 22636
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 15838 22624 15844 22636
rect 15059 22596 15844 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 16666 22624 16672 22636
rect 16627 22596 16672 22624
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 19058 22624 19064 22636
rect 18432 22596 19064 22624
rect 18432 22565 18460 22596
rect 19058 22584 19064 22596
rect 19116 22624 19122 22636
rect 19242 22624 19248 22636
rect 19116 22596 19248 22624
rect 19116 22584 19122 22596
rect 19242 22584 19248 22596
rect 19300 22624 19306 22636
rect 20180 22633 20208 22664
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 24872 22701 24900 22732
rect 24857 22695 24915 22701
rect 20404 22664 22048 22692
rect 20404 22652 20410 22664
rect 20073 22627 20131 22633
rect 20073 22624 20085 22627
rect 19300 22596 20085 22624
rect 19300 22584 19306 22596
rect 20073 22593 20085 22596
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20806 22624 20812 22636
rect 20767 22596 20812 22624
rect 20165 22587 20223 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 22020 22633 22048 22664
rect 24857 22661 24869 22695
rect 24903 22661 24915 22695
rect 27154 22692 27160 22704
rect 27115 22664 27160 22692
rect 24857 22655 24915 22661
rect 27154 22652 27160 22664
rect 27212 22652 27218 22704
rect 31726 22692 31754 22732
rect 47670 22720 47676 22732
rect 47728 22720 47734 22772
rect 37366 22692 37372 22704
rect 31726 22664 37372 22692
rect 37366 22652 37372 22664
rect 37424 22652 37430 22704
rect 45370 22692 45376 22704
rect 45331 22664 45376 22692
rect 45370 22652 45376 22664
rect 45428 22652 45434 22704
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 16945 22559 17003 22565
rect 12759 22528 12848 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 12820 22500 12848 22528
rect 16945 22525 16957 22559
rect 16991 22556 17003 22559
rect 18417 22559 18475 22565
rect 16991 22528 18276 22556
rect 16991 22525 17003 22528
rect 16945 22519 17003 22525
rect 12802 22448 12808 22500
rect 12860 22448 12866 22500
rect 18248 22488 18276 22528
rect 18417 22525 18429 22559
rect 18463 22525 18475 22559
rect 19150 22556 19156 22568
rect 19111 22528 19156 22556
rect 18417 22519 18475 22525
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 21836 22556 21864 22587
rect 22462 22584 22468 22636
rect 22520 22624 22526 22636
rect 23017 22627 23075 22633
rect 23017 22624 23029 22627
rect 22520 22596 23029 22624
rect 22520 22584 22526 22596
rect 23017 22593 23029 22596
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 25038 22584 25044 22636
rect 25096 22624 25102 22636
rect 25317 22627 25375 22633
rect 25317 22624 25329 22627
rect 25096 22596 25329 22624
rect 25096 22584 25102 22596
rect 25317 22593 25329 22596
rect 25363 22593 25375 22627
rect 43438 22624 43444 22636
rect 43399 22596 43444 22624
rect 25317 22587 25375 22593
rect 43438 22584 43444 22596
rect 43496 22584 43502 22636
rect 43714 22624 43720 22636
rect 43675 22596 43720 22624
rect 43714 22584 43720 22596
rect 43772 22584 43778 22636
rect 47578 22624 47584 22636
rect 47539 22596 47584 22624
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 23198 22556 23204 22568
rect 19904 22528 21864 22556
rect 23159 22528 23204 22556
rect 19904 22497 19932 22528
rect 23198 22516 23204 22528
rect 23256 22516 23262 22568
rect 25498 22516 25504 22568
rect 25556 22556 25562 22568
rect 25685 22559 25743 22565
rect 25685 22556 25697 22559
rect 25556 22528 25697 22556
rect 25556 22516 25562 22528
rect 25685 22525 25697 22528
rect 25731 22556 25743 22559
rect 25958 22556 25964 22568
rect 25731 22528 25964 22556
rect 25731 22525 25743 22528
rect 25685 22519 25743 22525
rect 25958 22516 25964 22528
rect 26016 22516 26022 22568
rect 26970 22556 26976 22568
rect 26931 22528 26976 22556
rect 26970 22516 26976 22528
rect 27028 22516 27034 22568
rect 27617 22559 27675 22565
rect 27617 22525 27629 22559
rect 27663 22525 27675 22559
rect 27617 22519 27675 22525
rect 44269 22559 44327 22565
rect 44269 22525 44281 22559
rect 44315 22556 44327 22559
rect 44542 22556 44548 22568
rect 44315 22528 44548 22556
rect 44315 22525 44327 22528
rect 44269 22519 44327 22525
rect 19429 22491 19487 22497
rect 19429 22488 19441 22491
rect 18248 22460 19441 22488
rect 19429 22457 19441 22460
rect 19475 22457 19487 22491
rect 19429 22451 19487 22457
rect 19889 22491 19947 22497
rect 19889 22457 19901 22491
rect 19935 22457 19947 22491
rect 19889 22451 19947 22457
rect 26602 22448 26608 22500
rect 26660 22488 26666 22500
rect 27632 22488 27660 22519
rect 44542 22516 44548 22528
rect 44600 22516 44606 22568
rect 45189 22559 45247 22565
rect 45189 22525 45201 22559
rect 45235 22556 45247 22559
rect 45554 22556 45560 22568
rect 45235 22528 45560 22556
rect 45235 22525 45247 22528
rect 45189 22519 45247 22525
rect 45554 22516 45560 22528
rect 45612 22516 45618 22568
rect 46566 22556 46572 22568
rect 46527 22528 46572 22556
rect 46566 22516 46572 22528
rect 46624 22516 46630 22568
rect 26660 22460 27660 22488
rect 26660 22448 26666 22460
rect 12986 22420 12992 22432
rect 12947 22392 12992 22420
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 15010 22380 15016 22432
rect 15068 22420 15074 22432
rect 15105 22423 15163 22429
rect 15105 22420 15117 22423
rect 15068 22392 15117 22420
rect 15068 22380 15074 22392
rect 15105 22389 15117 22392
rect 15151 22389 15163 22423
rect 15105 22383 15163 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 23198 22216 23204 22228
rect 23159 22188 23204 22216
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 2498 22040 2504 22092
rect 2556 22080 2562 22092
rect 10873 22083 10931 22089
rect 2556 22052 2774 22080
rect 2556 22040 2562 22052
rect 2746 21876 2774 22052
rect 10873 22049 10885 22083
rect 10919 22080 10931 22083
rect 11238 22080 11244 22092
rect 10919 22052 11244 22080
rect 10919 22049 10931 22052
rect 10873 22043 10931 22049
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 15010 22080 15016 22092
rect 14971 22052 15016 22080
rect 15010 22040 15016 22052
rect 15068 22040 15074 22092
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 16224 22052 26065 22080
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 14642 22012 14648 22024
rect 12676 21984 14648 22012
rect 12676 21972 12682 21984
rect 14642 21972 14648 21984
rect 14700 22012 14706 22024
rect 14829 22015 14887 22021
rect 14829 22012 14841 22015
rect 14700 21984 14841 22012
rect 14700 21972 14706 21984
rect 14829 21981 14841 21984
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 11054 21944 11060 21956
rect 11015 21916 11060 21944
rect 11054 21904 11060 21916
rect 11112 21904 11118 21956
rect 12710 21944 12716 21956
rect 12671 21916 12716 21944
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 16224 21876 16252 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 45278 22080 45284 22092
rect 45239 22052 45284 22080
rect 26053 22043 26111 22049
rect 45278 22040 45284 22052
rect 45336 22040 45342 22092
rect 45738 22040 45744 22092
rect 45796 22040 45802 22092
rect 46842 22080 46848 22092
rect 46803 22052 46848 22080
rect 46842 22040 46848 22052
rect 46900 22040 46906 22092
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 16669 22015 16727 22021
rect 16669 22012 16681 22015
rect 16540 21984 16681 22012
rect 16540 21972 16546 21984
rect 16669 21981 16681 21984
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19116 21984 19257 22012
rect 19116 21972 19122 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 20806 21972 20812 22024
rect 20864 22012 20870 22024
rect 21545 22015 21603 22021
rect 21545 22012 21557 22015
rect 20864 21984 21557 22012
rect 20864 21972 20870 21984
rect 21545 21981 21557 21984
rect 21591 21981 21603 22015
rect 21545 21975 21603 21981
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 22012 23167 22015
rect 23290 22012 23296 22024
rect 23155 21984 23296 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 23842 21972 23848 22024
rect 23900 22012 23906 22024
rect 24578 22012 24584 22024
rect 23900 21984 24584 22012
rect 23900 21972 23906 21984
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 25038 22012 25044 22024
rect 24999 21984 25044 22012
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 25869 22015 25927 22021
rect 25869 21981 25881 22015
rect 25915 21981 25927 22015
rect 44174 22012 44180 22024
rect 44135 21984 44180 22012
rect 25869 21975 25927 21981
rect 19426 21944 19432 21956
rect 19387 21916 19432 21944
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 21085 21947 21143 21953
rect 21085 21913 21097 21947
rect 21131 21944 21143 21947
rect 21266 21944 21272 21956
rect 21131 21916 21272 21944
rect 21131 21913 21143 21916
rect 21085 21907 21143 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 25884 21944 25912 21975
rect 44174 21972 44180 21984
rect 44232 21972 44238 22024
rect 44269 22015 44327 22021
rect 44269 21981 44281 22015
rect 44315 22012 44327 22015
rect 44910 22012 44916 22024
rect 44315 21984 44916 22012
rect 44315 21981 44327 21984
rect 44269 21975 44327 21981
rect 44910 21972 44916 21984
rect 44968 21972 44974 22024
rect 45005 22015 45063 22021
rect 45005 21981 45017 22015
rect 45051 22012 45063 22015
rect 45370 22012 45376 22024
rect 45051 21984 45376 22012
rect 45051 21981 45063 21984
rect 45005 21975 45063 21981
rect 45370 21972 45376 21984
rect 45428 21972 45434 22024
rect 26970 21944 26976 21956
rect 25884 21916 26976 21944
rect 26970 21904 26976 21916
rect 27028 21904 27034 21956
rect 27709 21947 27767 21953
rect 27709 21913 27721 21947
rect 27755 21944 27767 21947
rect 28994 21944 29000 21956
rect 27755 21916 29000 21944
rect 27755 21913 27767 21916
rect 27709 21907 27767 21913
rect 28994 21904 29000 21916
rect 29052 21904 29058 21956
rect 40678 21904 40684 21956
rect 40736 21944 40742 21956
rect 45756 21944 45784 22040
rect 46014 21972 46020 22024
rect 46072 22012 46078 22024
rect 46293 22015 46351 22021
rect 46293 22012 46305 22015
rect 46072 21984 46305 22012
rect 46072 21972 46078 21984
rect 46293 21981 46305 21984
rect 46339 21981 46351 22015
rect 46293 21975 46351 21981
rect 40736 21916 45784 21944
rect 46477 21947 46535 21953
rect 40736 21904 40742 21916
rect 46477 21913 46489 21947
rect 46523 21944 46535 21947
rect 47670 21944 47676 21956
rect 46523 21916 47676 21944
rect 46523 21913 46535 21916
rect 46477 21907 46535 21913
rect 47670 21904 47676 21916
rect 47728 21904 47734 21956
rect 2746 21848 16252 21876
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 21637 21879 21695 21885
rect 21637 21876 21649 21879
rect 21416 21848 21649 21876
rect 21416 21836 21422 21848
rect 21637 21845 21649 21848
rect 21683 21845 21695 21879
rect 21637 21839 21695 21845
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25133 21879 25191 21885
rect 25133 21876 25145 21879
rect 25096 21848 25145 21876
rect 25096 21836 25102 21848
rect 25133 21845 25145 21848
rect 25179 21845 25191 21879
rect 25133 21839 25191 21845
rect 43714 21836 43720 21888
rect 43772 21876 43778 21888
rect 43809 21879 43867 21885
rect 43809 21876 43821 21879
rect 43772 21848 43821 21876
rect 43772 21836 43778 21848
rect 43809 21845 43821 21848
rect 43855 21845 43867 21879
rect 44450 21876 44456 21888
rect 44411 21848 44456 21876
rect 43809 21839 43867 21845
rect 44450 21836 44456 21848
rect 44508 21836 44514 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 15381 21675 15439 21681
rect 15381 21672 15393 21675
rect 11112 21644 15393 21672
rect 11112 21632 11118 21644
rect 15381 21641 15393 21644
rect 15427 21641 15439 21675
rect 15381 21635 15439 21641
rect 17696 21644 18276 21672
rect 11974 21604 11980 21616
rect 7944 21576 11980 21604
rect 7944 21545 7972 21576
rect 11974 21564 11980 21576
rect 12032 21564 12038 21616
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 13265 21607 13323 21613
rect 13265 21604 13277 21607
rect 13044 21576 13277 21604
rect 13044 21564 13050 21576
rect 13265 21573 13277 21576
rect 13311 21573 13323 21607
rect 13265 21567 13323 21573
rect 13906 21564 13912 21616
rect 13964 21564 13970 21616
rect 7929 21539 7987 21545
rect 7929 21505 7941 21539
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21505 10471 21539
rect 10413 21499 10471 21505
rect 8113 21471 8171 21477
rect 8113 21437 8125 21471
rect 8159 21468 8171 21471
rect 9030 21468 9036 21480
rect 8159 21440 9036 21468
rect 8159 21437 8171 21440
rect 8113 21431 8171 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 3602 21360 3608 21412
rect 3660 21400 3666 21412
rect 9140 21400 9168 21431
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10428 21468 10456 21499
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 11112 21508 11529 21536
rect 11112 21496 11118 21508
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 11698 21496 11704 21548
rect 11756 21536 11762 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 11756 21508 12173 21536
rect 11756 21496 11762 21508
rect 12161 21505 12173 21508
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 12802 21536 12808 21548
rect 12391 21508 12808 21536
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21536 15347 21539
rect 15654 21536 15660 21548
rect 15335 21508 15660 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 15654 21496 15660 21508
rect 15712 21536 15718 21548
rect 17696 21536 17724 21644
rect 18138 21604 18144 21616
rect 17972 21576 18144 21604
rect 17972 21545 18000 21576
rect 18138 21564 18144 21576
rect 18196 21564 18202 21616
rect 18248 21604 18276 21644
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 20622 21672 20628 21684
rect 20312 21644 20628 21672
rect 20312 21632 20318 21644
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 21913 21675 21971 21681
rect 21913 21641 21925 21675
rect 21959 21672 21971 21675
rect 22094 21672 22100 21684
rect 21959 21644 22100 21672
rect 21959 21641 21971 21644
rect 21913 21635 21971 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 44174 21672 44180 21684
rect 42812 21644 44180 21672
rect 25038 21604 25044 21616
rect 18248 21576 25044 21604
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 25685 21607 25743 21613
rect 25685 21573 25697 21607
rect 25731 21604 25743 21607
rect 40678 21604 40684 21616
rect 25731 21576 40684 21604
rect 25731 21573 25743 21576
rect 25685 21567 25743 21573
rect 40678 21564 40684 21576
rect 40736 21564 40742 21616
rect 15712 21508 17724 21536
rect 17957 21539 18015 21545
rect 15712 21496 15718 21508
rect 17957 21505 17969 21539
rect 18003 21505 18015 21539
rect 20254 21536 20260 21548
rect 20167 21508 20260 21536
rect 17957 21499 18015 21505
rect 20254 21496 20260 21508
rect 20312 21536 20318 21548
rect 20312 21508 20576 21536
rect 20312 21496 20318 21508
rect 12986 21468 12992 21480
rect 9732 21440 12434 21468
rect 12947 21440 12992 21468
rect 9732 21428 9738 21440
rect 3660 21372 9168 21400
rect 12406 21400 12434 21440
rect 12986 21428 12992 21440
rect 13044 21428 13050 21480
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14700 21440 14749 21468
rect 14700 21428 14706 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 18141 21471 18199 21477
rect 18141 21437 18153 21471
rect 18187 21437 18199 21471
rect 18414 21468 18420 21480
rect 18375 21440 18420 21468
rect 18141 21431 18199 21437
rect 12894 21400 12900 21412
rect 12406 21372 12900 21400
rect 3660 21360 3666 21372
rect 12894 21360 12900 21372
rect 12952 21400 12958 21412
rect 18156 21400 18184 21431
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 20349 21403 20407 21409
rect 20349 21400 20361 21403
rect 12952 21372 13124 21400
rect 18156 21372 20361 21400
rect 12952 21360 12958 21372
rect 13096 21344 13124 21372
rect 20349 21369 20361 21372
rect 20395 21369 20407 21403
rect 20548 21400 20576 21508
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21600 21508 21833 21536
rect 21600 21496 21606 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 23109 21539 23167 21545
rect 23109 21505 23121 21539
rect 23155 21536 23167 21539
rect 23474 21536 23480 21548
rect 23155 21508 23480 21536
rect 23155 21505 23167 21508
rect 23109 21499 23167 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 25590 21496 25596 21548
rect 25648 21536 25654 21548
rect 42812 21545 42840 21644
rect 44174 21632 44180 21644
rect 44232 21632 44238 21684
rect 47670 21672 47676 21684
rect 47631 21644 47676 21672
rect 47670 21632 47676 21644
rect 47728 21632 47734 21684
rect 42889 21607 42947 21613
rect 42889 21573 42901 21607
rect 42935 21604 42947 21607
rect 42935 21576 46152 21604
rect 42935 21573 42947 21576
rect 42889 21567 42947 21573
rect 26145 21539 26203 21545
rect 26145 21536 26157 21539
rect 25648 21508 26157 21536
rect 25648 21496 25654 21508
rect 26145 21505 26157 21508
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 42797 21539 42855 21545
rect 42797 21505 42809 21539
rect 42843 21505 42855 21539
rect 42797 21499 42855 21505
rect 42981 21539 43039 21545
rect 42981 21505 42993 21539
rect 43027 21536 43039 21539
rect 43714 21536 43720 21548
rect 43027 21508 43720 21536
rect 43027 21505 43039 21508
rect 42981 21499 43039 21505
rect 43714 21496 43720 21508
rect 43772 21496 43778 21548
rect 44450 21536 44456 21548
rect 44411 21508 44456 21536
rect 44450 21496 44456 21508
rect 44508 21496 44514 21548
rect 44542 21496 44548 21548
rect 44600 21536 44606 21548
rect 44600 21508 44645 21536
rect 44600 21496 44606 21508
rect 44910 21496 44916 21548
rect 44968 21536 44974 21548
rect 45370 21536 45376 21548
rect 44968 21508 45376 21536
rect 44968 21496 44974 21508
rect 45370 21496 45376 21508
rect 45428 21536 45434 21548
rect 46124 21545 46152 21576
rect 45925 21539 45983 21545
rect 45925 21536 45937 21539
rect 45428 21508 45937 21536
rect 45428 21496 45434 21508
rect 45925 21505 45937 21508
rect 45971 21505 45983 21539
rect 45925 21499 45983 21505
rect 46109 21539 46167 21545
rect 46109 21505 46121 21539
rect 46155 21505 46167 21539
rect 47578 21536 47584 21548
rect 47539 21508 47584 21536
rect 46109 21499 46167 21505
rect 47578 21496 47584 21508
rect 47636 21496 47642 21548
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 23845 21471 23903 21477
rect 23845 21468 23857 21471
rect 20772 21440 23857 21468
rect 20772 21428 20778 21440
rect 23124 21412 23152 21440
rect 23845 21437 23857 21440
rect 23891 21437 23903 21471
rect 24026 21468 24032 21480
rect 23987 21440 24032 21468
rect 23845 21431 23903 21437
rect 24026 21428 24032 21440
rect 24084 21428 24090 21480
rect 46845 21471 46903 21477
rect 46845 21437 46857 21471
rect 46891 21437 46903 21471
rect 46845 21431 46903 21437
rect 20548 21372 22094 21400
rect 20349 21363 20407 21369
rect 10226 21332 10232 21344
rect 10187 21304 10232 21332
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 11606 21332 11612 21344
rect 11567 21304 11612 21332
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 12158 21332 12164 21344
rect 12119 21304 12164 21332
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 13078 21292 13084 21344
rect 13136 21292 13142 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 20530 21332 20536 21344
rect 19392 21304 20536 21332
rect 19392 21292 19398 21304
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 22066 21332 22094 21372
rect 23106 21360 23112 21412
rect 23164 21360 23170 21412
rect 26970 21360 26976 21412
rect 27028 21400 27034 21412
rect 44729 21403 44787 21409
rect 44729 21400 44741 21403
rect 27028 21372 44741 21400
rect 27028 21360 27034 21372
rect 44729 21369 44741 21372
rect 44775 21369 44787 21403
rect 44729 21363 44787 21369
rect 46014 21360 46020 21412
rect 46072 21400 46078 21412
rect 46860 21400 46888 21431
rect 46072 21372 46888 21400
rect 46072 21360 46078 21372
rect 23290 21332 23296 21344
rect 22066 21304 23296 21332
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 24762 21292 24768 21344
rect 24820 21332 24826 21344
rect 26329 21335 26387 21341
rect 26329 21332 26341 21335
rect 24820 21304 26341 21332
rect 24820 21292 24826 21304
rect 26329 21301 26341 21304
rect 26375 21301 26387 21335
rect 26329 21295 26387 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 11974 21128 11980 21140
rect 9140 21100 11560 21128
rect 11935 21100 11980 21128
rect 3510 21020 3516 21072
rect 3568 21060 3574 21072
rect 9140 21060 9168 21100
rect 3568 21032 9168 21060
rect 11532 21060 11560 21100
rect 11974 21088 11980 21100
rect 12032 21088 12038 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 13081 21131 13139 21137
rect 13081 21128 13093 21131
rect 13044 21100 13093 21128
rect 13044 21088 13050 21100
rect 13081 21097 13093 21100
rect 13127 21097 13139 21131
rect 13081 21091 13139 21097
rect 19337 21131 19395 21137
rect 19337 21097 19349 21131
rect 19383 21128 19395 21131
rect 19426 21128 19432 21140
rect 19383 21100 19432 21128
rect 19383 21097 19395 21100
rect 19337 21091 19395 21097
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 24026 21128 24032 21140
rect 23799 21100 24032 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 43714 21128 43720 21140
rect 43675 21100 43720 21128
rect 43714 21088 43720 21100
rect 43772 21088 43778 21140
rect 44174 21088 44180 21140
rect 44232 21128 44238 21140
rect 45649 21131 45707 21137
rect 45649 21128 45661 21131
rect 44232 21100 45661 21128
rect 44232 21088 44238 21100
rect 45649 21097 45661 21100
rect 45695 21097 45707 21131
rect 45649 21091 45707 21097
rect 20901 21063 20959 21069
rect 11532 21032 12434 21060
rect 3568 21020 3574 21032
rect 10226 20992 10232 21004
rect 10187 20964 10232 20992
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20992 10563 20995
rect 12158 20992 12164 21004
rect 10551 20964 12164 20992
rect 10551 20961 10563 20964
rect 10505 20955 10563 20961
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 12406 20992 12434 21032
rect 20901 21029 20913 21063
rect 20947 21060 20959 21063
rect 23106 21060 23112 21072
rect 20947 21032 21496 21060
rect 23067 21032 23112 21060
rect 20947 21029 20959 21032
rect 20901 21023 20959 21029
rect 20070 20992 20076 21004
rect 12406 20964 20076 20992
rect 20070 20952 20076 20964
rect 20128 20952 20134 21004
rect 20346 20952 20352 21004
rect 20404 20992 20410 21004
rect 20441 20995 20499 21001
rect 20441 20992 20453 20995
rect 20404 20964 20453 20992
rect 20404 20952 20410 20964
rect 20441 20961 20453 20964
rect 20487 20961 20499 20995
rect 21358 20992 21364 21004
rect 21319 20964 21364 20992
rect 20441 20955 20499 20961
rect 21358 20952 21364 20964
rect 21416 20952 21422 21004
rect 21468 20992 21496 21032
rect 23106 21020 23112 21032
rect 23164 21020 23170 21072
rect 23216 21032 28994 21060
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 21468 20964 21649 20992
rect 21637 20961 21649 20964
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 22922 20952 22928 21004
rect 22980 20992 22986 21004
rect 23216 20992 23244 21032
rect 26602 20992 26608 21004
rect 22980 20964 23244 20992
rect 26563 20964 26608 20992
rect 22980 20952 22986 20964
rect 26602 20952 26608 20964
rect 26660 20952 26666 21004
rect 8478 20884 8484 20936
rect 8536 20924 8542 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8536 20896 8953 20924
rect 8536 20884 8542 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9585 20927 9643 20933
rect 9585 20893 9597 20927
rect 9631 20924 9643 20927
rect 9674 20924 9680 20936
rect 9631 20896 9680 20924
rect 9631 20893 9643 20896
rect 9585 20887 9643 20893
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 13081 20927 13139 20933
rect 13081 20924 13093 20927
rect 12952 20896 13093 20924
rect 12952 20884 12958 20896
rect 13081 20893 13093 20896
rect 13127 20893 13139 20927
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 13081 20887 13139 20893
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 13096 20788 13124 20887
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20924 16819 20927
rect 17770 20924 17776 20936
rect 16807 20896 17776 20924
rect 16807 20893 16819 20896
rect 16761 20887 16819 20893
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 20254 20924 20260 20936
rect 19291 20896 20260 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20924 20591 20927
rect 20714 20924 20720 20936
rect 20579 20896 20720 20924
rect 20579 20893 20591 20896
rect 20533 20887 20591 20893
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 23290 20884 23296 20936
rect 23348 20924 23354 20936
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 23348 20896 23673 20924
rect 23348 20884 23354 20896
rect 23661 20893 23673 20896
rect 23707 20893 23719 20927
rect 24762 20924 24768 20936
rect 24723 20896 24768 20924
rect 23661 20887 23719 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 26145 20927 26203 20933
rect 26145 20893 26157 20927
rect 26191 20893 26203 20927
rect 28966 20924 28994 21032
rect 29362 20952 29368 21004
rect 29420 20992 29426 21004
rect 29733 20995 29791 21001
rect 29733 20992 29745 20995
rect 29420 20964 29745 20992
rect 29420 20952 29426 20964
rect 29733 20961 29745 20964
rect 29779 20961 29791 20995
rect 47210 20992 47216 21004
rect 29733 20955 29791 20961
rect 43640 20964 47216 20992
rect 43640 20933 43668 20964
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 28966 20896 29561 20924
rect 26145 20887 26203 20893
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 43625 20927 43683 20933
rect 43625 20893 43637 20927
rect 43671 20893 43683 20927
rect 43625 20887 43683 20893
rect 43809 20927 43867 20933
rect 43809 20893 43821 20927
rect 43855 20893 43867 20927
rect 43809 20887 43867 20893
rect 13630 20816 13636 20868
rect 13688 20856 13694 20868
rect 13688 20828 16988 20856
rect 13688 20816 13694 20828
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13096 20760 14289 20788
rect 14277 20757 14289 20760
rect 14323 20757 14335 20791
rect 16850 20788 16856 20800
rect 16811 20760 16856 20788
rect 14277 20751 14335 20757
rect 16850 20748 16856 20760
rect 16908 20748 16914 20800
rect 16960 20788 16988 20828
rect 22094 20816 22100 20868
rect 22152 20816 22158 20868
rect 25130 20816 25136 20868
rect 25188 20856 25194 20868
rect 25409 20859 25467 20865
rect 25409 20856 25421 20859
rect 25188 20828 25421 20856
rect 25188 20816 25194 20828
rect 25409 20825 25421 20828
rect 25455 20825 25467 20859
rect 25409 20819 25467 20825
rect 25148 20788 25176 20816
rect 16960 20760 25176 20788
rect 26160 20788 26188 20887
rect 26326 20856 26332 20868
rect 26287 20828 26332 20856
rect 26326 20816 26332 20828
rect 26384 20816 26390 20868
rect 31386 20856 31392 20868
rect 31347 20828 31392 20856
rect 31386 20816 31392 20828
rect 31444 20816 31450 20868
rect 43824 20856 43852 20887
rect 43898 20884 43904 20936
rect 43956 20924 43962 20936
rect 44269 20927 44327 20933
rect 44269 20924 44281 20927
rect 43956 20896 44281 20924
rect 43956 20884 43962 20896
rect 44269 20893 44281 20896
rect 44315 20893 44327 20927
rect 44269 20887 44327 20893
rect 44358 20884 44364 20936
rect 44416 20924 44422 20936
rect 45296 20933 45324 20964
rect 47210 20952 47216 20964
rect 47268 20952 47274 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 44453 20927 44511 20933
rect 44453 20924 44465 20927
rect 44416 20896 44465 20924
rect 44416 20884 44422 20896
rect 44453 20893 44465 20896
rect 44499 20893 44511 20927
rect 44453 20887 44511 20893
rect 45281 20927 45339 20933
rect 45281 20893 45293 20927
rect 45327 20893 45339 20927
rect 46290 20924 46296 20936
rect 46251 20896 46296 20924
rect 45281 20887 45339 20893
rect 46290 20884 46296 20896
rect 46348 20884 46354 20936
rect 44726 20856 44732 20868
rect 43824 20828 44732 20856
rect 44726 20816 44732 20828
rect 44784 20856 44790 20868
rect 45465 20859 45523 20865
rect 45465 20856 45477 20859
rect 44784 20828 45477 20856
rect 44784 20816 44790 20828
rect 45465 20825 45477 20828
rect 45511 20825 45523 20859
rect 45465 20819 45523 20825
rect 46477 20859 46535 20865
rect 46477 20825 46489 20859
rect 46523 20856 46535 20859
rect 47670 20856 47676 20868
rect 46523 20828 47676 20856
rect 46523 20825 46535 20828
rect 46477 20819 46535 20825
rect 47670 20816 47676 20828
rect 47728 20816 47734 20868
rect 28350 20788 28356 20800
rect 26160 20760 28356 20788
rect 28350 20748 28356 20760
rect 28408 20748 28414 20800
rect 44450 20788 44456 20800
rect 44411 20760 44456 20788
rect 44450 20748 44456 20760
rect 44508 20748 44514 20800
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 3786 20544 3792 20596
rect 3844 20584 3850 20596
rect 13081 20587 13139 20593
rect 3844 20556 12112 20584
rect 3844 20544 3850 20556
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 8205 20519 8263 20525
rect 8205 20516 8217 20519
rect 7515 20488 8217 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 8205 20485 8217 20488
rect 8251 20485 8263 20519
rect 8205 20479 8263 20485
rect 11517 20519 11575 20525
rect 11517 20485 11529 20519
rect 11563 20516 11575 20519
rect 11974 20516 11980 20528
rect 11563 20488 11980 20516
rect 11563 20485 11575 20488
rect 11517 20479 11575 20485
rect 11974 20476 11980 20488
rect 12032 20476 12038 20528
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20448 7435 20451
rect 7834 20448 7840 20460
rect 7423 20420 7840 20448
rect 7423 20417 7435 20420
rect 7377 20411 7435 20417
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8570 20380 8576 20392
rect 8067 20352 8432 20380
rect 8531 20352 8576 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8404 20312 8432 20352
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 11716 20380 11744 20411
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12084 20448 12112 20556
rect 13081 20553 13093 20587
rect 13127 20584 13139 20587
rect 13722 20584 13728 20596
rect 13127 20556 13728 20584
rect 13127 20553 13139 20556
rect 13081 20547 13139 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 13906 20584 13912 20596
rect 13867 20556 13912 20584
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 18414 20584 18420 20596
rect 15344 20556 18420 20584
rect 15344 20544 15350 20556
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 20165 20587 20223 20593
rect 20165 20553 20177 20587
rect 20211 20584 20223 20587
rect 20346 20584 20352 20596
rect 20211 20556 20352 20584
rect 20211 20553 20223 20556
rect 20165 20547 20223 20553
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22152 20556 22197 20584
rect 22152 20544 22158 20556
rect 26326 20544 26332 20596
rect 26384 20584 26390 20596
rect 27065 20587 27123 20593
rect 27065 20584 27077 20587
rect 26384 20556 27077 20584
rect 26384 20544 26390 20556
rect 27065 20553 27077 20556
rect 27111 20553 27123 20587
rect 40678 20584 40684 20596
rect 27065 20547 27123 20553
rect 35866 20556 40684 20584
rect 12158 20476 12164 20528
rect 12216 20516 12222 20528
rect 12713 20519 12771 20525
rect 12713 20516 12725 20519
rect 12216 20488 12725 20516
rect 12216 20476 12222 20488
rect 12713 20485 12725 20488
rect 12759 20485 12771 20519
rect 12713 20479 12771 20485
rect 12929 20519 12987 20525
rect 12929 20485 12941 20519
rect 12975 20516 12987 20519
rect 13630 20516 13636 20528
rect 12975 20488 13636 20516
rect 12975 20485 12987 20488
rect 12929 20479 12987 20485
rect 13630 20476 13636 20488
rect 13688 20476 13694 20528
rect 16850 20516 16856 20528
rect 16811 20488 16856 20516
rect 16850 20476 16856 20488
rect 16908 20476 16914 20528
rect 19981 20519 20039 20525
rect 19981 20485 19993 20519
rect 20027 20516 20039 20519
rect 20806 20516 20812 20528
rect 20027 20488 20812 20516
rect 20027 20485 20039 20488
rect 19981 20479 20039 20485
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 25038 20476 25044 20528
rect 25096 20516 25102 20528
rect 25774 20516 25780 20528
rect 25096 20488 25780 20516
rect 25096 20476 25102 20488
rect 25774 20476 25780 20488
rect 25832 20516 25838 20528
rect 27798 20516 27804 20528
rect 25832 20488 27016 20516
rect 27759 20488 27804 20516
rect 25832 20476 25838 20488
rect 11848 20420 11893 20448
rect 12084 20420 13768 20448
rect 11848 20408 11854 20420
rect 11882 20380 11888 20392
rect 11716 20352 11888 20380
rect 11882 20340 11888 20352
rect 11940 20380 11946 20392
rect 11940 20352 12434 20380
rect 11940 20340 11946 20352
rect 11238 20312 11244 20324
rect 8404 20284 11244 20312
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 11517 20315 11575 20321
rect 11517 20281 11529 20315
rect 11563 20312 11575 20315
rect 11698 20312 11704 20324
rect 11563 20284 11704 20312
rect 11563 20281 11575 20284
rect 11517 20275 11575 20281
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 4982 20204 4988 20256
rect 5040 20244 5046 20256
rect 12158 20244 12164 20256
rect 5040 20216 12164 20244
rect 5040 20204 5046 20216
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12406 20244 12434 20352
rect 13740 20312 13768 20420
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 13872 20420 13917 20448
rect 13872 20408 13878 20420
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 14884 20420 15761 20448
rect 14884 20408 14890 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20714 20448 20720 20460
rect 20119 20420 20720 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20714 20408 20720 20420
rect 20772 20448 20778 20460
rect 21082 20448 21088 20460
rect 20772 20420 21088 20448
rect 20772 20408 20778 20420
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 21542 20408 21548 20460
rect 21600 20448 21606 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21600 20420 22017 20448
rect 21600 20408 21606 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 23474 20448 23480 20460
rect 23387 20420 23480 20448
rect 22005 20411 22063 20417
rect 23474 20408 23480 20420
rect 23532 20448 23538 20460
rect 24762 20448 24768 20460
rect 23532 20420 24768 20448
rect 23532 20408 23538 20420
rect 24762 20408 24768 20420
rect 24820 20408 24826 20460
rect 26142 20448 26148 20460
rect 26103 20420 26148 20448
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 26602 20448 26608 20460
rect 26283 20420 26608 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 26988 20457 27016 20488
rect 27798 20476 27804 20488
rect 27856 20476 27862 20528
rect 26973 20451 27031 20457
rect 26973 20417 26985 20451
rect 27019 20417 27031 20451
rect 26973 20411 27031 20417
rect 29546 20408 29552 20460
rect 29604 20448 29610 20460
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 29604 20420 30389 20448
rect 29604 20408 29610 20420
rect 30377 20417 30389 20420
rect 30423 20448 30435 20451
rect 35866 20448 35894 20556
rect 40678 20544 40684 20556
rect 40736 20544 40742 20596
rect 45922 20584 45928 20596
rect 43824 20556 45928 20584
rect 39132 20488 40540 20516
rect 39132 20457 39160 20488
rect 30423 20420 35894 20448
rect 39117 20451 39175 20457
rect 30423 20417 30435 20420
rect 30377 20411 30435 20417
rect 39117 20417 39129 20451
rect 39163 20417 39175 20451
rect 40512 20448 40540 20488
rect 42794 20448 42800 20460
rect 40512 20420 42800 20448
rect 39117 20411 39175 20417
rect 42794 20408 42800 20420
rect 42852 20408 42858 20460
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 16632 20352 16681 20380
rect 16632 20340 16638 20352
rect 16669 20349 16681 20352
rect 16715 20349 16727 20383
rect 16669 20343 16727 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17144 20312 17172 20343
rect 17770 20340 17776 20392
rect 17828 20380 17834 20392
rect 23658 20380 23664 20392
rect 17828 20352 23664 20380
rect 17828 20340 17834 20352
rect 23658 20340 23664 20352
rect 23716 20380 23722 20392
rect 23753 20383 23811 20389
rect 23753 20380 23765 20383
rect 23716 20352 23765 20380
rect 23716 20340 23722 20352
rect 23753 20349 23765 20352
rect 23799 20349 23811 20383
rect 24946 20380 24952 20392
rect 24907 20352 24952 20380
rect 23753 20343 23811 20349
rect 24946 20340 24952 20352
rect 25004 20340 25010 20392
rect 27614 20380 27620 20392
rect 27575 20352 27620 20380
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 28994 20380 29000 20392
rect 28955 20352 29000 20380
rect 28994 20340 29000 20352
rect 29052 20340 29058 20392
rect 31386 20340 31392 20392
rect 31444 20380 31450 20392
rect 39298 20380 39304 20392
rect 31444 20352 39068 20380
rect 39259 20352 39304 20380
rect 31444 20340 31450 20352
rect 13740 20284 17172 20312
rect 19242 20272 19248 20324
rect 19300 20312 19306 20324
rect 19797 20315 19855 20321
rect 19797 20312 19809 20315
rect 19300 20284 19809 20312
rect 19300 20272 19306 20284
rect 19797 20281 19809 20284
rect 19843 20281 19855 20315
rect 22922 20312 22928 20324
rect 19797 20275 19855 20281
rect 19904 20284 22928 20312
rect 12897 20247 12955 20253
rect 12897 20244 12909 20247
rect 12406 20216 12909 20244
rect 12897 20213 12909 20216
rect 12943 20213 12955 20247
rect 15930 20244 15936 20256
rect 15891 20216 15936 20244
rect 12897 20207 12955 20213
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 19904 20244 19932 20284
rect 22922 20272 22928 20284
rect 22980 20272 22986 20324
rect 24964 20312 24992 20340
rect 39040 20312 39068 20352
rect 39298 20340 39304 20352
rect 39356 20340 39362 20392
rect 39577 20383 39635 20389
rect 39577 20349 39589 20383
rect 39623 20349 39635 20383
rect 43824 20380 43852 20556
rect 45922 20544 45928 20556
rect 45980 20544 45986 20596
rect 47670 20584 47676 20596
rect 47631 20556 47676 20584
rect 47670 20544 47676 20556
rect 47728 20544 47734 20596
rect 45373 20519 45431 20525
rect 45373 20485 45385 20519
rect 45419 20516 45431 20519
rect 45462 20516 45468 20528
rect 45419 20488 45468 20516
rect 45419 20485 45431 20488
rect 45373 20479 45431 20485
rect 45462 20476 45468 20488
rect 45520 20476 45526 20528
rect 45738 20476 45744 20528
rect 45796 20516 45802 20528
rect 45796 20488 46980 20516
rect 45796 20476 45802 20488
rect 46952 20460 46980 20488
rect 46934 20408 46940 20460
rect 46992 20448 46998 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 46992 20420 47593 20448
rect 46992 20408 46998 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 39577 20343 39635 20349
rect 41386 20352 43852 20380
rect 39592 20312 39620 20343
rect 24964 20284 35894 20312
rect 39040 20284 39620 20312
rect 17184 20216 19932 20244
rect 17184 20204 17190 20216
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 20349 20247 20407 20253
rect 20349 20244 20361 20247
rect 20036 20216 20361 20244
rect 20036 20204 20042 20216
rect 20349 20213 20361 20216
rect 20395 20213 20407 20247
rect 20349 20207 20407 20213
rect 20530 20204 20536 20256
rect 20588 20244 20594 20256
rect 23014 20244 23020 20256
rect 20588 20216 23020 20244
rect 20588 20204 20594 20216
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 26421 20247 26479 20253
rect 26421 20213 26433 20247
rect 26467 20244 26479 20247
rect 28258 20244 28264 20256
rect 26467 20216 28264 20244
rect 26467 20213 26479 20216
rect 26421 20207 26479 20213
rect 28258 20204 28264 20216
rect 28316 20204 28322 20256
rect 30466 20244 30472 20256
rect 30427 20216 30472 20244
rect 30466 20204 30472 20216
rect 30524 20204 30530 20256
rect 35866 20244 35894 20284
rect 41386 20244 41414 20352
rect 44174 20340 44180 20392
rect 44232 20380 44238 20392
rect 44269 20383 44327 20389
rect 44269 20380 44281 20383
rect 44232 20352 44281 20380
rect 44232 20340 44238 20352
rect 44269 20349 44281 20352
rect 44315 20349 44327 20383
rect 44269 20343 44327 20349
rect 44358 20340 44364 20392
rect 44416 20380 44422 20392
rect 45189 20383 45247 20389
rect 45189 20380 45201 20383
rect 44416 20352 45201 20380
rect 44416 20340 44422 20352
rect 45189 20349 45201 20352
rect 45235 20349 45247 20383
rect 45189 20343 45247 20349
rect 46566 20340 46572 20392
rect 46624 20380 46630 20392
rect 47029 20383 47087 20389
rect 47029 20380 47041 20383
rect 46624 20352 47041 20380
rect 46624 20340 46630 20352
rect 47029 20349 47041 20352
rect 47075 20380 47087 20383
rect 47946 20380 47952 20392
rect 47075 20352 47952 20380
rect 47075 20349 47087 20352
rect 47029 20343 47087 20349
rect 47946 20340 47952 20352
rect 48004 20340 48010 20392
rect 44450 20272 44456 20324
rect 44508 20312 44514 20324
rect 44545 20315 44603 20321
rect 44545 20312 44557 20315
rect 44508 20284 44557 20312
rect 44508 20272 44514 20284
rect 44545 20281 44557 20284
rect 44591 20281 44603 20315
rect 44545 20275 44603 20281
rect 35866 20216 41414 20244
rect 43806 20204 43812 20256
rect 43864 20244 43870 20256
rect 44729 20247 44787 20253
rect 44729 20244 44741 20247
rect 43864 20216 44741 20244
rect 43864 20204 43870 20216
rect 44729 20213 44741 20216
rect 44775 20213 44787 20247
rect 44729 20207 44787 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 9756 20043 9814 20049
rect 9756 20009 9768 20043
rect 9802 20040 9814 20043
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 9802 20012 11713 20040
rect 9802 20009 9814 20012
rect 9756 20003 9814 20009
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 15286 20040 15292 20052
rect 12032 20012 15292 20040
rect 12032 20000 12038 20012
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 17126 20040 17132 20052
rect 15396 20012 17132 20040
rect 1762 19932 1768 19984
rect 1820 19972 1826 19984
rect 15396 19972 15424 20012
rect 17126 20000 17132 20012
rect 17184 20000 17190 20052
rect 26602 20040 26608 20052
rect 17236 20012 22094 20040
rect 26563 20012 26608 20040
rect 1820 19944 2774 19972
rect 1820 19932 1826 19944
rect 2746 19904 2774 19944
rect 10796 19944 15424 19972
rect 10796 19904 10824 19944
rect 11238 19904 11244 19916
rect 2746 19876 10824 19904
rect 11199 19876 11244 19904
rect 11238 19864 11244 19876
rect 11296 19904 11302 19916
rect 11296 19876 12112 19904
rect 11296 19864 11302 19876
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19805 9551 19839
rect 9493 19799 9551 19805
rect 9508 19768 9536 19799
rect 10870 19796 10876 19848
rect 10928 19796 10934 19848
rect 11882 19836 11888 19848
rect 11843 19808 11888 19836
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 11974 19796 11980 19848
rect 12032 19796 12038 19848
rect 12084 19836 12112 19876
rect 12158 19864 12164 19916
rect 12216 19904 12222 19916
rect 17236 19904 17264 20012
rect 12216 19876 17264 19904
rect 19521 19907 19579 19913
rect 12216 19864 12222 19876
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20530 19904 20536 19916
rect 19567 19876 20536 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 12084 19808 12265 19836
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14826 19836 14832 19848
rect 14139 19808 14832 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 9674 19768 9680 19780
rect 9508 19740 9680 19768
rect 9674 19728 9680 19740
rect 9732 19728 9738 19780
rect 11992 19768 12020 19796
rect 11072 19740 12020 19768
rect 3970 19660 3976 19712
rect 4028 19700 4034 19712
rect 11072 19700 11100 19740
rect 12158 19728 12164 19780
rect 12216 19768 12222 19780
rect 12360 19768 12388 19799
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 16666 19796 16672 19848
rect 16724 19796 16730 19848
rect 17770 19836 17776 19848
rect 17731 19808 17776 19836
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 21542 19836 21548 19848
rect 19245 19799 19303 19805
rect 20824 19808 21548 19836
rect 15562 19768 15568 19780
rect 12216 19740 12388 19768
rect 15523 19740 15568 19768
rect 12216 19728 12222 19740
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 19260 19768 19288 19799
rect 19426 19768 19432 19780
rect 19260 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 4028 19672 11100 19700
rect 4028 19660 4034 19672
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11848 19672 11897 19700
rect 11848 19660 11854 19672
rect 11885 19669 11897 19672
rect 11931 19700 11943 19703
rect 11974 19700 11980 19712
rect 11931 19672 11980 19700
rect 11931 19669 11943 19672
rect 11885 19663 11943 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 13814 19700 13820 19712
rect 12308 19672 13820 19700
rect 12308 19660 12314 19672
rect 13814 19660 13820 19672
rect 13872 19700 13878 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 13872 19672 14289 19700
rect 13872 19660 13878 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14277 19663 14335 19669
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 16574 19700 16580 19712
rect 15804 19672 16580 19700
rect 15804 19660 15810 19672
rect 16574 19660 16580 19672
rect 16632 19700 16638 19712
rect 17037 19703 17095 19709
rect 17037 19700 17049 19703
rect 16632 19672 17049 19700
rect 16632 19660 16638 19672
rect 17037 19669 17049 19672
rect 17083 19669 17095 19703
rect 17862 19700 17868 19712
rect 17823 19672 17868 19700
rect 17037 19663 17095 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 18046 19660 18052 19712
rect 18104 19700 18110 19712
rect 20824 19700 20852 19808
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 22066 19836 22094 20012
rect 26602 20000 26608 20012
rect 26660 20000 26666 20052
rect 31386 19972 31392 19984
rect 26436 19944 31392 19972
rect 26436 19904 26464 19944
rect 31386 19932 31392 19944
rect 31444 19932 31450 19984
rect 44174 19932 44180 19984
rect 44232 19972 44238 19984
rect 44232 19944 45600 19972
rect 44232 19932 44238 19944
rect 27798 19904 27804 19916
rect 24596 19876 26464 19904
rect 24596 19845 24624 19876
rect 26436 19848 26464 19876
rect 27632 19876 27804 19904
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 22066 19808 24409 19836
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24412 19768 24440 19799
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 25133 19839 25191 19845
rect 25133 19836 25145 19839
rect 24820 19808 25145 19836
rect 24820 19796 24826 19808
rect 25133 19805 25145 19808
rect 25179 19805 25191 19839
rect 26237 19839 26295 19845
rect 26237 19836 26249 19839
rect 25133 19799 25191 19805
rect 25332 19808 26249 19836
rect 25332 19780 25360 19808
rect 26237 19805 26249 19808
rect 26283 19805 26295 19839
rect 26237 19799 26295 19805
rect 26418 19796 26424 19848
rect 26476 19836 26482 19848
rect 27430 19836 27436 19848
rect 26476 19808 26569 19836
rect 27391 19808 27436 19836
rect 26476 19796 26482 19808
rect 27430 19796 27436 19808
rect 27488 19796 27494 19848
rect 27632 19845 27660 19876
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 30466 19904 30472 19916
rect 30427 19876 30472 19904
rect 30466 19864 30472 19876
rect 30524 19864 30530 19916
rect 40589 19907 40647 19913
rect 40589 19873 40601 19907
rect 40635 19904 40647 19907
rect 44358 19904 44364 19916
rect 40635 19876 44364 19904
rect 40635 19873 40647 19876
rect 40589 19867 40647 19873
rect 44358 19864 44364 19876
rect 44416 19864 44422 19916
rect 44450 19864 44456 19916
rect 44508 19904 44514 19916
rect 44508 19876 45232 19904
rect 44508 19864 44514 19876
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19805 27675 19839
rect 28258 19836 28264 19848
rect 28219 19808 28264 19836
rect 27617 19799 27675 19805
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 30285 19839 30343 19845
rect 30285 19805 30297 19839
rect 30331 19805 30343 19839
rect 43806 19836 43812 19848
rect 43767 19808 43812 19836
rect 30285 19799 30343 19805
rect 25314 19768 25320 19780
rect 24412 19740 25320 19768
rect 25314 19728 25320 19740
rect 25372 19728 25378 19780
rect 25406 19728 25412 19780
rect 25464 19768 25470 19780
rect 25501 19771 25559 19777
rect 25501 19768 25513 19771
rect 25464 19740 25513 19768
rect 25464 19728 25470 19740
rect 25501 19737 25513 19740
rect 25547 19737 25559 19771
rect 25501 19731 25559 19737
rect 27709 19771 27767 19777
rect 27709 19737 27721 19771
rect 27755 19768 27767 19771
rect 27798 19768 27804 19780
rect 27755 19740 27804 19768
rect 27755 19737 27767 19740
rect 27709 19731 27767 19737
rect 27798 19728 27804 19740
rect 27856 19728 27862 19780
rect 30300 19768 30328 19799
rect 43806 19796 43812 19808
rect 43864 19796 43870 19848
rect 44085 19839 44143 19845
rect 44085 19805 44097 19839
rect 44131 19836 44143 19839
rect 44818 19836 44824 19848
rect 44131 19808 44824 19836
rect 44131 19805 44143 19808
rect 44085 19799 44143 19805
rect 44818 19796 44824 19808
rect 44876 19836 44882 19848
rect 45204 19845 45232 19876
rect 45370 19864 45376 19916
rect 45428 19904 45434 19916
rect 45572 19913 45600 19944
rect 45465 19907 45523 19913
rect 45465 19904 45477 19907
rect 45428 19876 45477 19904
rect 45428 19864 45434 19876
rect 45465 19873 45477 19876
rect 45511 19873 45523 19907
rect 45465 19867 45523 19873
rect 45557 19907 45615 19913
rect 45557 19873 45569 19907
rect 45603 19873 45615 19907
rect 45557 19867 45615 19873
rect 46477 19907 46535 19913
rect 46477 19873 46489 19907
rect 46523 19904 46535 19907
rect 48038 19904 48044 19916
rect 46523 19876 48044 19904
rect 46523 19873 46535 19876
rect 46477 19867 46535 19873
rect 48038 19864 48044 19876
rect 48096 19864 48102 19916
rect 45005 19839 45063 19845
rect 45005 19836 45017 19839
rect 44876 19808 45017 19836
rect 44876 19796 44882 19808
rect 45005 19805 45017 19808
rect 45051 19805 45063 19839
rect 45005 19799 45063 19805
rect 45189 19839 45247 19845
rect 45189 19805 45201 19839
rect 45235 19805 45247 19839
rect 45189 19799 45247 19805
rect 46293 19839 46351 19845
rect 46293 19805 46305 19839
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 31938 19768 31944 19780
rect 30300 19740 31944 19768
rect 31938 19728 31944 19740
rect 31996 19728 32002 19780
rect 32122 19768 32128 19780
rect 32083 19740 32128 19768
rect 32122 19728 32128 19740
rect 32180 19728 32186 19780
rect 40770 19768 40776 19780
rect 40731 19740 40776 19768
rect 40770 19728 40776 19740
rect 40828 19728 40834 19780
rect 42426 19768 42432 19780
rect 42387 19740 42432 19768
rect 42426 19728 42432 19740
rect 42484 19728 42490 19780
rect 46308 19768 46336 19799
rect 43824 19740 46336 19768
rect 20990 19700 20996 19712
rect 18104 19672 20852 19700
rect 20951 19672 20996 19700
rect 18104 19660 18110 19672
rect 20990 19660 20996 19672
rect 21048 19660 21054 19712
rect 21542 19660 21548 19712
rect 21600 19700 21606 19712
rect 21637 19703 21695 19709
rect 21637 19700 21649 19703
rect 21600 19672 21649 19700
rect 21600 19660 21606 19672
rect 21637 19669 21649 19672
rect 21683 19669 21695 19703
rect 21637 19663 21695 19669
rect 24581 19703 24639 19709
rect 24581 19669 24593 19703
rect 24627 19700 24639 19703
rect 26142 19700 26148 19712
rect 24627 19672 26148 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 26142 19660 26148 19672
rect 26200 19660 26206 19712
rect 28350 19700 28356 19712
rect 28311 19672 28356 19700
rect 28350 19660 28356 19672
rect 28408 19660 28414 19712
rect 40586 19660 40592 19712
rect 40644 19700 40650 19712
rect 43824 19700 43852 19740
rect 48038 19728 48044 19780
rect 48096 19768 48102 19780
rect 48133 19771 48191 19777
rect 48133 19768 48145 19771
rect 48096 19740 48145 19768
rect 48096 19728 48102 19740
rect 48133 19737 48145 19740
rect 48179 19737 48191 19771
rect 48133 19731 48191 19737
rect 40644 19672 43852 19700
rect 40644 19660 40650 19672
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 10870 19496 10876 19508
rect 10831 19468 10876 19496
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11882 19496 11888 19508
rect 11843 19468 11888 19496
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 16761 19499 16819 19505
rect 16761 19496 16773 19499
rect 16724 19468 16773 19496
rect 16724 19456 16730 19468
rect 16761 19465 16773 19468
rect 16807 19465 16819 19499
rect 19242 19496 19248 19508
rect 16761 19459 16819 19465
rect 17696 19468 19248 19496
rect 11238 19388 11244 19440
rect 11296 19428 11302 19440
rect 11517 19431 11575 19437
rect 11517 19428 11529 19431
rect 11296 19400 11529 19428
rect 11296 19388 11302 19400
rect 11517 19397 11529 19400
rect 11563 19397 11575 19431
rect 11517 19391 11575 19397
rect 11733 19431 11791 19437
rect 11733 19397 11745 19431
rect 11779 19428 11791 19431
rect 11779 19400 11928 19428
rect 11779 19397 11791 19400
rect 11733 19391 11791 19397
rect 11900 19372 11928 19400
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 11054 19360 11060 19372
rect 10827 19332 11060 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12342 19360 12348 19372
rect 12303 19332 12348 19360
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12529 19363 12587 19369
rect 12529 19360 12541 19363
rect 12452 19332 12541 19360
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 12452 19292 12480 19332
rect 12529 19329 12541 19332
rect 12575 19329 12587 19363
rect 15746 19360 15752 19372
rect 15707 19332 15752 19360
rect 12529 19323 12587 19329
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 17696 19369 17724 19468
rect 19242 19456 19248 19468
rect 19300 19496 19306 19508
rect 20990 19496 20996 19508
rect 19300 19468 20996 19496
rect 19300 19456 19306 19468
rect 17862 19428 17868 19440
rect 17823 19400 17868 19428
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15988 19332 16681 19360
rect 15988 19320 15994 19332
rect 16669 19329 16681 19332
rect 16715 19360 16727 19363
rect 17681 19363 17739 19369
rect 16715 19332 17632 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 12216 19264 12480 19292
rect 15841 19295 15899 19301
rect 12216 19252 12222 19264
rect 15841 19261 15853 19295
rect 15887 19292 15899 19295
rect 16022 19292 16028 19304
rect 15887 19264 16028 19292
rect 15887 19261 15899 19264
rect 15841 19255 15899 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 17604 19292 17632 19332
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 20158 19363 20216 19369
rect 20158 19329 20170 19363
rect 20204 19358 20216 19363
rect 20272 19358 20300 19468
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21082 19456 21088 19508
rect 21140 19496 21146 19508
rect 21177 19499 21235 19505
rect 21177 19496 21189 19499
rect 21140 19468 21189 19496
rect 21140 19456 21146 19468
rect 21177 19465 21189 19468
rect 21223 19465 21235 19499
rect 21177 19459 21235 19465
rect 27614 19456 27620 19508
rect 27672 19496 27678 19508
rect 28074 19496 28080 19508
rect 27672 19468 28080 19496
rect 27672 19456 27678 19468
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 31938 19456 31944 19508
rect 31996 19496 32002 19508
rect 40586 19496 40592 19508
rect 31996 19468 40592 19496
rect 31996 19456 32002 19468
rect 40586 19456 40592 19468
rect 40644 19456 40650 19508
rect 40770 19496 40776 19508
rect 40731 19468 40776 19496
rect 40770 19456 40776 19468
rect 40828 19456 40834 19508
rect 44082 19456 44088 19508
rect 44140 19496 44146 19508
rect 45830 19496 45836 19508
rect 44140 19468 45836 19496
rect 44140 19456 44146 19468
rect 45830 19456 45836 19468
rect 45888 19496 45894 19508
rect 46474 19496 46480 19508
rect 45888 19468 46480 19496
rect 45888 19456 45894 19468
rect 46474 19456 46480 19468
rect 46532 19456 46538 19508
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 21818 19428 21824 19440
rect 20404 19400 21312 19428
rect 21779 19400 21824 19428
rect 20404 19388 20410 19400
rect 20204 19330 20300 19358
rect 20204 19329 20216 19330
rect 20158 19323 20216 19329
rect 20806 19320 20812 19372
rect 20864 19360 20870 19372
rect 21284 19369 21312 19400
rect 21818 19388 21824 19400
rect 21876 19388 21882 19440
rect 23014 19428 23020 19440
rect 22051 19397 22109 19403
rect 22975 19400 23020 19428
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20864 19332 21005 19360
rect 20864 19320 20870 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22051 19363 22063 19397
rect 22097 19363 22109 19397
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 43254 19428 43260 19440
rect 35866 19400 43260 19428
rect 22051 19360 22109 19363
rect 25222 19360 25228 19372
rect 21315 19357 22109 19360
rect 21315 19332 22094 19357
rect 25183 19332 25228 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 18046 19292 18052 19304
rect 17604 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19261 18291 19295
rect 18233 19255 18291 19261
rect 20257 19295 20315 19301
rect 20257 19261 20269 19295
rect 20303 19261 20315 19295
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 20257 19255 20315 19261
rect 3418 19184 3424 19236
rect 3476 19224 3482 19236
rect 3476 19196 15516 19224
rect 3476 19184 3482 19196
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 11790 19156 11796 19168
rect 11747 19128 11796 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 12894 19156 12900 19168
rect 12391 19128 12900 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 15488 19156 15516 19196
rect 15562 19184 15568 19236
rect 15620 19224 15626 19236
rect 16117 19227 16175 19233
rect 16117 19224 16129 19227
rect 15620 19196 16129 19224
rect 15620 19184 15626 19196
rect 16117 19193 16129 19196
rect 16163 19193 16175 19227
rect 16117 19187 16175 19193
rect 18248 19156 18276 19255
rect 20272 19224 20300 19255
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 21008 19292 21036 19323
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 25314 19320 25320 19372
rect 25372 19360 25378 19372
rect 25961 19363 26019 19369
rect 25372 19332 25417 19360
rect 25372 19320 25378 19332
rect 25961 19329 25973 19363
rect 26007 19360 26019 19363
rect 26418 19360 26424 19372
rect 26007 19332 26424 19360
rect 26007 19329 26019 19332
rect 25961 19323 26019 19329
rect 26418 19320 26424 19332
rect 26476 19320 26482 19372
rect 27709 19363 27767 19369
rect 27709 19329 27721 19363
rect 27755 19360 27767 19363
rect 28442 19360 28448 19372
rect 27755 19332 28448 19360
rect 27755 19329 27767 19332
rect 27709 19323 27767 19329
rect 21818 19292 21824 19304
rect 21008 19264 21824 19292
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22922 19292 22928 19304
rect 22883 19264 22928 19292
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 23750 19292 23756 19304
rect 23711 19264 23756 19292
rect 23750 19252 23756 19264
rect 23808 19252 23814 19304
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 26053 19295 26111 19301
rect 26053 19292 26065 19295
rect 24912 19264 26065 19292
rect 24912 19252 24918 19264
rect 26053 19261 26065 19264
rect 26099 19261 26111 19295
rect 26053 19255 26111 19261
rect 26329 19295 26387 19301
rect 26329 19261 26341 19295
rect 26375 19292 26387 19295
rect 27724 19292 27752 19323
rect 28442 19320 28448 19332
rect 28500 19360 28506 19372
rect 28629 19363 28687 19369
rect 28629 19360 28641 19363
rect 28500 19332 28641 19360
rect 28500 19320 28506 19332
rect 28629 19329 28641 19332
rect 28675 19329 28687 19363
rect 28629 19323 28687 19329
rect 28718 19320 28724 19372
rect 28776 19360 28782 19372
rect 28905 19363 28963 19369
rect 28905 19360 28917 19363
rect 28776 19332 28917 19360
rect 28776 19320 28782 19332
rect 28905 19329 28917 19332
rect 28951 19329 28963 19363
rect 28905 19323 28963 19329
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19360 29791 19363
rect 35866 19360 35894 19400
rect 43254 19388 43260 19400
rect 43312 19388 43318 19440
rect 47578 19428 47584 19440
rect 43732 19400 47584 19428
rect 40678 19360 40684 19372
rect 29779 19332 35894 19360
rect 40639 19332 40684 19360
rect 29779 19329 29791 19332
rect 29733 19323 29791 19329
rect 40678 19320 40684 19332
rect 40736 19360 40742 19372
rect 43732 19360 43760 19400
rect 47578 19388 47584 19400
rect 47636 19388 47642 19440
rect 43898 19360 43904 19372
rect 40736 19332 43760 19360
rect 43859 19332 43904 19360
rect 40736 19320 40742 19332
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 44082 19360 44088 19372
rect 44043 19332 44088 19360
rect 44082 19320 44088 19332
rect 44140 19320 44146 19372
rect 44174 19320 44180 19372
rect 44232 19320 44238 19372
rect 45002 19360 45008 19372
rect 44963 19332 45008 19360
rect 45002 19320 45008 19332
rect 45060 19320 45066 19372
rect 26375 19264 27752 19292
rect 27801 19295 27859 19301
rect 26375 19261 26387 19264
rect 26329 19255 26387 19261
rect 27801 19261 27813 19295
rect 27847 19292 27859 19295
rect 27982 19292 27988 19304
rect 27847 19264 27988 19292
rect 27847 19261 27859 19264
rect 27801 19255 27859 19261
rect 27982 19252 27988 19264
rect 28040 19252 28046 19304
rect 28810 19252 28816 19304
rect 28868 19292 28874 19304
rect 29365 19295 29423 19301
rect 29365 19292 29377 19295
rect 28868 19264 29377 19292
rect 28868 19252 28874 19264
rect 29365 19261 29377 19264
rect 29411 19261 29423 19295
rect 29365 19255 29423 19261
rect 43993 19295 44051 19301
rect 43993 19261 44005 19295
rect 44039 19292 44051 19295
rect 44192 19292 44220 19320
rect 44039 19264 44220 19292
rect 44039 19261 44051 19264
rect 43993 19255 44051 19261
rect 44266 19252 44272 19304
rect 44324 19292 44330 19304
rect 44729 19295 44787 19301
rect 44729 19292 44741 19295
rect 44324 19264 44741 19292
rect 44324 19252 44330 19264
rect 44729 19261 44741 19264
rect 44775 19261 44787 19295
rect 45554 19292 45560 19304
rect 45515 19264 45560 19292
rect 44729 19255 44787 19261
rect 45554 19252 45560 19264
rect 45612 19252 45618 19304
rect 46290 19252 46296 19304
rect 46348 19292 46354 19304
rect 47765 19295 47823 19301
rect 47765 19292 47777 19295
rect 46348 19264 47777 19292
rect 46348 19252 46354 19264
rect 47765 19261 47777 19264
rect 47811 19261 47823 19295
rect 47765 19255 47823 19261
rect 20714 19224 20720 19236
rect 20272 19196 20720 19224
rect 20714 19184 20720 19196
rect 20772 19224 20778 19236
rect 22189 19227 22247 19233
rect 22189 19224 22201 19227
rect 20772 19196 22201 19224
rect 20772 19184 20778 19196
rect 22189 19193 22201 19196
rect 22235 19193 22247 19227
rect 22189 19187 22247 19193
rect 30009 19227 30067 19233
rect 30009 19193 30021 19227
rect 30055 19224 30067 19227
rect 44174 19224 44180 19236
rect 30055 19196 44180 19224
rect 30055 19193 30067 19196
rect 30009 19187 30067 19193
rect 44174 19184 44180 19196
rect 44232 19184 44238 19236
rect 20990 19156 20996 19168
rect 15488 19128 18276 19156
rect 20951 19128 20996 19156
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21140 19128 22017 19156
rect 21140 19116 21146 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 46290 19116 46296 19168
rect 46348 19156 46354 19168
rect 47029 19159 47087 19165
rect 47029 19156 47041 19159
rect 46348 19128 47041 19156
rect 46348 19116 46354 19128
rect 47029 19125 47041 19128
rect 47075 19125 47087 19159
rect 47029 19119 47087 19125
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2004 18924 2329 18952
rect 2004 18912 2010 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 11977 18955 12035 18961
rect 11977 18952 11989 18955
rect 11940 18924 11989 18952
rect 11940 18912 11946 18924
rect 11977 18921 11989 18924
rect 12023 18921 12035 18955
rect 12158 18952 12164 18964
rect 12119 18924 12164 18952
rect 11977 18915 12035 18921
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13688 18924 14289 18952
rect 13688 18912 13694 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 15749 18955 15807 18961
rect 15749 18952 15761 18955
rect 15344 18924 15761 18952
rect 15344 18912 15350 18924
rect 15749 18921 15761 18924
rect 15795 18921 15807 18955
rect 19426 18952 19432 18964
rect 19387 18924 19432 18952
rect 15749 18915 15807 18921
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 22281 18955 22339 18961
rect 22281 18952 22293 18955
rect 21876 18924 22293 18952
rect 21876 18912 21882 18924
rect 22281 18921 22293 18924
rect 22327 18921 22339 18955
rect 27982 18952 27988 18964
rect 27943 18924 27988 18952
rect 22281 18915 22339 18921
rect 27982 18912 27988 18924
rect 28040 18912 28046 18964
rect 31938 18952 31944 18964
rect 31899 18924 31944 18952
rect 31938 18912 31944 18924
rect 31996 18912 32002 18964
rect 44266 18952 44272 18964
rect 44227 18924 44272 18952
rect 44266 18912 44272 18924
rect 44324 18912 44330 18964
rect 14461 18887 14519 18893
rect 14461 18853 14473 18887
rect 14507 18853 14519 18887
rect 14461 18847 14519 18853
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12897 18819 12955 18825
rect 12897 18816 12909 18819
rect 12032 18788 12909 18816
rect 12032 18776 12038 18788
rect 12897 18785 12909 18788
rect 12943 18785 12955 18819
rect 14476 18816 14504 18847
rect 16022 18844 16028 18896
rect 16080 18884 16086 18896
rect 19978 18884 19984 18896
rect 16080 18856 19984 18884
rect 16080 18844 16086 18856
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 23845 18887 23903 18893
rect 23845 18853 23857 18887
rect 23891 18884 23903 18887
rect 24854 18884 24860 18896
rect 23891 18856 24860 18884
rect 23891 18853 23903 18856
rect 23845 18847 23903 18853
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 27798 18884 27804 18896
rect 27759 18856 27804 18884
rect 27798 18844 27804 18856
rect 27856 18844 27862 18896
rect 43349 18887 43407 18893
rect 43349 18884 43361 18887
rect 35866 18856 43361 18884
rect 23477 18819 23535 18825
rect 12897 18779 12955 18785
rect 13464 18788 14504 18816
rect 15764 18788 19380 18816
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 2314 18748 2320 18760
rect 2271 18720 2320 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 2314 18708 2320 18720
rect 2372 18748 2378 18760
rect 7558 18748 7564 18760
rect 2372 18720 7564 18748
rect 2372 18708 2378 18720
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 11054 18748 11060 18760
rect 11015 18720 11060 18748
rect 11054 18708 11060 18720
rect 11112 18748 11118 18760
rect 12250 18748 12256 18760
rect 11112 18720 12256 18748
rect 11112 18708 11118 18720
rect 12250 18708 12256 18720
rect 12308 18748 12314 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 12308 18720 13369 18748
rect 12308 18708 12314 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 11790 18680 11796 18692
rect 11751 18652 11796 18680
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 12009 18683 12067 18689
rect 12009 18649 12021 18683
rect 12055 18680 12067 18683
rect 12713 18683 12771 18689
rect 12713 18680 12725 18683
rect 12055 18652 12725 18680
rect 12055 18649 12067 18652
rect 12009 18643 12067 18649
rect 12713 18649 12725 18652
rect 12759 18680 12771 18683
rect 13464 18680 13492 18788
rect 15764 18760 15792 18788
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 14921 18751 14979 18757
rect 14921 18748 14933 18751
rect 14884 18720 14933 18748
rect 14884 18708 14890 18720
rect 14921 18717 14933 18720
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 15746 18748 15752 18760
rect 15703 18720 15752 18748
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 17586 18748 17592 18760
rect 17547 18720 17592 18748
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 19352 18757 19380 18788
rect 23477 18785 23489 18819
rect 23523 18816 23535 18819
rect 23750 18816 23756 18828
rect 23523 18788 23756 18816
rect 23523 18785 23535 18788
rect 23477 18779 23535 18785
rect 23750 18776 23756 18788
rect 23808 18816 23814 18828
rect 23808 18788 24532 18816
rect 23808 18776 23814 18788
rect 24504 18760 24532 18788
rect 25222 18776 25228 18828
rect 25280 18816 25286 18828
rect 26053 18819 26111 18825
rect 26053 18816 26065 18819
rect 25280 18788 26065 18816
rect 25280 18776 25286 18788
rect 26053 18785 26065 18788
rect 26099 18785 26111 18819
rect 28442 18816 28448 18828
rect 28403 18788 28448 18816
rect 26053 18779 26111 18785
rect 28442 18776 28448 18788
rect 28500 18776 28506 18828
rect 19337 18751 19395 18757
rect 19337 18717 19349 18751
rect 19383 18748 19395 18751
rect 19426 18748 19432 18760
rect 19383 18720 19432 18748
rect 19383 18717 19395 18720
rect 19337 18711 19395 18717
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20036 18720 20545 18748
rect 20036 18708 20042 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 24486 18748 24492 18760
rect 24447 18720 24492 18748
rect 23661 18711 23719 18717
rect 12759 18652 13492 18680
rect 12759 18649 12771 18652
rect 12713 18643 12771 18649
rect 13906 18640 13912 18692
rect 13964 18680 13970 18692
rect 14093 18683 14151 18689
rect 14093 18680 14105 18683
rect 13964 18652 14105 18680
rect 13964 18640 13970 18652
rect 14093 18649 14105 18652
rect 14139 18680 14151 18683
rect 14550 18680 14556 18692
rect 14139 18652 14556 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 18230 18680 18236 18692
rect 18191 18652 18236 18680
rect 18230 18640 18236 18652
rect 18288 18680 18294 18692
rect 20806 18680 20812 18692
rect 18288 18652 20668 18680
rect 20767 18652 20812 18680
rect 18288 18640 18294 18652
rect 20640 18624 20668 18652
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 21542 18640 21548 18692
rect 21600 18640 21606 18692
rect 23676 18680 23704 18711
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 26142 18748 26148 18760
rect 26103 18720 26148 18748
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 27525 18751 27583 18757
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 27614 18748 27620 18760
rect 27571 18720 27620 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 27614 18708 27620 18720
rect 27672 18748 27678 18760
rect 28629 18751 28687 18757
rect 28629 18748 28641 18751
rect 27672 18720 28641 18748
rect 27672 18708 27678 18720
rect 28629 18717 28641 18720
rect 28675 18748 28687 18751
rect 28718 18748 28724 18760
rect 28675 18720 28724 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 28718 18708 28724 18720
rect 28776 18708 28782 18760
rect 28905 18751 28963 18757
rect 28905 18717 28917 18751
rect 28951 18748 28963 18751
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 28951 18720 30113 18748
rect 28951 18717 28963 18720
rect 28905 18711 28963 18717
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18748 31079 18751
rect 35866 18748 35894 18856
rect 43349 18853 43361 18856
rect 43395 18853 43407 18887
rect 43349 18847 43407 18853
rect 45097 18887 45155 18893
rect 45097 18853 45109 18887
rect 45143 18853 45155 18887
rect 45097 18847 45155 18853
rect 45112 18816 45140 18847
rect 46290 18816 46296 18828
rect 43272 18788 45140 18816
rect 46251 18788 46296 18816
rect 43272 18760 43300 18788
rect 46290 18776 46296 18788
rect 46348 18776 46354 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 43254 18748 43260 18760
rect 31067 18720 35894 18748
rect 43215 18720 43260 18748
rect 31067 18717 31079 18720
rect 31021 18711 31079 18717
rect 43254 18708 43260 18720
rect 43312 18708 43318 18760
rect 43533 18751 43591 18757
rect 43533 18717 43545 18751
rect 43579 18717 43591 18751
rect 44174 18748 44180 18760
rect 44135 18720 44180 18748
rect 43533 18711 43591 18717
rect 24688 18680 24716 18708
rect 25222 18680 25228 18692
rect 23676 18652 24716 18680
rect 25183 18652 25228 18680
rect 25222 18640 25228 18652
rect 25280 18640 25286 18692
rect 27798 18640 27804 18692
rect 27856 18680 27862 18692
rect 28810 18680 28816 18692
rect 27856 18652 28816 18680
rect 27856 18640 27862 18652
rect 28810 18640 28816 18652
rect 28868 18680 28874 18692
rect 28997 18683 29055 18689
rect 28997 18680 29009 18683
rect 28868 18652 29009 18680
rect 28868 18640 28874 18652
rect 28997 18649 29009 18652
rect 29043 18649 29055 18683
rect 43548 18680 43576 18711
rect 44174 18708 44180 18720
rect 44232 18708 44238 18760
rect 44361 18751 44419 18757
rect 44361 18717 44373 18751
rect 44407 18748 44419 18751
rect 44910 18748 44916 18760
rect 44407 18720 44916 18748
rect 44407 18717 44419 18720
rect 44361 18711 44419 18717
rect 44376 18680 44404 18711
rect 44910 18708 44916 18720
rect 44968 18708 44974 18760
rect 45005 18751 45063 18757
rect 45005 18717 45017 18751
rect 45051 18717 45063 18751
rect 45186 18748 45192 18760
rect 45147 18720 45192 18748
rect 45005 18711 45063 18717
rect 43548 18652 44404 18680
rect 45020 18680 45048 18711
rect 45186 18708 45192 18720
rect 45244 18708 45250 18760
rect 45094 18680 45100 18692
rect 45020 18652 45100 18680
rect 28997 18643 29055 18649
rect 45094 18640 45100 18652
rect 45152 18640 45158 18692
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18612 11207 18615
rect 11238 18612 11244 18624
rect 11195 18584 11244 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 13446 18612 13452 18624
rect 13407 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 14293 18615 14351 18621
rect 14293 18612 14305 18615
rect 13872 18584 14305 18612
rect 13872 18572 13878 18584
rect 14293 18581 14305 18584
rect 14339 18612 14351 18615
rect 14734 18612 14740 18624
rect 14339 18584 14740 18612
rect 14339 18581 14351 18584
rect 14293 18575 14351 18581
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15105 18615 15163 18621
rect 15105 18581 15117 18615
rect 15151 18612 15163 18615
rect 15470 18612 15476 18624
rect 15151 18584 15476 18612
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 26513 18615 26571 18621
rect 26513 18612 26525 18615
rect 26292 18584 26525 18612
rect 26292 18572 26298 18584
rect 26513 18581 26525 18584
rect 26559 18581 26571 18615
rect 26513 18575 26571 18581
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 19889 18411 19947 18417
rect 1995 18380 16988 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 7558 18300 7564 18352
rect 7616 18340 7622 18352
rect 12526 18340 12532 18352
rect 7616 18312 12532 18340
rect 7616 18300 7622 18312
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 12894 18340 12900 18352
rect 12855 18312 12900 18340
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 13446 18300 13452 18352
rect 13504 18300 13510 18352
rect 16025 18343 16083 18349
rect 16025 18309 16037 18343
rect 16071 18340 16083 18343
rect 16853 18343 16911 18349
rect 16853 18340 16865 18343
rect 16071 18312 16865 18340
rect 16071 18309 16083 18312
rect 16025 18303 16083 18309
rect 16853 18309 16865 18312
rect 16899 18309 16911 18343
rect 16960 18340 16988 18380
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 19978 18408 19984 18420
rect 19935 18380 19984 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 20806 18408 20812 18420
rect 20579 18380 20812 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 27890 18408 27896 18420
rect 27448 18380 27896 18408
rect 20070 18340 20076 18352
rect 16960 18312 20076 18340
rect 16853 18303 16911 18309
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 20990 18340 20996 18352
rect 20456 18312 20996 18340
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 11882 18272 11888 18284
rect 11843 18244 11888 18272
rect 11701 18235 11759 18241
rect 8570 18204 8576 18216
rect 8531 18176 8576 18204
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 8754 18204 8760 18216
rect 8715 18176 8760 18204
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18173 9091 18207
rect 11716 18204 11744 18235
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 15930 18272 15936 18284
rect 12032 18244 12077 18272
rect 15891 18244 15936 18272
rect 12032 18232 12038 18244
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16040 18244 16681 18272
rect 11790 18204 11796 18216
rect 11703 18176 11796 18204
rect 9033 18167 9091 18173
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 9048 18136 9076 18167
rect 11790 18164 11796 18176
rect 11848 18204 11854 18216
rect 12618 18204 12624 18216
rect 11848 18176 12480 18204
rect 12579 18176 12624 18204
rect 11848 18164 11854 18176
rect 4948 18108 9076 18136
rect 11701 18139 11759 18145
rect 4948 18096 4954 18108
rect 11701 18105 11713 18139
rect 11747 18136 11759 18139
rect 12342 18136 12348 18148
rect 11747 18108 12348 18136
rect 11747 18105 11759 18108
rect 11701 18099 11759 18105
rect 12342 18096 12348 18108
rect 12400 18096 12406 18148
rect 12452 18068 12480 18176
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18204 14427 18207
rect 16040 18204 16068 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 19061 18275 19119 18281
rect 19061 18272 19073 18275
rect 18104 18244 19073 18272
rect 18104 18232 18110 18244
rect 19061 18241 19073 18244
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 20456 18281 20484 18312
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 27448 18340 27476 18380
rect 27890 18368 27896 18380
rect 27948 18368 27954 18420
rect 47670 18408 47676 18420
rect 41386 18380 47164 18408
rect 47631 18380 47676 18408
rect 27614 18340 27620 18352
rect 27356 18312 27476 18340
rect 27575 18312 27620 18340
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19484 18244 19809 18272
rect 19484 18232 19490 18244
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18272 20683 18275
rect 20714 18272 20720 18284
rect 20671 18244 20720 18272
rect 20671 18241 20683 18244
rect 20625 18235 20683 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 23293 18275 23351 18281
rect 23293 18272 23305 18275
rect 21876 18244 23305 18272
rect 21876 18232 21882 18244
rect 23293 18241 23305 18244
rect 23339 18241 23351 18275
rect 25774 18272 25780 18284
rect 25735 18244 25780 18272
rect 23293 18235 23351 18241
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 27356 18281 27384 18312
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 41386 18340 41414 18380
rect 45002 18340 45008 18352
rect 31726 18312 41414 18340
rect 44652 18312 45008 18340
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18241 27399 18275
rect 27341 18235 27399 18241
rect 27430 18232 27436 18284
rect 27488 18272 27494 18284
rect 28074 18272 28080 18284
rect 27488 18244 27581 18272
rect 28035 18244 28080 18272
rect 27488 18232 27494 18244
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 14415 18176 16068 18204
rect 18509 18207 18567 18213
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 18598 18204 18604 18216
rect 18555 18176 18604 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 14384 18068 14412 18167
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18204 19211 18207
rect 20162 18204 20168 18216
rect 19199 18176 20168 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 23474 18204 23480 18216
rect 23435 18176 23480 18204
rect 23474 18164 23480 18176
rect 23532 18164 23538 18216
rect 25130 18204 25136 18216
rect 25091 18176 25136 18204
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 26326 18164 26332 18216
rect 26384 18204 26390 18216
rect 27448 18204 27476 18232
rect 28258 18204 28264 18216
rect 26384 18176 27476 18204
rect 28219 18176 28264 18204
rect 26384 18164 26390 18176
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 29914 18204 29920 18216
rect 29875 18176 29920 18204
rect 29914 18164 29920 18176
rect 29972 18164 29978 18216
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 31726 18136 31754 18312
rect 44174 18272 44180 18284
rect 44135 18244 44180 18272
rect 44174 18232 44180 18244
rect 44232 18232 44238 18284
rect 44652 18281 44680 18312
rect 45002 18300 45008 18312
rect 45060 18340 45066 18352
rect 46293 18343 46351 18349
rect 46293 18340 46305 18343
rect 45060 18312 46305 18340
rect 45060 18300 45066 18312
rect 46293 18309 46305 18312
rect 46339 18309 46351 18343
rect 46293 18303 46351 18309
rect 44637 18275 44695 18281
rect 44637 18241 44649 18275
rect 44683 18241 44695 18275
rect 44910 18272 44916 18284
rect 44871 18244 44916 18272
rect 44637 18235 44695 18241
rect 44910 18232 44916 18244
rect 44968 18232 44974 18284
rect 45922 18272 45928 18284
rect 45883 18244 45928 18272
rect 45922 18232 45928 18244
rect 45980 18232 45986 18284
rect 46109 18275 46167 18281
rect 46109 18241 46121 18275
rect 46155 18241 46167 18275
rect 46109 18235 46167 18241
rect 44450 18164 44456 18216
rect 44508 18204 44514 18216
rect 45281 18207 45339 18213
rect 45281 18204 45293 18207
rect 44508 18176 45293 18204
rect 44508 18164 44514 18176
rect 45281 18173 45293 18176
rect 45327 18204 45339 18207
rect 46124 18204 46152 18235
rect 46842 18232 46848 18284
rect 46900 18272 46906 18284
rect 47029 18275 47087 18281
rect 47029 18272 47041 18275
rect 46900 18244 47041 18272
rect 46900 18232 46906 18244
rect 47029 18241 47041 18244
rect 47075 18241 47087 18275
rect 47136 18272 47164 18380
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 47394 18272 47400 18284
rect 47136 18244 47400 18272
rect 47029 18235 47087 18241
rect 47394 18232 47400 18244
rect 47452 18272 47458 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47452 18244 47593 18272
rect 47452 18232 47458 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 45327 18176 46152 18204
rect 45327 18173 45339 18176
rect 45281 18167 45339 18173
rect 25464 18108 31754 18136
rect 25464 18096 25470 18108
rect 44818 18096 44824 18148
rect 44876 18136 44882 18148
rect 45373 18139 45431 18145
rect 45373 18136 45385 18139
rect 44876 18108 45385 18136
rect 44876 18096 44882 18108
rect 45373 18105 45385 18108
rect 45419 18105 45431 18139
rect 45373 18099 45431 18105
rect 12452 18040 14412 18068
rect 21450 18028 21456 18080
rect 21508 18068 21514 18080
rect 25590 18068 25596 18080
rect 21508 18040 25596 18068
rect 21508 18028 21514 18040
rect 25590 18028 25596 18040
rect 25648 18028 25654 18080
rect 25866 18068 25872 18080
rect 25827 18040 25872 18068
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 45094 18028 45100 18080
rect 45152 18068 45158 18080
rect 46845 18071 46903 18077
rect 46845 18068 46857 18071
rect 45152 18040 46857 18068
rect 45152 18028 45158 18040
rect 46845 18037 46857 18040
rect 46891 18037 46903 18071
rect 46845 18031 46903 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 12618 17864 12624 17876
rect 2746 17836 12434 17864
rect 12579 17836 12624 17864
rect 2130 17756 2136 17808
rect 2188 17796 2194 17808
rect 2746 17796 2774 17836
rect 2188 17768 2774 17796
rect 8297 17799 8355 17805
rect 2188 17756 2194 17768
rect 8297 17765 8309 17799
rect 8343 17796 8355 17799
rect 8754 17796 8760 17808
rect 8343 17768 8760 17796
rect 8343 17765 8355 17768
rect 8297 17759 8355 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 12406 17796 12434 17836
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 15930 17824 15936 17876
rect 15988 17864 15994 17876
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 15988 17836 16681 17864
rect 15988 17824 15994 17836
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 18230 17864 18236 17876
rect 16669 17827 16727 17833
rect 17880 17836 18236 17864
rect 17880 17796 17908 17836
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 23474 17864 23480 17876
rect 23435 17836 23480 17864
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 28077 17867 28135 17873
rect 24136 17836 26004 17864
rect 24136 17796 24164 17836
rect 8864 17768 9352 17796
rect 12406 17768 17908 17796
rect 17972 17768 24164 17796
rect 25976 17796 26004 17836
rect 28077 17833 28089 17867
rect 28123 17864 28135 17867
rect 28258 17864 28264 17876
rect 28123 17836 28264 17864
rect 28123 17833 28135 17836
rect 28077 17827 28135 17833
rect 28258 17824 28264 17836
rect 28316 17824 28322 17876
rect 44450 17864 44456 17876
rect 44411 17836 44456 17864
rect 44450 17824 44456 17836
rect 44508 17824 44514 17876
rect 44910 17824 44916 17876
rect 44968 17864 44974 17876
rect 45281 17867 45339 17873
rect 45281 17864 45293 17867
rect 44968 17836 45293 17864
rect 44968 17824 44974 17836
rect 45281 17833 45293 17836
rect 45327 17833 45339 17867
rect 45281 17827 45339 17833
rect 44634 17796 44640 17808
rect 25976 17768 44640 17796
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 8864 17728 8892 17768
rect 9030 17728 9036 17740
rect 4028 17700 8892 17728
rect 8991 17700 9036 17728
rect 4028 17688 4034 17700
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17660 8263 17663
rect 8478 17660 8484 17672
rect 8251 17632 8484 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8628 17632 9137 17660
rect 8628 17620 8634 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 2004 17496 2237 17524
rect 2004 17484 2010 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 9140 17524 9168 17623
rect 9324 17592 9352 17768
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 10229 17731 10287 17737
rect 10229 17728 10241 17731
rect 9539 17700 10241 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 10229 17697 10241 17700
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 17972 17737 18000 17768
rect 44634 17756 44640 17768
rect 44692 17796 44698 17808
rect 47394 17796 47400 17808
rect 44692 17768 47400 17796
rect 44692 17756 44698 17768
rect 47394 17756 47400 17768
rect 47452 17756 47458 17808
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 14516 17700 17969 17728
rect 14516 17688 14522 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 19996 17700 21496 17728
rect 9950 17660 9956 17672
rect 9911 17632 9956 17660
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12400 17632 12633 17660
rect 12400 17620 12406 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 14090 17660 14096 17672
rect 14003 17632 14096 17660
rect 12621 17623 12679 17629
rect 14090 17620 14096 17632
rect 14148 17660 14154 17672
rect 16577 17663 16635 17669
rect 14148 17632 16528 17660
rect 14148 17620 14154 17632
rect 10502 17592 10508 17604
rect 9324 17564 10508 17592
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 11238 17552 11244 17604
rect 11296 17552 11302 17604
rect 11701 17527 11759 17533
rect 11701 17524 11713 17527
rect 9140 17496 11713 17524
rect 2225 17487 2283 17493
rect 11701 17493 11713 17496
rect 11747 17524 11759 17527
rect 11882 17524 11888 17536
rect 11747 17496 11888 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 14274 17524 14280 17536
rect 14235 17496 14280 17524
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 16500 17524 16528 17632
rect 16577 17629 16589 17663
rect 16623 17660 16635 17663
rect 17497 17663 17555 17669
rect 17497 17660 17509 17663
rect 16623 17632 17509 17660
rect 16623 17629 16635 17632
rect 16577 17623 16635 17629
rect 17497 17629 17509 17632
rect 17543 17660 17555 17663
rect 17586 17660 17592 17672
rect 17543 17632 17592 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 17586 17620 17592 17632
rect 17644 17662 17650 17672
rect 19245 17663 19303 17669
rect 17644 17660 17724 17662
rect 17644 17634 18828 17660
rect 17644 17620 17650 17634
rect 17696 17632 18828 17634
rect 18800 17592 18828 17632
rect 19245 17629 19257 17663
rect 19291 17660 19303 17663
rect 19334 17660 19340 17672
rect 19291 17632 19340 17660
rect 19291 17629 19303 17632
rect 19245 17623 19303 17629
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 19996 17669 20024 17700
rect 21468 17672 21496 17700
rect 25866 17688 25872 17740
rect 25924 17728 25930 17740
rect 26142 17728 26148 17740
rect 25924 17700 25966 17728
rect 26103 17700 26148 17728
rect 25924 17688 25930 17700
rect 26142 17688 26148 17700
rect 26200 17688 26206 17740
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17660 20959 17663
rect 20990 17660 20996 17672
rect 20947 17632 20996 17660
rect 20947 17629 20959 17632
rect 20901 17623 20959 17629
rect 20824 17592 20852 17623
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22204 17632 22293 17660
rect 22094 17592 22100 17604
rect 18800 17564 20760 17592
rect 20824 17564 22100 17592
rect 19242 17524 19248 17536
rect 16500 17496 19248 17524
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19426 17524 19432 17536
rect 19387 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 20036 17496 20177 17524
rect 20036 17484 20042 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20732 17524 20760 17564
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 21637 17527 21695 17533
rect 21637 17524 21649 17527
rect 20732 17496 21649 17524
rect 20165 17487 20223 17493
rect 21637 17493 21649 17496
rect 21683 17524 21695 17527
rect 22204 17524 22232 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 23348 17632 23397 17660
rect 23348 17620 23354 17632
rect 23385 17629 23397 17632
rect 23431 17660 23443 17663
rect 23658 17660 23664 17672
rect 23431 17632 23664 17660
rect 23431 17629 23443 17632
rect 23385 17623 23443 17629
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 25685 17663 25743 17669
rect 25685 17629 25697 17663
rect 25731 17629 25743 17663
rect 25685 17623 25743 17629
rect 27985 17663 28043 17669
rect 27985 17629 27997 17663
rect 28031 17629 28043 17663
rect 44082 17660 44088 17672
rect 44043 17632 44088 17660
rect 27985 17623 28043 17629
rect 25700 17592 25728 17623
rect 26234 17592 26240 17604
rect 25700 17564 26240 17592
rect 26234 17552 26240 17564
rect 26292 17552 26298 17604
rect 21683 17496 22232 17524
rect 22373 17527 22431 17533
rect 21683 17493 21695 17496
rect 21637 17487 21695 17493
rect 22373 17493 22385 17527
rect 22419 17524 22431 17527
rect 23014 17524 23020 17536
rect 22419 17496 23020 17524
rect 22419 17493 22431 17496
rect 22373 17487 22431 17493
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 28000 17524 28028 17623
rect 44082 17620 44088 17632
rect 44140 17620 44146 17672
rect 44266 17660 44272 17672
rect 44227 17632 44272 17660
rect 44266 17620 44272 17632
rect 44324 17620 44330 17672
rect 45005 17663 45063 17669
rect 45005 17629 45017 17663
rect 45051 17660 45063 17663
rect 45094 17660 45100 17672
rect 45051 17632 45100 17660
rect 45051 17629 45063 17632
rect 45005 17623 45063 17629
rect 45094 17620 45100 17632
rect 45152 17620 45158 17672
rect 46290 17660 46296 17672
rect 46251 17632 46296 17660
rect 46290 17620 46296 17632
rect 46348 17620 46354 17672
rect 45186 17592 45192 17604
rect 45147 17564 45192 17592
rect 45186 17552 45192 17564
rect 45244 17552 45250 17604
rect 46477 17595 46535 17601
rect 46477 17561 46489 17595
rect 46523 17592 46535 17595
rect 47670 17592 47676 17604
rect 46523 17564 47676 17592
rect 46523 17561 46535 17564
rect 46477 17555 46535 17561
rect 47670 17552 47676 17564
rect 47728 17552 47734 17604
rect 48130 17592 48136 17604
rect 48091 17564 48136 17592
rect 48130 17552 48136 17564
rect 48188 17552 48194 17604
rect 25832 17496 28028 17524
rect 25832 17484 25838 17496
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 14 17280 20 17332
rect 72 17320 78 17332
rect 72 17292 2774 17320
rect 72 17280 78 17292
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 2746 17252 2774 17292
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10008 17292 10609 17320
rect 10008 17280 10014 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 10597 17283 10655 17289
rect 10686 17280 10692 17332
rect 10744 17320 10750 17332
rect 10744 17292 22048 17320
rect 10744 17280 10750 17292
rect 12434 17252 12440 17264
rect 2746 17224 6316 17252
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2038 17116 2044 17128
rect 1811 17088 2044 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2774 17076 2780 17128
rect 2832 17116 2838 17128
rect 2832 17088 2877 17116
rect 2832 17076 2838 17088
rect 6288 17048 6316 17224
rect 7944 17224 12440 17252
rect 7944 17193 7972 17224
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 20990 17252 20996 17264
rect 20746 17224 20996 17252
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22020 17252 22048 17292
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22646 17320 22652 17332
rect 22152 17292 22652 17320
rect 22152 17280 22158 17292
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 26142 17320 26148 17332
rect 22756 17292 26148 17320
rect 22756 17252 22784 17292
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 44361 17323 44419 17329
rect 44361 17289 44373 17323
rect 44407 17320 44419 17323
rect 45922 17320 45928 17332
rect 44407 17292 45928 17320
rect 44407 17289 44419 17292
rect 44361 17283 44419 17289
rect 45922 17280 45928 17292
rect 45980 17280 45986 17332
rect 47670 17320 47676 17332
rect 47631 17292 47676 17320
rect 47670 17280 47676 17292
rect 47728 17280 47734 17332
rect 23014 17252 23020 17264
rect 22020 17224 22784 17252
rect 22975 17224 23020 17252
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 43530 17212 43536 17264
rect 43588 17252 43594 17264
rect 44082 17252 44088 17264
rect 43588 17224 44088 17252
rect 43588 17212 43594 17224
rect 44082 17212 44088 17224
rect 44140 17252 44146 17264
rect 44140 17224 44496 17252
rect 44140 17212 44146 17224
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17184 10563 17187
rect 12342 17184 12348 17196
rect 10551 17156 12348 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 12342 17144 12348 17156
rect 12400 17184 12406 17196
rect 14185 17187 14243 17193
rect 14185 17184 14197 17187
rect 12400 17156 14197 17184
rect 12400 17144 12406 17156
rect 14185 17153 14197 17156
rect 14231 17184 14243 17187
rect 14274 17184 14280 17196
rect 14231 17156 14280 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 14274 17144 14280 17156
rect 14332 17184 14338 17196
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 14332 17156 14933 17184
rect 14332 17144 14338 17156
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15528 17156 15669 17184
rect 15528 17144 15534 17156
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 16761 17187 16819 17193
rect 16761 17153 16773 17187
rect 16807 17184 16819 17187
rect 16850 17184 16856 17196
rect 16807 17156 16856 17184
rect 16807 17153 16819 17156
rect 16761 17147 16819 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17586 17184 17592 17196
rect 17547 17156 17592 17184
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22278 17184 22284 17196
rect 22051 17156 22284 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26292 17156 26985 17184
rect 26292 17144 26298 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 44266 17184 44272 17196
rect 44179 17156 44272 17184
rect 26973 17147 27031 17153
rect 44266 17144 44272 17156
rect 44324 17144 44330 17196
rect 44468 17193 44496 17224
rect 44453 17187 44511 17193
rect 44453 17153 44465 17187
rect 44499 17153 44511 17187
rect 44453 17147 44511 17153
rect 46290 17144 46296 17196
rect 46348 17184 46354 17196
rect 47029 17187 47087 17193
rect 47029 17184 47041 17187
rect 46348 17156 47041 17184
rect 46348 17144 46354 17156
rect 47029 17153 47041 17156
rect 47075 17153 47087 17187
rect 47029 17147 47087 17153
rect 47394 17144 47400 17196
rect 47452 17184 47458 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47452 17156 47593 17184
rect 47452 17144 47458 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 8110 17116 8116 17128
rect 8071 17088 8116 17116
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 8404 17048 8432 17079
rect 9030 17076 9036 17128
rect 9088 17116 9094 17128
rect 11974 17116 11980 17128
rect 9088 17088 11980 17116
rect 9088 17076 9094 17088
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 12526 17076 12532 17128
rect 12584 17116 12590 17128
rect 17770 17116 17776 17128
rect 12584 17088 17776 17116
rect 12584 17076 12590 17088
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 19242 17116 19248 17128
rect 19203 17088 19248 17116
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17116 19579 17119
rect 20254 17116 20260 17128
rect 19567 17088 20260 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17085 21327 17119
rect 21269 17079 21327 17085
rect 22833 17119 22891 17125
rect 22833 17085 22845 17119
rect 22879 17116 22891 17119
rect 23566 17116 23572 17128
rect 22879 17088 23572 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 6288 17020 8432 17048
rect 8478 17008 8484 17060
rect 8536 17048 8542 17060
rect 15930 17048 15936 17060
rect 8536 17020 15936 17048
rect 8536 17008 8542 17020
rect 15930 17008 15936 17020
rect 15988 17008 15994 17060
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 12710 16980 12716 16992
rect 4028 16952 12716 16980
rect 4028 16940 4034 16952
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 14366 16980 14372 16992
rect 14327 16952 14372 16980
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 14921 16983 14979 16989
rect 14921 16980 14933 16983
rect 14700 16952 14933 16980
rect 14700 16940 14706 16952
rect 14921 16949 14933 16952
rect 14967 16949 14979 16983
rect 14921 16943 14979 16949
rect 15654 16940 15660 16992
rect 15712 16980 15718 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 15712 16952 15761 16980
rect 15712 16940 15718 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 15749 16943 15807 16949
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 17034 16980 17040 16992
rect 16899 16952 17040 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 21284 16980 21312 17079
rect 23566 17076 23572 17088
rect 23624 17076 23630 17128
rect 24673 17119 24731 17125
rect 24673 17085 24685 17119
rect 24719 17085 24731 17119
rect 24673 17079 24731 17085
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27246 17116 27252 17128
rect 27203 17088 27252 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 24688 17048 24716 17079
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 28813 17119 28871 17125
rect 28813 17085 28825 17119
rect 28859 17116 28871 17119
rect 28994 17116 29000 17128
rect 28859 17088 29000 17116
rect 28859 17085 28871 17088
rect 28813 17079 28871 17085
rect 28994 17076 29000 17088
rect 29052 17076 29058 17128
rect 44284 17116 44312 17144
rect 46566 17116 46572 17128
rect 44284 17088 46572 17116
rect 46566 17076 46572 17088
rect 46624 17076 46630 17128
rect 46658 17048 46664 17060
rect 24688 17020 46664 17048
rect 46658 17008 46664 17020
rect 46716 17008 46722 17060
rect 19392 16952 21312 16980
rect 21821 16983 21879 16989
rect 19392 16940 19398 16952
rect 21821 16949 21833 16983
rect 21867 16980 21879 16983
rect 22094 16980 22100 16992
rect 21867 16952 22100 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 8110 16736 8116 16788
rect 8168 16776 8174 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 8168 16748 8217 16776
rect 8168 16736 8174 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 13541 16779 13599 16785
rect 13541 16745 13553 16779
rect 13587 16776 13599 16779
rect 13630 16776 13636 16788
rect 13587 16748 13636 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 18138 16776 18144 16788
rect 17828 16748 18144 16776
rect 17828 16736 17834 16748
rect 18138 16736 18144 16748
rect 18196 16776 18202 16788
rect 18196 16748 22094 16776
rect 18196 16736 18202 16748
rect 19242 16668 19248 16720
rect 19300 16668 19306 16720
rect 22066 16708 22094 16748
rect 47486 16708 47492 16720
rect 22066 16680 47492 16708
rect 47486 16668 47492 16680
rect 47544 16668 47550 16720
rect 8202 16640 8208 16652
rect 8128 16612 8208 16640
rect 8128 16581 8156 16612
rect 8202 16600 8208 16612
rect 8260 16640 8266 16652
rect 14458 16640 14464 16652
rect 8260 16612 14464 16640
rect 8260 16600 8266 16612
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 14642 16640 14648 16652
rect 14603 16612 14648 16640
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 14918 16640 14924 16652
rect 14879 16612 14924 16640
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 16390 16640 16396 16652
rect 16303 16612 16396 16640
rect 16390 16600 16396 16612
rect 16448 16640 16454 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16448 16612 16865 16640
rect 16448 16600 16454 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 16853 16603 16911 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 19260 16640 19288 16668
rect 28994 16640 29000 16652
rect 19260 16612 29000 16640
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11974 16572 11980 16584
rect 11287 16544 11652 16572
rect 11935 16544 11980 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11330 16504 11336 16516
rect 11291 16476 11336 16504
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 11624 16504 11652 16544
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12250 16572 12256 16584
rect 12211 16544 12256 16572
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12492 16544 13001 16572
rect 12492 16532 12498 16544
rect 12989 16541 13001 16544
rect 13035 16572 13047 16575
rect 13262 16572 13268 16584
rect 13035 16544 13268 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18472 16544 19257 16572
rect 18472 16532 18478 16544
rect 19245 16541 19257 16544
rect 19291 16572 19303 16575
rect 19978 16572 19984 16584
rect 19291 16544 19984 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19978 16532 19984 16544
rect 20036 16572 20042 16584
rect 20809 16575 20867 16581
rect 20809 16572 20821 16575
rect 20036 16544 20821 16572
rect 20036 16532 20042 16544
rect 20809 16541 20821 16544
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21784 16544 21925 16572
rect 21784 16532 21790 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 22646 16572 22652 16584
rect 22559 16544 22652 16572
rect 21913 16535 21971 16541
rect 22646 16532 22652 16544
rect 22704 16572 22710 16584
rect 23382 16572 23388 16584
rect 22704 16544 23388 16572
rect 22704 16532 22710 16544
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 27338 16572 27344 16584
rect 27299 16544 27344 16572
rect 27338 16532 27344 16544
rect 27396 16532 27402 16584
rect 12342 16504 12348 16516
rect 11624 16476 12348 16504
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 13280 16476 15148 16504
rect 11790 16436 11796 16448
rect 11751 16408 11796 16436
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 13170 16436 13176 16448
rect 13131 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13280 16445 13308 16476
rect 15120 16448 15148 16476
rect 15654 16464 15660 16516
rect 15712 16464 15718 16516
rect 18690 16504 18696 16516
rect 18651 16476 18696 16504
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 20073 16507 20131 16513
rect 20073 16473 20085 16507
rect 20119 16504 20131 16507
rect 20162 16504 20168 16516
rect 20119 16476 20168 16504
rect 20119 16473 20131 16476
rect 20073 16467 20131 16473
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 21361 16507 21419 16513
rect 21361 16473 21373 16507
rect 21407 16504 21419 16507
rect 21450 16504 21456 16516
rect 21407 16476 21456 16504
rect 21407 16473 21419 16476
rect 21361 16467 21419 16473
rect 21450 16464 21456 16476
rect 21508 16464 21514 16516
rect 26050 16504 26056 16516
rect 21560 16476 26056 16504
rect 13265 16439 13323 16445
rect 13265 16405 13277 16439
rect 13311 16405 13323 16439
rect 13265 16399 13323 16405
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 13412 16408 13457 16436
rect 13412 16396 13418 16408
rect 15102 16396 15108 16448
rect 15160 16396 15166 16448
rect 20180 16436 20208 16464
rect 21560 16436 21588 16476
rect 26050 16464 26056 16476
rect 26108 16504 26114 16516
rect 40678 16504 40684 16516
rect 26108 16476 40684 16504
rect 26108 16464 26114 16476
rect 40678 16464 40684 16476
rect 40736 16464 40742 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 46750 16504 46756 16516
rect 46523 16476 46756 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 46750 16464 46756 16476
rect 46808 16464 46814 16516
rect 48130 16504 48136 16516
rect 48091 16476 48136 16504
rect 48130 16464 48136 16476
rect 48188 16464 48194 16516
rect 20180 16408 21588 16436
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 22097 16439 22155 16445
rect 22097 16436 22109 16439
rect 21876 16408 22109 16436
rect 21876 16396 21882 16408
rect 22097 16405 22109 16408
rect 22143 16405 22155 16439
rect 22738 16436 22744 16448
rect 22699 16408 22744 16436
rect 22097 16399 22155 16405
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 27525 16439 27583 16445
rect 27525 16405 27537 16439
rect 27571 16436 27583 16439
rect 27614 16436 27620 16448
rect 27571 16408 27620 16436
rect 27571 16405 27583 16408
rect 27525 16399 27583 16405
rect 27614 16396 27620 16408
rect 27672 16436 27678 16448
rect 28534 16436 28540 16448
rect 27672 16408 28540 16436
rect 27672 16396 27678 16408
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 13262 16232 13268 16244
rect 13223 16204 13268 16232
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 15470 16232 15476 16244
rect 14200 16204 15476 16232
rect 11790 16164 11796 16176
rect 11751 16136 11796 16164
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 13817 16167 13875 16173
rect 13817 16164 13829 16167
rect 13018 16136 13829 16164
rect 13817 16133 13829 16136
rect 13863 16133 13875 16167
rect 13817 16127 13875 16133
rect 11330 16056 11336 16108
rect 11388 16096 11394 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11388 16068 11529 16096
rect 11388 16056 11394 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 14200 16096 14228 16204
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 46382 16232 46388 16244
rect 18748 16204 46388 16232
rect 18748 16192 18754 16204
rect 46382 16192 46388 16204
rect 46440 16192 46446 16244
rect 46750 16232 46756 16244
rect 46711 16204 46756 16232
rect 46750 16192 46756 16204
rect 46808 16192 46814 16244
rect 15930 16164 15936 16176
rect 15870 16136 15936 16164
rect 15930 16124 15936 16136
rect 15988 16124 15994 16176
rect 17129 16167 17187 16173
rect 17129 16133 17141 16167
rect 17175 16164 17187 16167
rect 17865 16167 17923 16173
rect 17865 16164 17877 16167
rect 17175 16136 17877 16164
rect 17175 16133 17187 16136
rect 17129 16127 17187 16133
rect 17865 16133 17877 16136
rect 17911 16133 17923 16167
rect 17865 16127 17923 16133
rect 22094 16124 22100 16176
rect 22152 16164 22158 16176
rect 22152 16136 22197 16164
rect 22152 16124 22158 16136
rect 22738 16124 22744 16176
rect 22796 16124 22802 16176
rect 23382 16124 23388 16176
rect 23440 16164 23446 16176
rect 27614 16164 27620 16176
rect 23440 16136 27620 16164
rect 23440 16124 23446 16136
rect 14366 16096 14372 16108
rect 13771 16068 14228 16096
rect 14327 16068 14372 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16908 16068 17049 16096
rect 16908 16056 16914 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 17037 16059 17095 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 21818 16096 21824 16108
rect 21779 16068 21824 16096
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 24044 16105 24072 16136
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 38194 16164 38200 16176
rect 35866 16136 38200 16164
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 25409 16099 25467 16105
rect 25409 16065 25421 16099
rect 25455 16096 25467 16099
rect 35866 16096 35894 16136
rect 38194 16124 38200 16136
rect 38252 16124 38258 16176
rect 25455 16068 35894 16096
rect 25455 16065 25467 16068
rect 25409 16059 25467 16065
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 14090 16028 14096 16040
rect 13228 16000 14096 16028
rect 13228 15988 13234 16000
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 14642 16028 14648 16040
rect 14603 16000 14648 16028
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 16117 16031 16175 16037
rect 16117 16028 16129 16031
rect 15160 16000 16129 16028
rect 15160 15988 15166 16000
rect 16117 15997 16129 16000
rect 16163 16028 16175 16031
rect 17681 16031 17739 16037
rect 17681 16028 17693 16031
rect 16163 16000 17693 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 17681 15997 17693 16000
rect 17727 15997 17739 16031
rect 19518 16028 19524 16040
rect 19479 16000 19524 16028
rect 17681 15991 17739 15997
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 20346 16028 20352 16040
rect 19812 16000 20352 16028
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 19812 15892 19840 16000
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 21450 15988 21456 16040
rect 21508 16028 21514 16040
rect 25424 16028 25452 16059
rect 40678 16056 40684 16108
rect 40736 16096 40742 16108
rect 46661 16099 46719 16105
rect 46661 16096 46673 16099
rect 40736 16068 46673 16096
rect 40736 16056 40742 16068
rect 46661 16065 46673 16068
rect 46707 16065 46719 16099
rect 47762 16096 47768 16108
rect 47723 16068 47768 16096
rect 46661 16059 46719 16065
rect 47762 16056 47768 16068
rect 47820 16056 47826 16108
rect 21508 16000 25452 16028
rect 21508 15988 21514 16000
rect 3016 15864 19840 15892
rect 3016 15852 3022 15864
rect 21082 15852 21088 15904
rect 21140 15892 21146 15904
rect 22186 15892 22192 15904
rect 21140 15864 22192 15892
rect 21140 15852 21146 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23566 15892 23572 15904
rect 23527 15864 23572 15892
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 24026 15852 24032 15904
rect 24084 15892 24090 15904
rect 24121 15895 24179 15901
rect 24121 15892 24133 15895
rect 24084 15864 24133 15892
rect 24084 15852 24090 15864
rect 24121 15861 24133 15864
rect 24167 15861 24179 15895
rect 25498 15892 25504 15904
rect 25459 15864 25504 15892
rect 24121 15855 24179 15861
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 13354 15688 13360 15700
rect 13267 15660 13360 15688
rect 13354 15648 13360 15660
rect 13412 15688 13418 15700
rect 15378 15688 15384 15700
rect 13412 15660 15384 15688
rect 13412 15648 13418 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 15930 15688 15936 15700
rect 15891 15660 15936 15688
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 20254 15688 20260 15700
rect 20215 15660 20260 15688
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 46934 15688 46940 15700
rect 20404 15660 46940 15688
rect 20404 15648 20410 15660
rect 46934 15648 46940 15660
rect 46992 15648 46998 15700
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 14645 15623 14703 15629
rect 14645 15620 14657 15623
rect 12308 15592 14657 15620
rect 12308 15580 12314 15592
rect 14645 15589 14657 15592
rect 14691 15589 14703 15623
rect 14645 15583 14703 15589
rect 15105 15623 15163 15629
rect 15105 15589 15117 15623
rect 15151 15620 15163 15623
rect 15194 15620 15200 15632
rect 15151 15592 15200 15620
rect 15151 15589 15163 15592
rect 15105 15583 15163 15589
rect 15194 15580 15200 15592
rect 15252 15580 15258 15632
rect 19518 15580 19524 15632
rect 19576 15620 19582 15632
rect 19576 15592 31754 15620
rect 19576 15580 19582 15592
rect 14090 15552 14096 15564
rect 14003 15524 14096 15552
rect 14090 15512 14096 15524
rect 14148 15552 14154 15564
rect 16390 15552 16396 15564
rect 14148 15524 16396 15552
rect 14148 15512 14154 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 20714 15552 20720 15564
rect 20180 15524 20720 15552
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 2041 15447 2099 15453
rect 13188 15456 14289 15484
rect 13188 15425 13216 15456
rect 14277 15453 14289 15456
rect 14323 15484 14335 15487
rect 15102 15484 15108 15496
rect 14323 15456 15108 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 13173 15419 13231 15425
rect 13173 15385 13185 15419
rect 13219 15385 13231 15419
rect 14461 15419 14519 15425
rect 14461 15416 14473 15419
rect 13173 15379 13231 15385
rect 13464 15388 14473 15416
rect 13262 15308 13268 15360
rect 13320 15348 13326 15360
rect 13373 15351 13431 15357
rect 13373 15348 13385 15351
rect 13320 15320 13385 15348
rect 13320 15308 13326 15320
rect 13373 15317 13385 15320
rect 13419 15348 13431 15351
rect 13464 15348 13492 15388
rect 14461 15385 14473 15388
rect 14507 15416 14519 15419
rect 15396 15416 15424 15447
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15838 15484 15844 15496
rect 15528 15456 15844 15484
rect 15528 15444 15534 15456
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 20180 15493 20208 15524
rect 20714 15512 20720 15524
rect 20772 15552 20778 15564
rect 21726 15552 21732 15564
rect 20772 15524 21732 15552
rect 20772 15512 20778 15524
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 21910 15512 21916 15564
rect 21968 15552 21974 15564
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 21968 15524 22017 15552
rect 21968 15512 21974 15524
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 25498 15552 25504 15564
rect 25459 15524 25504 15552
rect 22005 15515 22063 15521
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 27154 15552 27160 15564
rect 27115 15524 27160 15552
rect 27154 15512 27160 15524
rect 27212 15512 27218 15564
rect 31726 15552 31754 15592
rect 45554 15552 45560 15564
rect 31726 15524 45560 15552
rect 45554 15512 45560 15524
rect 45612 15512 45618 15564
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 20165 15447 20223 15453
rect 14507 15388 15424 15416
rect 18233 15419 18291 15425
rect 14507 15385 14519 15388
rect 14461 15379 14519 15385
rect 18233 15385 18245 15419
rect 18279 15416 18291 15419
rect 18414 15416 18420 15428
rect 18279 15388 18420 15416
rect 18279 15385 18291 15388
rect 18233 15379 18291 15385
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 13419 15320 13492 15348
rect 13541 15351 13599 15357
rect 13419 15317 13431 15320
rect 13373 15311 13431 15317
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13998 15348 14004 15360
rect 13587 15320 14004 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 14369 15351 14427 15357
rect 14369 15317 14381 15351
rect 14415 15348 14427 15351
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 14415 15320 15301 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 15289 15317 15301 15320
rect 15335 15348 15347 15351
rect 15378 15348 15384 15360
rect 15335 15320 15384 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 18325 15351 18383 15357
rect 18325 15348 18337 15351
rect 16908 15320 18337 15348
rect 16908 15308 16914 15320
rect 18325 15317 18337 15320
rect 18371 15317 18383 15351
rect 18325 15311 18383 15317
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 20180 15348 20208 15447
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22925 15487 22983 15493
rect 22152 15456 22197 15484
rect 22152 15444 22158 15456
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 21269 15419 21327 15425
rect 21269 15385 21281 15419
rect 21315 15416 21327 15419
rect 21358 15416 21364 15428
rect 21315 15388 21364 15416
rect 21315 15385 21327 15388
rect 21269 15379 21327 15385
rect 21358 15376 21364 15388
rect 21416 15376 21422 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22940 15416 22968 15447
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 25317 15487 25375 15493
rect 25317 15484 25329 15487
rect 24452 15456 25329 15484
rect 24452 15444 24458 15456
rect 25317 15453 25329 15456
rect 25363 15453 25375 15487
rect 25317 15447 25375 15453
rect 22244 15388 22968 15416
rect 22244 15376 22250 15388
rect 19659 15320 20208 15348
rect 21453 15351 21511 15357
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 21453 15317 21465 15351
rect 21499 15348 21511 15351
rect 22002 15348 22008 15360
rect 21499 15320 22008 15348
rect 21499 15317 21511 15320
rect 21453 15311 21511 15317
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22462 15348 22468 15360
rect 22423 15320 22468 15348
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 23017 15351 23075 15357
rect 23017 15348 23029 15351
rect 22704 15320 23029 15348
rect 22704 15308 22710 15320
rect 23017 15317 23029 15320
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14700 15116 15025 15144
rect 14700 15104 14706 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15013 15107 15071 15113
rect 21726 15104 21732 15156
rect 21784 15144 21790 15156
rect 22186 15144 22192 15156
rect 21784 15116 22192 15144
rect 21784 15104 21790 15116
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 24394 15144 24400 15156
rect 24355 15116 24400 15144
rect 24394 15104 24400 15116
rect 24452 15104 24458 15156
rect 13906 15076 13912 15088
rect 13188 15048 13912 15076
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 13188 15017 13216 15048
rect 13906 15036 13912 15048
rect 13964 15036 13970 15088
rect 15194 15076 15200 15088
rect 14936 15048 15200 15076
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 14977 13231 15011
rect 13173 14971 13231 14977
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 13814 15008 13820 15020
rect 13311 14980 13820 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14090 15008 14096 15020
rect 14051 14980 14096 15008
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14936 15017 14964 15048
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 21177 15079 21235 15085
rect 21177 15045 21189 15079
rect 21223 15076 21235 15079
rect 21910 15076 21916 15088
rect 21223 15048 21916 15076
rect 21223 15045 21235 15048
rect 21177 15039 21235 15045
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 18322 15008 18328 15020
rect 18283 14980 18328 15008
rect 15105 14971 15163 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 13998 14940 14004 14952
rect 2832 14912 2877 14940
rect 13959 14912 14004 14940
rect 2832 14900 2838 14912
rect 13998 14900 14004 14912
rect 14056 14940 14062 14952
rect 15120 14940 15148 14971
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 21082 15008 21088 15020
rect 21043 14980 21088 15008
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 21358 15008 21364 15020
rect 21315 14980 21364 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 21836 15017 21864 15048
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 22462 15036 22468 15088
rect 22520 15076 22526 15088
rect 22925 15079 22983 15085
rect 22925 15076 22937 15079
rect 22520 15048 22937 15076
rect 22520 15036 22526 15048
rect 22925 15045 22937 15048
rect 22971 15045 22983 15079
rect 22925 15039 22983 15045
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 14977 21879 15011
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 21821 14971 21879 14977
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22278 15008 22284 15020
rect 22235 14980 22284 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22646 15008 22652 15020
rect 22607 14980 22652 15008
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 24026 14968 24032 15020
rect 24084 14968 24090 15020
rect 14056 14912 15148 14940
rect 18601 14943 18659 14949
rect 14056 14900 14062 14912
rect 18601 14909 18613 14943
rect 18647 14940 18659 14943
rect 18690 14940 18696 14952
rect 18647 14912 18696 14940
rect 18647 14909 18659 14912
rect 18601 14903 18659 14909
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 23566 14940 23572 14952
rect 22066 14912 23572 14940
rect 14461 14875 14519 14881
rect 14461 14841 14473 14875
rect 14507 14872 14519 14875
rect 14918 14872 14924 14884
rect 14507 14844 14924 14872
rect 14507 14841 14519 14844
rect 14461 14835 14519 14841
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 22066 14872 22094 14912
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 18380 14844 22094 14872
rect 18380 14832 18386 14844
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 13320 14776 13461 14804
rect 13320 14764 13326 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 13449 14767 13507 14773
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 22094 14804 22100 14816
rect 20956 14776 22100 14804
rect 20956 14764 20962 14776
rect 22094 14764 22100 14776
rect 22152 14804 22158 14816
rect 24394 14804 24400 14816
rect 22152 14776 24400 14804
rect 22152 14764 22158 14776
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 24946 14600 24952 14612
rect 2746 14572 24952 14600
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 2746 14396 2774 14572
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 13872 14504 17877 14532
rect 13872 14492 13878 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 21082 14532 21088 14544
rect 17865 14495 17923 14501
rect 20732 14504 21088 14532
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 17770 14464 17776 14476
rect 13964 14436 17776 14464
rect 13964 14424 13970 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 20732 14473 20760 14504
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 20956 14436 21001 14464
rect 20956 14424 20962 14436
rect 2188 14368 2774 14396
rect 2188 14356 2194 14368
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17497 14399 17555 14405
rect 17092 14368 17448 14396
rect 17092 14356 17098 14368
rect 17310 14328 17316 14340
rect 17271 14300 17316 14328
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17420 14328 17448 14368
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 18322 14396 18328 14408
rect 17543 14368 18328 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14396 20131 14399
rect 20162 14396 20168 14408
rect 20119 14368 20168 14396
rect 20119 14365 20131 14368
rect 20073 14359 20131 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 21634 14396 21640 14408
rect 21039 14368 21640 14396
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 17420 14300 17693 14328
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 20824 14328 20852 14359
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 21358 14328 21364 14340
rect 18748 14300 21364 14328
rect 18748 14288 18754 14300
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17184 14232 17601 14260
rect 17184 14220 17190 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17589 14223 17647 14229
rect 19889 14263 19947 14269
rect 19889 14229 19901 14263
rect 19935 14260 19947 14263
rect 19978 14260 19984 14272
rect 19935 14232 19984 14260
rect 19935 14229 19947 14232
rect 19889 14223 19947 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20533 14263 20591 14269
rect 20533 14260 20545 14263
rect 20128 14232 20545 14260
rect 20128 14220 20134 14232
rect 20533 14229 20545 14232
rect 20579 14229 20591 14263
rect 20533 14223 20591 14229
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 17126 14016 17132 14028
rect 17184 14056 17190 14068
rect 17184 14028 17816 14056
rect 17184 14016 17190 14028
rect 16758 13988 16764 14000
rect 16719 13960 16764 13988
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 16977 13991 17035 13997
rect 16977 13957 16989 13991
rect 17023 13988 17035 13991
rect 17678 13988 17684 14000
rect 17023 13960 17684 13988
rect 17023 13957 17035 13960
rect 16977 13951 17035 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 17788 13988 17816 14028
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18969 14059 19027 14065
rect 18969 14056 18981 14059
rect 17920 14028 18981 14056
rect 17920 14016 17926 14028
rect 18969 14025 18981 14028
rect 19015 14025 19027 14059
rect 20162 14056 20168 14068
rect 20123 14028 20168 14056
rect 18969 14019 19027 14025
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 21876 14028 22385 14056
rect 21876 14016 21882 14028
rect 22373 14025 22385 14028
rect 22419 14025 22431 14059
rect 22373 14019 22431 14025
rect 17957 13991 18015 13997
rect 17957 13988 17969 13991
rect 17788 13960 17969 13988
rect 17957 13957 17969 13960
rect 18003 13957 18015 13991
rect 18782 13988 18788 14000
rect 18743 13960 18788 13988
rect 17957 13951 18015 13957
rect 18782 13948 18788 13960
rect 18840 13988 18846 14000
rect 20898 13988 20904 14000
rect 18840 13960 20904 13988
rect 18840 13948 18846 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15804 13892 15853 13920
rect 15804 13880 15810 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 18690 13920 18696 13932
rect 17819 13892 18696 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 18690 13880 18696 13892
rect 18748 13920 18754 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18748 13892 18889 13920
rect 18748 13880 18754 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 20714 13920 20720 13932
rect 18877 13883 18935 13889
rect 19076 13892 19840 13920
rect 20675 13892 20720 13920
rect 17310 13812 17316 13864
rect 17368 13852 17374 13864
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17368 13824 17601 13852
rect 17368 13812 17374 13824
rect 17589 13821 17601 13824
rect 17635 13852 17647 13855
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17635 13824 17816 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 4798 13716 4804 13728
rect 3844 13688 4804 13716
rect 3844 13676 3850 13688
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 16025 13719 16083 13725
rect 16025 13685 16037 13719
rect 16071 13716 16083 13719
rect 16574 13716 16580 13728
rect 16071 13688 16580 13716
rect 16071 13685 16083 13688
rect 16025 13679 16083 13685
rect 16574 13676 16580 13688
rect 16632 13676 16638 13728
rect 16945 13719 17003 13725
rect 16945 13685 16957 13719
rect 16991 13716 17003 13719
rect 17218 13716 17224 13728
rect 16991 13688 17224 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 17788 13716 17816 13824
rect 17880 13824 18153 13852
rect 17880 13796 17908 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18141 13815 18199 13821
rect 18248 13824 18613 13852
rect 17862 13744 17868 13796
rect 17920 13744 17926 13796
rect 18248 13716 18276 13824
rect 18601 13821 18613 13824
rect 18647 13852 18659 13855
rect 19076 13852 19104 13892
rect 18647 13824 19104 13852
rect 19153 13855 19211 13861
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 19153 13821 19165 13855
rect 19199 13852 19211 13855
rect 19334 13852 19340 13864
rect 19199 13824 19340 13852
rect 19199 13821 19211 13824
rect 19153 13815 19211 13821
rect 19334 13812 19340 13824
rect 19392 13852 19398 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19392 13824 19717 13852
rect 19392 13812 19398 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19812 13852 19840 13892
rect 20714 13880 20720 13892
rect 20772 13920 20778 13932
rect 20990 13920 20996 13932
rect 20772 13892 20996 13920
rect 20772 13880 20778 13892
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 27338 13920 27344 13932
rect 22235 13892 27344 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 21634 13852 21640 13864
rect 19812 13824 21640 13852
rect 19705 13815 19763 13821
rect 21634 13812 21640 13824
rect 21692 13812 21698 13864
rect 20070 13784 20076 13796
rect 20031 13756 20076 13784
rect 20070 13744 20076 13756
rect 20128 13744 20134 13796
rect 17788 13688 18276 13716
rect 20714 13676 20720 13728
rect 20772 13716 20778 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20772 13688 20821 13716
rect 20772 13676 20778 13688
rect 20809 13685 20821 13688
rect 20855 13685 20867 13719
rect 20809 13679 20867 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 21634 13472 21640 13524
rect 21692 13512 21698 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21692 13484 22109 13512
rect 21692 13472 21698 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17828 13416 17908 13444
rect 17828 13404 17834 13416
rect 13262 13376 13268 13388
rect 13223 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 13587 13348 14381 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 14369 13345 14381 13348
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 14090 13308 14096 13320
rect 14051 13280 14096 13308
rect 13173 13271 13231 13277
rect 13188 13172 13216 13271
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 16390 13308 16396 13320
rect 16351 13280 16396 13308
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 17880 13308 17908 13416
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 19484 13416 19809 13444
rect 19484 13404 19490 13416
rect 19797 13413 19809 13416
rect 19843 13413 19855 13447
rect 19797 13407 19855 13413
rect 19334 13376 19340 13388
rect 19295 13348 19340 13376
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20714 13376 20720 13388
rect 20395 13348 20720 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 17880 13280 19441 13308
rect 19429 13277 19441 13280
rect 19475 13308 19487 13311
rect 19475 13280 19564 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 14826 13200 14832 13252
rect 14884 13200 14890 13252
rect 16666 13240 16672 13252
rect 16627 13212 16672 13240
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 18230 13240 18236 13252
rect 17894 13212 18236 13240
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 15378 13172 15384 13184
rect 13188 13144 15384 13172
rect 15378 13132 15384 13144
rect 15436 13172 15442 13184
rect 15841 13175 15899 13181
rect 15841 13172 15853 13175
rect 15436 13144 15853 13172
rect 15436 13132 15442 13144
rect 15841 13141 15853 13144
rect 15887 13141 15899 13175
rect 15841 13135 15899 13141
rect 17310 13132 17316 13184
rect 17368 13172 17374 13184
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 17368 13144 18153 13172
rect 17368 13132 17374 13144
rect 18141 13141 18153 13144
rect 18187 13141 18199 13175
rect 19536 13172 19564 13280
rect 19978 13200 19984 13252
rect 20036 13240 20042 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 20036 13212 20637 13240
rect 20036 13200 20042 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 21910 13240 21916 13252
rect 21850 13212 21916 13240
rect 20625 13203 20683 13209
rect 21910 13200 21916 13212
rect 21968 13200 21974 13252
rect 20898 13172 20904 13184
rect 19536 13144 20904 13172
rect 18141 13135 18199 13141
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 14090 12968 14096 12980
rect 14051 12940 14096 12968
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 14826 12968 14832 12980
rect 14783 12940 14832 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 16448 12940 16865 12968
rect 16448 12928 16454 12940
rect 16853 12937 16865 12940
rect 16899 12937 16911 12971
rect 16853 12931 16911 12937
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 17276 12940 17601 12968
rect 17276 12928 17282 12940
rect 17589 12937 17601 12940
rect 17635 12968 17647 12971
rect 17770 12968 17776 12980
rect 17635 12940 17776 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 19334 12968 19340 12980
rect 19076 12940 19340 12968
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 17310 12900 17316 12912
rect 16816 12872 17316 12900
rect 16816 12860 16822 12872
rect 17310 12860 17316 12872
rect 17368 12900 17374 12912
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 17368 12872 17417 12900
rect 17368 12860 17374 12872
rect 17405 12869 17417 12872
rect 17451 12869 17463 12903
rect 19076 12900 19104 12940
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 19518 12900 19524 12912
rect 17405 12863 17463 12869
rect 17696 12872 19104 12900
rect 19168 12872 19524 12900
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15194 12832 15200 12844
rect 14691 12804 15200 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 14108 12764 14136 12795
rect 15194 12792 15200 12804
rect 15252 12832 15258 12844
rect 15838 12832 15844 12844
rect 15252 12804 15844 12832
rect 15252 12792 15258 12804
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 17696 12841 17724 12872
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12801 17739 12835
rect 17681 12795 17739 12801
rect 18141 12835 18199 12841
rect 18141 12801 18153 12835
rect 18187 12832 18199 12835
rect 18230 12832 18236 12844
rect 18187 12804 18236 12832
rect 18187 12801 18199 12804
rect 18141 12795 18199 12801
rect 16574 12764 16580 12776
rect 14108 12736 16580 12764
rect 16574 12724 16580 12736
rect 16632 12764 16638 12776
rect 16684 12764 16712 12795
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 19168 12841 19196 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 20162 12860 20168 12912
rect 20220 12860 20226 12912
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21818 12832 21824 12844
rect 20772 12804 21824 12832
rect 20772 12792 20778 12804
rect 21818 12792 21824 12804
rect 21876 12792 21882 12844
rect 19426 12764 19432 12776
rect 16632 12736 16712 12764
rect 19387 12736 19432 12764
rect 16632 12724 16638 12736
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 30006 12696 30012 12708
rect 2746 12668 18368 12696
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 2746 12628 2774 12668
rect 1627 12600 2774 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 17000 12600 17417 12628
rect 17000 12588 17006 12600
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 18340 12628 18368 12668
rect 20456 12668 30012 12696
rect 20456 12628 20484 12668
rect 30006 12656 30012 12668
rect 30064 12656 30070 12708
rect 47762 12628 47768 12640
rect 18340 12600 20484 12628
rect 47723 12600 47768 12628
rect 17405 12591 17463 12597
rect 47762 12588 47768 12600
rect 47820 12588 47826 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 16724 12396 16957 12424
rect 16724 12384 16730 12396
rect 16945 12393 16957 12396
rect 16991 12393 17003 12427
rect 19518 12424 19524 12436
rect 19479 12396 19524 12424
rect 16945 12387 17003 12393
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 20220 12396 20269 12424
rect 20220 12384 20226 12396
rect 20257 12393 20269 12396
rect 20303 12393 20315 12427
rect 20257 12387 20315 12393
rect 20990 12288 20996 12300
rect 19444 12260 20996 12288
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15194 12220 15200 12232
rect 14783 12192 15200 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17218 12220 17224 12232
rect 17175 12192 17224 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17218 12180 17224 12192
rect 17276 12220 17282 12232
rect 17862 12220 17868 12232
rect 17276 12192 17868 12220
rect 17276 12180 17282 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 19444 12229 19472 12260
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12288 46351 12291
rect 47762 12288 47768 12300
rect 46339 12260 47768 12288
rect 46339 12257 46351 12260
rect 46293 12251 46351 12257
rect 47762 12248 47768 12260
rect 47820 12248 47826 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 20622 12220 20628 12232
rect 20211 12192 20628 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 18230 12112 18236 12164
rect 18288 12152 18294 12164
rect 20180 12152 20208 12183
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 18288 12124 20208 12152
rect 46477 12155 46535 12161
rect 18288 12112 18294 12124
rect 46477 12121 46489 12155
rect 46523 12152 46535 12155
rect 47670 12152 47676 12164
rect 46523 12124 47676 12152
rect 46523 12121 46535 12124
rect 46477 12115 46535 12121
rect 47670 12112 47676 12124
rect 47728 12112 47734 12164
rect 14829 12087 14887 12093
rect 14829 12053 14841 12087
rect 14875 12084 14887 12087
rect 15194 12084 15200 12096
rect 14875 12056 15200 12084
rect 14875 12053 14887 12056
rect 14829 12047 14887 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 47670 11880 47676 11892
rect 47631 11852 47676 11880
rect 47670 11840 47676 11852
rect 47728 11840 47734 11892
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 16761 11815 16819 11821
rect 16761 11812 16773 11815
rect 15620 11784 16773 11812
rect 15620 11772 15626 11784
rect 16761 11781 16773 11784
rect 16807 11781 16819 11815
rect 16761 11775 16819 11781
rect 16942 11772 16948 11824
rect 17000 11821 17006 11824
rect 17000 11815 17019 11821
rect 17007 11781 17019 11815
rect 17000 11775 17019 11781
rect 17000 11772 17006 11775
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 14231 11716 15853 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 15841 11713 15853 11716
rect 15887 11744 15899 11747
rect 16574 11744 16580 11756
rect 15887 11716 16580 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16574 11704 16580 11716
rect 16632 11744 16638 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 16632 11716 17601 11744
rect 16632 11704 16638 11716
rect 17589 11713 17601 11716
rect 17635 11713 17647 11747
rect 17589 11707 17647 11713
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 47581 11747 47639 11753
rect 47581 11744 47593 11747
rect 26016 11716 47593 11744
rect 26016 11704 26022 11716
rect 47581 11713 47593 11716
rect 47627 11713 47639 11747
rect 47581 11707 47639 11713
rect 17770 11608 17776 11620
rect 16960 11580 17776 11608
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13872 11512 14013 11540
rect 13872 11500 13878 11512
rect 14001 11509 14013 11512
rect 14047 11509 14059 11543
rect 16022 11540 16028 11552
rect 15983 11512 16028 11540
rect 14001 11503 14059 11509
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16960 11549 16988 11580
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 16945 11543 17003 11549
rect 16945 11509 16957 11543
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17129 11543 17187 11549
rect 17129 11540 17141 11543
rect 17092 11512 17141 11540
rect 17092 11500 17098 11512
rect 17129 11509 17141 11512
rect 17175 11509 17187 11543
rect 17678 11540 17684 11552
rect 17639 11512 17684 11540
rect 17129 11503 17187 11509
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 15654 11336 15660 11348
rect 14752 11308 15660 11336
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 14752 11141 14780 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 15488 11240 16160 11268
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13320 11104 14473 11132
rect 13320 11092 13326 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15488 11132 15516 11240
rect 16022 11200 16028 11212
rect 15983 11172 16028 11200
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 16132 11200 16160 11240
rect 16666 11200 16672 11212
rect 16132 11172 16672 11200
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 46293 11203 46351 11209
rect 46293 11169 46305 11203
rect 46339 11200 46351 11203
rect 47762 11200 47768 11212
rect 46339 11172 47768 11200
rect 46339 11169 46351 11172
rect 46293 11163 46351 11169
rect 47762 11160 47768 11172
rect 47820 11160 47826 11212
rect 15427 11104 15516 11132
rect 15565 11135 15623 11141
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 15654 11132 15660 11144
rect 15611 11104 15660 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14240 11036 14780 11064
rect 14240 11024 14246 11036
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 14148 10968 14289 10996
rect 14148 10956 14154 10968
rect 14277 10965 14289 10968
rect 14323 10965 14335 10999
rect 14752 10996 14780 11036
rect 14936 10996 14964 11095
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 18230 11132 18236 11144
rect 18191 11104 18236 11132
rect 18230 11092 18236 11104
rect 18288 11132 18294 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18288 11104 19257 11132
rect 18288 11092 18294 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 15473 11067 15531 11073
rect 15473 11033 15485 11067
rect 15519 11064 15531 11067
rect 16301 11067 16359 11073
rect 16301 11064 16313 11067
rect 15519 11036 16313 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 16301 11033 16313 11036
rect 16347 11033 16359 11067
rect 18325 11067 18383 11073
rect 18325 11064 18337 11067
rect 17526 11036 18337 11064
rect 16301 11027 16359 11033
rect 18325 11033 18337 11036
rect 18371 11033 18383 11067
rect 18325 11027 18383 11033
rect 19337 11067 19395 11073
rect 19337 11033 19349 11067
rect 19383 11064 19395 11067
rect 19426 11064 19432 11076
rect 19383 11036 19432 11064
rect 19383 11033 19395 11036
rect 19337 11027 19395 11033
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 25958 11064 25964 11076
rect 24912 11036 25964 11064
rect 24912 11024 24918 11036
rect 25958 11024 25964 11036
rect 26016 11024 26022 11076
rect 46474 11064 46480 11076
rect 46435 11036 46480 11064
rect 46474 11024 46480 11036
rect 46532 11024 46538 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 15562 10996 15568 11008
rect 14752 10968 15568 10996
rect 14277 10959 14335 10965
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 17770 10996 17776 11008
rect 17731 10968 17776 10996
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 15562 10792 15568 10804
rect 15523 10764 15568 10792
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 46474 10752 46480 10804
rect 46532 10792 46538 10804
rect 46845 10795 46903 10801
rect 46845 10792 46857 10795
rect 46532 10764 46857 10792
rect 46532 10752 46538 10764
rect 46845 10761 46857 10764
rect 46891 10761 46903 10795
rect 46845 10755 46903 10761
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 4890 10724 4896 10736
rect 2832 10696 4896 10724
rect 2832 10684 2838 10696
rect 4890 10684 4896 10696
rect 4948 10684 4954 10736
rect 14090 10724 14096 10736
rect 14051 10696 14096 10724
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 19426 10724 19432 10736
rect 19366 10696 19432 10724
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 15194 10616 15200 10668
rect 15252 10616 15258 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 17000 10628 17049 10656
rect 17000 10616 17006 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17678 10616 17684 10668
rect 17736 10656 17742 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17736 10628 17877 10656
rect 17736 10616 17742 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 46753 10659 46811 10665
rect 46753 10656 46765 10659
rect 23348 10628 46765 10656
rect 23348 10616 23354 10628
rect 46753 10625 46765 10628
rect 46799 10625 46811 10659
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 46753 10619 46811 10625
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 17218 10588 17224 10600
rect 17175 10560 17224 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17972 10560 18153 10588
rect 17405 10523 17463 10529
rect 17405 10489 17417 10523
rect 17451 10520 17463 10523
rect 17972 10520 18000 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 17451 10492 18000 10520
rect 17451 10489 17463 10492
rect 17405 10483 17463 10489
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19484 10424 19625 10452
rect 19484 10412 19490 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 46290 10452 46296 10464
rect 46251 10424 46296 10452
rect 19613 10415 19671 10421
rect 46290 10412 46296 10424
rect 46348 10412 46354 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 16724 10220 17693 10248
rect 16724 10208 16730 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17862 10180 17868 10192
rect 17000 10152 17868 10180
rect 17000 10140 17006 10152
rect 17862 10140 17868 10152
rect 17920 10140 17926 10192
rect 15378 10112 15384 10124
rect 15339 10084 15384 10112
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 17218 10072 17224 10124
rect 17276 10072 17282 10124
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 17236 10044 17264 10072
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 17236 10016 17969 10044
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 15562 9976 15568 9988
rect 15523 9948 15568 9976
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 17221 9979 17279 9985
rect 17221 9945 17233 9979
rect 17267 9976 17279 9979
rect 17586 9976 17592 9988
rect 17267 9948 17592 9976
rect 17267 9945 17279 9948
rect 17221 9939 17279 9945
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 17681 9979 17739 9985
rect 17681 9945 17693 9979
rect 17727 9976 17739 9979
rect 17770 9976 17776 9988
rect 17727 9948 17776 9976
rect 17727 9945 17739 9948
rect 17681 9939 17739 9945
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17696 9908 17724 9939
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 17862 9936 17868 9988
rect 17920 9976 17926 9988
rect 46477 9979 46535 9985
rect 17920 9948 17965 9976
rect 17920 9936 17926 9948
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 16632 9880 17724 9908
rect 16632 9868 16638 9880
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 16971 9707 17029 9713
rect 16971 9673 16983 9707
rect 17017 9704 17029 9707
rect 17218 9704 17224 9716
rect 17017 9676 17224 9704
rect 17017 9673 17029 9676
rect 16971 9667 17029 9673
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 19426 9704 19432 9716
rect 17920 9676 19432 9704
rect 17920 9664 17926 9676
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16632 9608 16773 9636
rect 16632 9596 16638 9608
rect 16761 9605 16773 9608
rect 16807 9605 16819 9639
rect 16761 9599 16819 9605
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 18693 9639 18751 9645
rect 18693 9636 18705 9639
rect 18472 9608 18705 9636
rect 18472 9596 18478 9608
rect 18693 9605 18705 9608
rect 18739 9605 18751 9639
rect 18693 9599 18751 9605
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 16908 9540 17601 9568
rect 16908 9528 16914 9540
rect 17589 9537 17601 9540
rect 17635 9568 17647 9571
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 17635 9540 18889 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 18877 9537 18889 9540
rect 18923 9568 18935 9571
rect 19242 9568 19248 9580
rect 18923 9540 19248 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19444 9577 19472 9664
rect 47670 9636 47676 9648
rect 47631 9608 47676 9636
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 46198 9568 46204 9580
rect 46159 9540 46204 9568
rect 19429 9531 19487 9537
rect 46198 9528 46204 9540
rect 46256 9528 46262 9580
rect 47486 9528 47492 9580
rect 47544 9568 47550 9580
rect 47581 9571 47639 9577
rect 47581 9568 47593 9571
rect 47544 9540 47593 9568
rect 47544 9528 47550 9540
rect 47581 9537 47593 9540
rect 47627 9537 47639 9571
rect 47581 9531 47639 9537
rect 19610 9500 19616 9512
rect 19571 9472 19616 9500
rect 19610 9460 19616 9472
rect 19668 9460 19674 9512
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 28994 9500 29000 9512
rect 21315 9472 29000 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 46474 9500 46480 9512
rect 46435 9472 46480 9500
rect 46474 9460 46480 9472
rect 46532 9460 46538 9512
rect 15654 9392 15660 9444
rect 15712 9432 15718 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 15712 9404 17141 9432
rect 15712 9392 15718 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 16942 9364 16948 9376
rect 16903 9336 16948 9364
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 17276 9336 17693 9364
rect 17276 9324 17282 9336
rect 17681 9333 17693 9336
rect 17727 9333 17739 9367
rect 17681 9327 17739 9333
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 15562 9160 15568 9172
rect 15519 9132 15568 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 19337 9163 19395 9169
rect 19337 9129 19349 9163
rect 19383 9160 19395 9163
rect 19610 9160 19616 9172
rect 19383 9132 19616 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 16758 9092 16764 9104
rect 15396 9064 16764 9092
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15396 8965 15424 9064
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 46382 9052 46388 9104
rect 46440 9092 46446 9104
rect 46440 9064 46980 9092
rect 46440 9052 46446 9064
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 18230 9024 18236 9036
rect 18191 8996 18236 9024
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 46474 9024 46480 9036
rect 46435 8996 46480 9024
rect 46474 8984 46480 8996
rect 46532 8984 46538 9036
rect 46952 9033 46980 9064
rect 46937 9027 46995 9033
rect 46937 8993 46949 9027
rect 46983 8993 46995 9027
rect 46937 8987 46995 8993
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15252 8928 15393 8956
rect 15252 8916 15258 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 19242 8956 19248 8968
rect 19203 8928 19248 8956
rect 15381 8919 15439 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 27154 8916 27160 8968
rect 27212 8956 27218 8968
rect 28350 8956 28356 8968
rect 27212 8928 28356 8956
rect 27212 8916 27218 8928
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 46290 8956 46296 8968
rect 46251 8928 46296 8956
rect 46290 8916 46296 8928
rect 46348 8916 46354 8968
rect 16758 8888 16764 8900
rect 16719 8860 16764 8888
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 17218 8548 17224 8560
rect 6886 8520 15700 8548
rect 17179 8520 17224 8548
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 6886 8344 6914 8520
rect 14182 8480 14188 8492
rect 14143 8452 14188 8480
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 14660 8344 14688 8375
rect 3384 8316 6914 8344
rect 12406 8316 14688 8344
rect 15672 8344 15700 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 47762 8548 47768 8560
rect 47723 8520 47768 8548
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 19242 8440 19248 8492
rect 19300 8480 19306 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19300 8452 19349 8480
rect 19300 8440 19306 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8412 17095 8415
rect 17402 8412 17408 8424
rect 17083 8384 17408 8412
rect 17083 8381 17095 8384
rect 17037 8375 17095 8381
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17512 8344 17540 8375
rect 15672 8316 17540 8344
rect 3384 8304 3390 8316
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 12406 8276 12434 8316
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 18012 8316 19441 8344
rect 18012 8304 18018 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 19429 8307 19487 8313
rect 30098 8304 30104 8356
rect 30156 8344 30162 8356
rect 47949 8347 48007 8353
rect 47949 8344 47961 8347
rect 30156 8316 47961 8344
rect 30156 8304 30162 8316
rect 47949 8313 47961 8316
rect 47995 8313 48007 8347
rect 47949 8307 48007 8313
rect 3200 8248 12434 8276
rect 3200 8236 3206 8248
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 45554 8276 45560 8288
rect 17644 8248 45560 8276
rect 17644 8236 17650 8248
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16758 8072 16764 8084
rect 16347 8044 16764 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 17126 8004 17132 8016
rect 16868 7976 17132 8004
rect 16868 7945 16896 7976
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17954 7936 17960 7948
rect 17083 7908 17960 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 18104 7908 18149 7936
rect 18104 7896 18110 7908
rect 46014 7896 46020 7948
rect 46072 7936 46078 7948
rect 46293 7939 46351 7945
rect 46293 7936 46305 7939
rect 46072 7908 46305 7936
rect 46072 7896 46078 7908
rect 46293 7905 46305 7908
rect 46339 7905 46351 7939
rect 48038 7936 48044 7948
rect 47999 7908 48044 7936
rect 46293 7899 46351 7905
rect 48038 7896 48044 7908
rect 48096 7896 48102 7948
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 15194 7868 15200 7880
rect 14323 7840 15200 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 16758 7868 16764 7880
rect 16255 7840 16764 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 46477 7803 46535 7809
rect 46477 7769 46489 7803
rect 46523 7800 46535 7803
rect 47486 7800 47492 7812
rect 46523 7772 47492 7800
rect 46523 7769 46535 7772
rect 46477 7763 46535 7769
rect 47486 7760 47492 7772
rect 47544 7760 47550 7812
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 18046 7528 18052 7540
rect 3660 7500 18052 7528
rect 3660 7488 3666 7500
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 1670 7420 1676 7472
rect 1728 7460 1734 7472
rect 44821 7463 44879 7469
rect 44821 7460 44833 7463
rect 1728 7432 44833 7460
rect 1728 7420 1734 7432
rect 44821 7429 44833 7432
rect 44867 7429 44879 7463
rect 44821 7423 44879 7429
rect 17218 7392 17224 7404
rect 17179 7364 17224 7392
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 17402 7324 17408 7336
rect 17363 7296 17408 7324
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 44729 7327 44787 7333
rect 44729 7293 44741 7327
rect 44775 7293 44787 7327
rect 45186 7324 45192 7336
rect 45147 7296 45192 7324
rect 44729 7287 44787 7293
rect 44744 7256 44772 7287
rect 45186 7284 45192 7296
rect 45244 7284 45250 7336
rect 47949 7259 48007 7265
rect 47949 7256 47961 7259
rect 44744 7228 47961 7256
rect 47949 7225 47961 7228
rect 47995 7225 48007 7259
rect 47949 7219 48007 7225
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17460 6956 17509 6984
rect 17460 6944 17466 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17954 6848 17960 6860
rect 3476 6820 17960 6848
rect 3476 6808 3482 6820
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 47302 6848 47308 6860
rect 47263 6820 47308 6848
rect 47302 6808 47308 6820
rect 47360 6808 47366 6860
rect 47486 6808 47492 6860
rect 47544 6848 47550 6860
rect 47581 6851 47639 6857
rect 47581 6848 47593 6851
rect 47544 6820 47593 6848
rect 47544 6808 47550 6820
rect 47581 6817 47593 6820
rect 47627 6817 47639 6851
rect 47581 6811 47639 6817
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16816 6752 17417 6780
rect 16816 6740 16822 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 48130 6304 48136 6316
rect 48091 6276 48136 6304
rect 48130 6264 48136 6276
rect 48188 6264 48194 6316
rect 47946 6100 47952 6112
rect 47907 6072 47952 6100
rect 47946 6060 47952 6072
rect 48004 6060 48010 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 46842 5720 46848 5772
rect 46900 5760 46906 5772
rect 47305 5763 47363 5769
rect 47305 5760 47317 5763
rect 46900 5732 47317 5760
rect 46900 5720 46906 5732
rect 47305 5729 47317 5732
rect 47351 5729 47363 5763
rect 47305 5723 47363 5729
rect 20809 5695 20867 5701
rect 20809 5661 20821 5695
rect 20855 5692 20867 5695
rect 21634 5692 21640 5704
rect 20855 5664 21640 5692
rect 20855 5661 20867 5664
rect 20809 5655 20867 5661
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 46566 5652 46572 5704
rect 46624 5692 46630 5704
rect 47581 5695 47639 5701
rect 47581 5692 47593 5695
rect 46624 5664 47593 5692
rect 46624 5652 46630 5664
rect 47581 5661 47593 5664
rect 47627 5661 47639 5695
rect 47581 5655 47639 5661
rect 20901 5559 20959 5565
rect 20901 5525 20913 5559
rect 20947 5556 20959 5559
rect 22186 5556 22192 5568
rect 20947 5528 22192 5556
rect 20947 5525 20959 5528
rect 20901 5519 20959 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 45830 5352 45836 5364
rect 45480 5324 45836 5352
rect 45480 5293 45508 5324
rect 45830 5312 45836 5324
rect 45888 5352 45894 5364
rect 46290 5352 46296 5364
rect 45888 5324 46296 5352
rect 45888 5312 45894 5324
rect 46290 5312 46296 5324
rect 46348 5312 46354 5364
rect 45465 5287 45523 5293
rect 45465 5253 45477 5287
rect 45511 5253 45523 5287
rect 45465 5247 45523 5253
rect 45557 5287 45615 5293
rect 45557 5253 45569 5287
rect 45603 5284 45615 5287
rect 47946 5284 47952 5296
rect 45603 5256 47952 5284
rect 45603 5253 45615 5256
rect 45557 5247 45615 5253
rect 47946 5244 47952 5256
rect 48004 5244 48010 5296
rect 18598 5216 18604 5228
rect 18559 5188 18604 5216
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 19978 5216 19984 5228
rect 19567 5188 19984 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 20346 5216 20352 5228
rect 20211 5188 20352 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 20990 5216 20996 5228
rect 20855 5188 20996 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5216 21879 5219
rect 22278 5216 22284 5228
rect 21867 5188 22284 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22480 5148 22508 5179
rect 46842 5176 46848 5228
rect 46900 5216 46906 5228
rect 47857 5219 47915 5225
rect 47857 5216 47869 5219
rect 46900 5188 47869 5216
rect 46900 5176 46906 5188
rect 47857 5185 47869 5188
rect 47903 5185 47915 5219
rect 47857 5179 47915 5185
rect 22152 5120 22508 5148
rect 45741 5151 45799 5157
rect 22152 5108 22158 5120
rect 45741 5117 45753 5151
rect 45787 5117 45799 5151
rect 45741 5111 45799 5117
rect 45186 5040 45192 5092
rect 45244 5080 45250 5092
rect 45756 5080 45784 5111
rect 45244 5052 45784 5080
rect 45244 5040 45250 5052
rect 18690 5012 18696 5024
rect 18651 4984 18696 5012
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 19610 5012 19616 5024
rect 19571 4984 19616 5012
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 5012 20315 5015
rect 20806 5012 20812 5024
rect 20303 4984 20812 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 20901 5015 20959 5021
rect 20901 4981 20913 5015
rect 20947 5012 20959 5015
rect 21542 5012 21548 5024
rect 20947 4984 21548 5012
rect 20947 4981 20959 4984
rect 20901 4975 20959 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22370 5012 22376 5024
rect 21959 4984 22376 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 23014 5012 23020 5024
rect 22603 4984 23020 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 27338 4972 27344 5024
rect 27396 5012 27402 5024
rect 48041 5015 48099 5021
rect 48041 5012 48053 5015
rect 27396 4984 48053 5012
rect 27396 4972 27402 4984
rect 48041 4981 48053 4984
rect 48087 4981 48099 5015
rect 48041 4975 48099 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 20346 4808 20352 4820
rect 20307 4780 20352 4808
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 20990 4808 20996 4820
rect 20951 4780 20996 4808
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 21634 4808 21640 4820
rect 21595 4780 21640 4808
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 22278 4808 22284 4820
rect 22239 4780 22284 4808
rect 22278 4768 22284 4780
rect 22336 4768 22342 4820
rect 46934 4740 46940 4752
rect 42720 4712 46940 4740
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 6972 4644 15301 4672
rect 6972 4632 6978 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9180 4576 9505 4604
rect 9180 4564 9186 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 9493 4567 9551 4573
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4604 19303 4607
rect 19334 4604 19340 4616
rect 19291 4576 19340 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 19668 4576 20269 4604
rect 19668 4564 19674 4576
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20864 4576 20913 4604
rect 20864 4564 20870 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 21542 4604 21548 4616
rect 21503 4576 21548 4604
rect 20901 4567 20959 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 22186 4604 22192 4616
rect 22147 4576 22192 4604
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 22830 4604 22836 4616
rect 22791 4576 22836 4604
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23477 4607 23535 4613
rect 23477 4573 23489 4607
rect 23523 4573 23535 4607
rect 39850 4604 39856 4616
rect 39811 4576 39856 4604
rect 23477 4567 23535 4573
rect 15473 4539 15531 4545
rect 15473 4505 15485 4539
rect 15519 4536 15531 4539
rect 15562 4536 15568 4548
rect 15519 4508 15568 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 17126 4536 17132 4548
rect 17087 4508 17132 4536
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 23492 4536 23520 4567
rect 39850 4564 39856 4576
rect 39908 4564 39914 4616
rect 42720 4613 42748 4712
rect 46934 4700 46940 4712
rect 46992 4700 46998 4752
rect 45830 4672 45836 4684
rect 45791 4644 45836 4672
rect 45830 4632 45836 4644
rect 45888 4632 45894 4684
rect 47026 4672 47032 4684
rect 46987 4644 47032 4672
rect 47026 4632 47032 4644
rect 47084 4632 47090 4684
rect 42705 4607 42763 4613
rect 42705 4573 42717 4607
rect 42751 4573 42763 4607
rect 42705 4567 42763 4573
rect 45186 4564 45192 4616
rect 45244 4604 45250 4616
rect 45373 4607 45431 4613
rect 45373 4604 45385 4607
rect 45244 4576 45385 4604
rect 45244 4564 45250 4576
rect 45373 4573 45385 4576
rect 45419 4573 45431 4607
rect 45373 4567 45431 4573
rect 46014 4536 46020 4548
rect 20824 4508 23520 4536
rect 45975 4508 46020 4536
rect 20824 4480 20852 4508
rect 46014 4496 46020 4508
rect 46072 4496 46078 4548
rect 18506 4468 18512 4480
rect 18467 4440 18512 4468
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 19337 4471 19395 4477
rect 19337 4437 19349 4471
rect 19383 4468 19395 4471
rect 20070 4468 20076 4480
rect 19383 4440 20076 4468
rect 19383 4437 19395 4440
rect 19337 4431 19395 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 20806 4428 20812 4480
rect 20864 4428 20870 4480
rect 22462 4428 22468 4480
rect 22520 4468 22526 4480
rect 22925 4471 22983 4477
rect 22925 4468 22937 4471
rect 22520 4440 22937 4468
rect 22520 4428 22526 4440
rect 22925 4437 22937 4440
rect 22971 4437 22983 4471
rect 23566 4468 23572 4480
rect 23527 4440 23572 4468
rect 22925 4431 22983 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 39942 4468 39948 4480
rect 39903 4440 39948 4468
rect 39942 4428 39948 4440
rect 40000 4428 40006 4480
rect 42794 4468 42800 4480
rect 42755 4440 42800 4468
rect 42794 4428 42800 4440
rect 42852 4428 42858 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 18233 4267 18291 4273
rect 18233 4233 18245 4267
rect 18279 4264 18291 4267
rect 18414 4264 18420 4276
rect 18279 4236 18420 4264
rect 18279 4233 18291 4236
rect 18233 4227 18291 4233
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 20165 4267 20223 4273
rect 20165 4264 20177 4267
rect 20036 4236 20177 4264
rect 20036 4224 20042 4236
rect 20165 4233 20177 4236
rect 20211 4233 20223 4267
rect 22830 4264 22836 4276
rect 22791 4236 22836 4264
rect 20165 4227 20223 4233
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 32950 4224 32956 4276
rect 33008 4264 33014 4276
rect 33229 4267 33287 4273
rect 33229 4264 33241 4267
rect 33008 4236 33241 4264
rect 33008 4224 33014 4236
rect 33229 4233 33241 4236
rect 33275 4233 33287 4267
rect 33229 4227 33287 4233
rect 39393 4267 39451 4273
rect 39393 4233 39405 4267
rect 39439 4264 39451 4267
rect 39850 4264 39856 4276
rect 39439 4236 39856 4264
rect 39439 4233 39451 4236
rect 39393 4227 39451 4233
rect 39850 4224 39856 4236
rect 39908 4224 39914 4276
rect 43070 4224 43076 4276
rect 43128 4264 43134 4276
rect 45830 4264 45836 4276
rect 43128 4236 45836 4264
rect 43128 4224 43134 4236
rect 45830 4224 45836 4236
rect 45888 4224 45894 4276
rect 17494 4156 17500 4208
rect 17552 4196 17558 4208
rect 21726 4196 21732 4208
rect 17552 4168 21732 4196
rect 17552 4156 17558 4168
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 21818 4156 21824 4208
rect 21876 4196 21882 4208
rect 22186 4196 22192 4208
rect 21876 4168 22192 4196
rect 21876 4156 21882 4168
rect 22186 4156 22192 4168
rect 22244 4156 22250 4208
rect 22370 4156 22376 4208
rect 22428 4196 22434 4208
rect 23661 4199 23719 4205
rect 22428 4168 22784 4196
rect 22428 4156 22434 4168
rect 8478 4128 8484 4140
rect 8439 4100 8484 4128
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 13633 4131 13691 4137
rect 11563 4100 12434 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2866 4060 2872 4072
rect 2179 4032 2872 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 1964 3992 1992 4023
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 9309 4063 9367 4069
rect 3016 4032 3061 4060
rect 3016 4020 3022 4032
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 10134 4060 10140 4072
rect 9355 4032 10140 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 3878 3992 3884 4004
rect 1964 3964 3884 3992
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 10244 3992 10272 4023
rect 9088 3964 10272 3992
rect 12406 3992 12434 4100
rect 13633 4097 13645 4131
rect 13679 4128 13691 4131
rect 17954 4128 17960 4140
rect 13679 4100 17960 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4128 18935 4131
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 18923 4100 19441 4128
rect 18923 4097 18935 4100
rect 18877 4091 18935 4097
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 20070 4128 20076 4140
rect 20031 4100 20076 4128
rect 19429 4091 19487 4097
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 18800 4060 18828 4091
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 21085 4131 21143 4137
rect 21085 4097 21097 4131
rect 21131 4128 21143 4131
rect 22462 4128 22468 4140
rect 21131 4100 22468 4128
rect 21131 4097 21143 4100
rect 21085 4091 21143 4097
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 22756 4137 22784 4168
rect 23661 4165 23673 4199
rect 23707 4196 23719 4199
rect 23842 4196 23848 4208
rect 23707 4168 23848 4196
rect 23707 4165 23719 4168
rect 23661 4159 23719 4165
rect 23842 4156 23848 4168
rect 23900 4156 23906 4208
rect 24486 4156 24492 4208
rect 24544 4196 24550 4208
rect 24581 4199 24639 4205
rect 24581 4196 24593 4199
rect 24544 4168 24593 4196
rect 24544 4156 24550 4168
rect 24581 4165 24593 4168
rect 24627 4165 24639 4199
rect 24581 4159 24639 4165
rect 25130 4156 25136 4208
rect 25188 4196 25194 4208
rect 25188 4168 25544 4196
rect 25188 4156 25194 4168
rect 22741 4131 22799 4137
rect 22741 4097 22753 4131
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 22922 4088 22928 4140
rect 22980 4128 22986 4140
rect 23382 4128 23388 4140
rect 22980 4100 23388 4128
rect 22980 4088 22986 4100
rect 23382 4088 23388 4100
rect 23440 4088 23446 4140
rect 25038 4128 25044 4140
rect 24412 4100 25044 4128
rect 17276 4032 18828 4060
rect 17276 4020 17282 4032
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19392 4032 19533 4060
rect 19392 4020 19398 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 22094 4060 22100 4072
rect 21223 4032 22100 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 23569 4063 23627 4069
rect 23569 4029 23581 4063
rect 23615 4060 23627 4063
rect 24412 4060 24440 4100
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 25406 4128 25412 4140
rect 25363 4100 25412 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 25516 4128 25544 4168
rect 32674 4156 32680 4208
rect 32732 4196 32738 4208
rect 40034 4196 40040 4208
rect 32732 4168 33272 4196
rect 32732 4156 32738 4168
rect 29178 4128 29184 4140
rect 25516 4100 29184 4128
rect 29178 4088 29184 4100
rect 29236 4088 29242 4140
rect 33134 4128 33140 4140
rect 31036 4100 31432 4128
rect 33095 4100 33140 4128
rect 23615 4032 24440 4060
rect 23615 4029 23627 4032
rect 23569 4023 23627 4029
rect 27614 4020 27620 4072
rect 27672 4060 27678 4072
rect 29086 4060 29092 4072
rect 27672 4032 29092 4060
rect 27672 4020 27678 4032
rect 29086 4020 29092 4032
rect 29144 4020 29150 4072
rect 29454 4060 29460 4072
rect 29415 4032 29460 4060
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 29641 4063 29699 4069
rect 29641 4029 29653 4063
rect 29687 4060 29699 4063
rect 30006 4060 30012 4072
rect 29687 4032 30012 4060
rect 29687 4029 29699 4032
rect 29641 4023 29699 4029
rect 30006 4020 30012 4032
rect 30064 4020 30070 4072
rect 21818 3992 21824 4004
rect 12406 3964 21824 3992
rect 9088 3952 9094 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 21928 3964 25544 3992
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8168 3896 8585 3924
rect 8168 3884 8174 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 10928 3896 11621 3924
rect 10928 3884 10934 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 13722 3924 13728 3936
rect 13683 3896 13728 3924
rect 11609 3887 11667 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 18230 3924 18236 3936
rect 14976 3896 18236 3924
rect 14976 3884 14982 3896
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19242 3924 19248 3936
rect 18840 3896 19248 3924
rect 18840 3884 18846 3896
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 21928 3924 21956 3964
rect 20496 3896 21956 3924
rect 20496 3884 20502 3896
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22281 3927 22339 3933
rect 22281 3924 22293 3927
rect 22060 3896 22293 3924
rect 22060 3884 22066 3896
rect 22281 3893 22293 3896
rect 22327 3893 22339 3927
rect 22281 3887 22339 3893
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 24820 3896 25421 3924
rect 24820 3884 24826 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25516 3924 25544 3964
rect 26970 3952 26976 4004
rect 27028 3992 27034 4004
rect 31036 3992 31064 4100
rect 31294 4060 31300 4072
rect 31255 4032 31300 4060
rect 31294 4020 31300 4032
rect 31352 4020 31358 4072
rect 27028 3964 31064 3992
rect 31404 3992 31432 4100
rect 33134 4088 33140 4100
rect 33192 4088 33198 4140
rect 33244 4128 33272 4168
rect 39132 4168 40040 4196
rect 39132 4128 39160 4168
rect 40034 4156 40040 4168
rect 40092 4156 40098 4208
rect 46658 4196 46664 4208
rect 40880 4168 41368 4196
rect 33244 4100 39160 4128
rect 39206 4088 39212 4140
rect 39264 4128 39270 4140
rect 39301 4131 39359 4137
rect 39301 4128 39313 4131
rect 39264 4100 39313 4128
rect 39264 4088 39270 4100
rect 39301 4097 39313 4100
rect 39347 4097 39359 4131
rect 39301 4091 39359 4097
rect 39574 4088 39580 4140
rect 39632 4128 39638 4140
rect 39945 4131 40003 4137
rect 39945 4128 39957 4131
rect 39632 4100 39957 4128
rect 39632 4088 39638 4100
rect 39945 4097 39957 4100
rect 39991 4097 40003 4131
rect 39945 4091 40003 4097
rect 31662 4020 31668 4072
rect 31720 4060 31726 4072
rect 40880 4060 40908 4168
rect 40954 4088 40960 4140
rect 41012 4128 41018 4140
rect 41233 4131 41291 4137
rect 41233 4128 41245 4131
rect 41012 4100 41245 4128
rect 41012 4088 41018 4100
rect 41233 4097 41245 4100
rect 41279 4097 41291 4131
rect 41340 4128 41368 4168
rect 43088 4168 44496 4196
rect 46619 4168 46664 4196
rect 43088 4128 43116 4168
rect 41340 4100 43116 4128
rect 44468 4128 44496 4168
rect 46658 4156 46664 4168
rect 46716 4156 46722 4208
rect 47762 4196 47768 4208
rect 47723 4168 47768 4196
rect 47762 4156 47768 4168
rect 47820 4156 47826 4208
rect 44468 4100 45048 4128
rect 41233 4091 41291 4097
rect 41046 4060 41052 4072
rect 31720 4032 40908 4060
rect 41007 4032 41052 4060
rect 31720 4020 31726 4032
rect 41046 4020 41052 4032
rect 41104 4060 41110 4072
rect 41322 4060 41328 4072
rect 41104 4032 41328 4060
rect 41104 4020 41110 4032
rect 41322 4020 41328 4032
rect 41380 4020 41386 4072
rect 41414 4020 41420 4072
rect 41472 4060 41478 4072
rect 43070 4060 43076 4072
rect 41472 4032 43076 4060
rect 41472 4020 41478 4032
rect 43070 4020 43076 4032
rect 43128 4020 43134 4072
rect 43257 4063 43315 4069
rect 43257 4029 43269 4063
rect 43303 4060 43315 4063
rect 43898 4060 43904 4072
rect 43303 4032 43904 4060
rect 43303 4029 43315 4032
rect 43257 4023 43315 4029
rect 43898 4020 43904 4032
rect 43956 4020 43962 4072
rect 44082 4020 44088 4072
rect 44140 4060 44146 4072
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 44140 4032 44189 4060
rect 44140 4020 44146 4032
rect 44177 4029 44189 4032
rect 44223 4029 44235 4063
rect 45020 4060 45048 4100
rect 45738 4088 45744 4140
rect 45796 4128 45802 4140
rect 45925 4131 45983 4137
rect 45925 4128 45937 4131
rect 45796 4100 45937 4128
rect 45796 4088 45802 4100
rect 45925 4097 45937 4100
rect 45971 4097 45983 4131
rect 45925 4091 45983 4097
rect 48041 4063 48099 4069
rect 48041 4060 48053 4063
rect 45020 4032 48053 4060
rect 44177 4023 44235 4029
rect 48041 4029 48053 4032
rect 48087 4029 48099 4063
rect 48041 4023 48099 4029
rect 46845 3995 46903 4001
rect 46845 3992 46857 3995
rect 31404 3964 40172 3992
rect 27028 3952 27034 3964
rect 33134 3924 33140 3936
rect 25516 3896 33140 3924
rect 25409 3887 25467 3893
rect 33134 3884 33140 3896
rect 33192 3884 33198 3936
rect 39114 3884 39120 3936
rect 39172 3924 39178 3936
rect 40037 3927 40095 3933
rect 40037 3924 40049 3927
rect 39172 3896 40049 3924
rect 39172 3884 39178 3896
rect 40037 3893 40049 3896
rect 40083 3893 40095 3927
rect 40144 3924 40172 3964
rect 41386 3964 42748 3992
rect 41386 3924 41414 3964
rect 40144 3896 41414 3924
rect 41693 3927 41751 3933
rect 40037 3887 40095 3893
rect 41693 3893 41705 3927
rect 41739 3924 41751 3927
rect 42426 3924 42432 3936
rect 41739 3896 42432 3924
rect 41739 3893 41751 3896
rect 41693 3887 41751 3893
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 42610 3924 42616 3936
rect 42571 3896 42616 3924
rect 42610 3884 42616 3896
rect 42668 3884 42674 3936
rect 42720 3924 42748 3964
rect 43272 3964 46857 3992
rect 43272 3924 43300 3964
rect 46845 3961 46857 3964
rect 46891 3961 46903 3995
rect 46845 3955 46903 3961
rect 42720 3896 43300 3924
rect 46017 3927 46075 3933
rect 46017 3893 46029 3927
rect 46063 3924 46075 3927
rect 46474 3924 46480 3936
rect 46063 3896 46480 3924
rect 46063 3893 46075 3896
rect 46017 3887 46075 3893
rect 46474 3884 46480 3896
rect 46532 3884 46538 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 2866 3720 2872 3732
rect 2827 3692 2872 3720
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3936 3692 3985 3720
rect 3936 3680 3942 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 3973 3683 4031 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 19337 3723 19395 3729
rect 19337 3720 19349 3723
rect 18196 3692 19349 3720
rect 18196 3680 18202 3692
rect 19337 3689 19349 3692
rect 19383 3689 19395 3723
rect 19337 3683 19395 3689
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 21266 3720 21272 3732
rect 19484 3692 21272 3720
rect 19484 3680 19490 3692
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 26988 3692 29040 3720
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 26988 3652 27016 3692
rect 3844 3624 27016 3652
rect 29012 3652 29040 3692
rect 29914 3680 29920 3732
rect 29972 3720 29978 3732
rect 39022 3720 39028 3732
rect 29972 3692 39028 3720
rect 29972 3680 29978 3692
rect 39022 3680 39028 3692
rect 39080 3680 39086 3732
rect 39206 3720 39212 3732
rect 39167 3692 39212 3720
rect 39206 3680 39212 3692
rect 39264 3680 39270 3732
rect 42334 3720 42340 3732
rect 39316 3692 42340 3720
rect 39316 3652 39344 3692
rect 42334 3680 42340 3692
rect 42392 3680 42398 3732
rect 43438 3680 43444 3732
rect 43496 3720 43502 3732
rect 44082 3720 44088 3732
rect 43496 3692 44088 3720
rect 43496 3680 43502 3692
rect 44082 3680 44088 3692
rect 44140 3680 44146 3732
rect 42242 3652 42248 3664
rect 29012 3624 39344 3652
rect 39408 3624 42248 3652
rect 3844 3612 3850 3624
rect 10870 3584 10876 3596
rect 2792 3556 9996 3584
rect 10831 3556 10876 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1762 3516 1768 3528
rect 1719 3488 1768 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 2130 3516 2136 3528
rect 2091 3488 2136 3516
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2792 3525 2820 3556
rect 5276 3525 5304 3556
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 5261 3479 5319 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 5399 3420 6101 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6089 3417 6101 3420
rect 6135 3417 6147 3451
rect 6089 3411 6147 3417
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 6512 3420 7757 3448
rect 6512 3408 6518 3420
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 7745 3411 7803 3417
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 9140 3448 9168 3479
rect 7984 3420 9168 3448
rect 7984 3408 7990 3420
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2004 3352 2237 3380
rect 2004 3340 2010 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 7248 3352 8309 3380
rect 7248 3340 7254 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 9968 3380 9996 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 11020 3556 11161 3584
rect 11020 3544 11026 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 18690 3584 18696 3596
rect 11149 3547 11207 3553
rect 17144 3556 18696 3584
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10686 3516 10692 3528
rect 10647 3488 10692 3516
rect 10045 3479 10103 3485
rect 10060 3448 10088 3479
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 17144 3525 17172 3556
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 21910 3584 21916 3596
rect 18800 3556 21916 3584
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13596 3488 14289 3516
rect 13596 3476 13602 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17770 3516 17776 3528
rect 17731 3488 17776 3516
rect 17129 3479 17187 3485
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18288 3488 18429 3516
rect 18288 3476 18294 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 15194 3448 15200 3460
rect 10060 3420 15200 3448
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 18800 3448 18828 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 25590 3584 25596 3596
rect 22244 3556 25596 3584
rect 22244 3544 22250 3556
rect 25590 3544 25596 3556
rect 25648 3544 25654 3596
rect 27154 3584 27160 3596
rect 27115 3556 27160 3584
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 27338 3544 27344 3596
rect 27396 3584 27402 3596
rect 27614 3584 27620 3596
rect 27396 3556 27441 3584
rect 27575 3556 27620 3584
rect 27396 3544 27402 3556
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 28994 3544 29000 3596
rect 29052 3584 29058 3596
rect 30926 3584 30932 3596
rect 29052 3556 30932 3584
rect 29052 3544 29058 3556
rect 30926 3544 30932 3556
rect 30984 3544 30990 3596
rect 31726 3556 33180 3584
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19334 3516 19340 3528
rect 19291 3488 19340 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 20070 3516 20076 3528
rect 20031 3488 20076 3516
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3485 22431 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 22373 3479 22431 3485
rect 17236 3420 18828 3448
rect 20257 3451 20315 3457
rect 17236 3380 17264 3420
rect 20257 3417 20269 3451
rect 20303 3448 20315 3451
rect 20990 3448 20996 3460
rect 20303 3420 20996 3448
rect 20303 3417 20315 3420
rect 20257 3411 20315 3417
rect 20990 3408 20996 3420
rect 21048 3408 21054 3460
rect 21082 3408 21088 3460
rect 21140 3448 21146 3460
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21140 3420 21925 3448
rect 21140 3408 21146 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 22388 3448 22416 3479
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23661 3519 23719 3525
rect 23661 3516 23673 3519
rect 23155 3488 23673 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23661 3485 23673 3488
rect 23707 3485 23719 3519
rect 23661 3479 23719 3485
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 24636 3488 25145 3516
rect 24636 3476 24642 3488
rect 25133 3485 25145 3488
rect 25179 3485 25191 3519
rect 31726 3516 31754 3556
rect 25133 3479 25191 3485
rect 28920 3488 31754 3516
rect 33152 3510 33180 3556
rect 33226 3544 33232 3596
rect 33284 3584 33290 3596
rect 39408 3584 39436 3624
rect 42242 3612 42248 3624
rect 42300 3612 42306 3664
rect 44726 3652 44732 3664
rect 42444 3624 44732 3652
rect 33284 3556 33329 3584
rect 37568 3556 39436 3584
rect 33284 3544 33290 3556
rect 35894 3516 35900 3528
rect 33244 3510 35900 3516
rect 33152 3488 35900 3510
rect 22388 3420 22600 3448
rect 21913 3411 21971 3417
rect 9968 3352 17264 3380
rect 17865 3383 17923 3389
rect 8297 3343 8355 3349
rect 17865 3349 17877 3383
rect 17911 3380 17923 3383
rect 18414 3380 18420 3392
rect 17911 3352 18420 3380
rect 17911 3349 17923 3352
rect 17865 3343 17923 3349
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 18509 3383 18567 3389
rect 18509 3349 18521 3383
rect 18555 3380 18567 3383
rect 18782 3380 18788 3392
rect 18555 3352 18788 3380
rect 18555 3349 18567 3352
rect 18509 3343 18567 3349
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 22094 3380 22100 3392
rect 20956 3352 22100 3380
rect 20956 3340 20962 3352
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 22186 3340 22192 3392
rect 22244 3380 22250 3392
rect 22465 3383 22523 3389
rect 22465 3380 22477 3383
rect 22244 3352 22477 3380
rect 22244 3340 22250 3352
rect 22465 3349 22477 3352
rect 22511 3349 22523 3383
rect 22572 3380 22600 3420
rect 22646 3408 22652 3460
rect 22704 3448 22710 3460
rect 25222 3448 25228 3460
rect 22704 3420 25228 3448
rect 22704 3408 22710 3420
rect 25222 3408 25228 3420
rect 25280 3408 25286 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 28920 3448 28948 3488
rect 33152 3482 33272 3488
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 35802 3448 35808 3460
rect 25372 3420 28948 3448
rect 29104 3420 35808 3448
rect 25372 3408 25378 3420
rect 23290 3380 23296 3392
rect 22572 3352 23296 3380
rect 22465 3343 22523 3349
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 23750 3380 23756 3392
rect 23711 3352 23756 3380
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 23842 3340 23848 3392
rect 23900 3380 23906 3392
rect 29104 3380 29132 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 36081 3451 36139 3457
rect 36081 3417 36093 3451
rect 36127 3448 36139 3451
rect 36170 3448 36176 3460
rect 36127 3420 36176 3448
rect 36127 3417 36139 3420
rect 36081 3411 36139 3417
rect 36170 3408 36176 3420
rect 36228 3408 36234 3460
rect 23900 3352 29132 3380
rect 23900 3340 23906 3352
rect 29178 3340 29184 3392
rect 29236 3380 29242 3392
rect 37568 3380 37596 3556
rect 39850 3544 39856 3596
rect 39908 3584 39914 3596
rect 39908 3556 39953 3584
rect 39908 3544 39914 3556
rect 40034 3544 40040 3596
rect 40092 3584 40098 3596
rect 40218 3584 40224 3596
rect 40092 3556 40224 3584
rect 40092 3544 40098 3556
rect 40218 3544 40224 3556
rect 40276 3584 40282 3596
rect 40313 3587 40371 3593
rect 40313 3584 40325 3587
rect 40276 3556 40325 3584
rect 40276 3544 40282 3556
rect 40313 3553 40325 3556
rect 40359 3553 40371 3587
rect 40313 3547 40371 3553
rect 40402 3544 40408 3596
rect 40460 3584 40466 3596
rect 42444 3584 42472 3624
rect 44726 3612 44732 3624
rect 44784 3652 44790 3664
rect 47026 3652 47032 3664
rect 44784 3624 47032 3652
rect 44784 3612 44790 3624
rect 47026 3612 47032 3624
rect 47084 3612 47090 3664
rect 42610 3584 42616 3596
rect 40460 3556 42472 3584
rect 42571 3556 42616 3584
rect 40460 3544 40466 3556
rect 42610 3544 42616 3556
rect 42668 3544 42674 3596
rect 42794 3584 42800 3596
rect 42755 3556 42800 3584
rect 42794 3544 42800 3556
rect 42852 3544 42858 3596
rect 43162 3584 43168 3596
rect 43123 3556 43168 3584
rect 43162 3544 43168 3556
rect 43220 3544 43226 3596
rect 45189 3587 45247 3593
rect 45189 3553 45201 3587
rect 45235 3584 45247 3587
rect 46293 3587 46351 3593
rect 46293 3584 46305 3587
rect 45235 3556 46305 3584
rect 45235 3553 45247 3556
rect 45189 3547 45247 3553
rect 46293 3553 46305 3556
rect 46339 3553 46351 3587
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46293 3547 46351 3553
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 45649 3519 45707 3525
rect 45649 3485 45661 3519
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 37737 3451 37795 3457
rect 37737 3417 37749 3451
rect 37783 3417 37795 3451
rect 37737 3411 37795 3417
rect 40037 3451 40095 3457
rect 40037 3417 40049 3451
rect 40083 3448 40095 3451
rect 40126 3448 40132 3460
rect 40083 3420 40132 3448
rect 40083 3417 40095 3420
rect 40037 3411 40095 3417
rect 29236 3352 37596 3380
rect 37752 3380 37780 3411
rect 40126 3408 40132 3420
rect 40184 3408 40190 3460
rect 41414 3408 41420 3460
rect 41472 3448 41478 3460
rect 43438 3448 43444 3460
rect 41472 3420 43444 3448
rect 41472 3408 41478 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 45664 3448 45692 3479
rect 47394 3448 47400 3460
rect 45664 3420 47400 3448
rect 47394 3408 47400 3420
rect 47452 3408 47458 3460
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 43530 3380 43536 3392
rect 37752 3352 43536 3380
rect 29236 3340 29242 3352
rect 43530 3340 43536 3352
rect 43588 3340 43594 3392
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 45741 3383 45799 3389
rect 45741 3380 45753 3383
rect 45428 3352 45753 3380
rect 45428 3340 45434 3352
rect 45741 3349 45753 3352
rect 45787 3349 45799 3383
rect 45741 3343 45799 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 17828 3148 18889 3176
rect 17828 3136 17834 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 23750 3176 23756 3188
rect 18877 3139 18935 3145
rect 19536 3148 23756 3176
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 8110 3108 8116 3120
rect 8071 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 13722 3108 13728 3120
rect 13683 3080 13728 3108
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 17184 3080 18368 3108
rect 17184 3068 17190 3080
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5960 3012 6561 3040
rect 5960 3000 5966 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 6549 3003 6607 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10744 3012 10977 3040
rect 10744 3000 10750 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 10965 3003 11023 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7800 2944 8401 2972
rect 7800 2932 7806 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 8389 2935 8447 2941
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 17773 2975 17831 2981
rect 17773 2972 17785 2975
rect 15252 2944 17785 2972
rect 15252 2932 15258 2944
rect 17773 2941 17785 2944
rect 17819 2941 17831 2975
rect 17773 2935 17831 2941
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 17678 2904 17684 2916
rect 8536 2876 17684 2904
rect 8536 2864 8542 2876
rect 17678 2864 17684 2876
rect 17736 2864 17742 2916
rect 17880 2904 17908 3003
rect 18230 2972 18236 2984
rect 18191 2944 18236 2972
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 18340 2972 18368 3080
rect 18414 3068 18420 3120
rect 18472 3108 18478 3120
rect 19150 3108 19156 3120
rect 18472 3080 19156 3108
rect 18472 3068 18478 3080
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19536 3049 19564 3148
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 25774 3176 25780 3188
rect 23860 3148 25780 3176
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20806 3108 20812 3120
rect 19659 3080 20812 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 20990 3108 20996 3120
rect 20951 3080 20996 3108
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22278 3068 22284 3120
rect 22336 3108 22342 3120
rect 23860 3108 23888 3148
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 28902 3136 28908 3188
rect 28960 3176 28966 3188
rect 32766 3176 32772 3188
rect 28960 3148 32772 3176
rect 28960 3136 28966 3148
rect 32766 3136 32772 3148
rect 32824 3136 32830 3188
rect 36170 3176 36176 3188
rect 36131 3148 36176 3176
rect 36170 3136 36176 3148
rect 36228 3136 36234 3188
rect 39574 3176 39580 3188
rect 39535 3148 39580 3176
rect 39574 3136 39580 3148
rect 39632 3136 39638 3188
rect 41414 3176 41420 3188
rect 39684 3148 41420 3176
rect 24762 3108 24768 3120
rect 22336 3080 23888 3108
rect 24723 3080 24768 3108
rect 22336 3068 22342 3080
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 24854 3068 24860 3120
rect 24912 3108 24918 3120
rect 24912 3080 32904 3108
rect 24912 3068 24918 3080
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20128 3012 20361 3040
rect 20128 3000 20134 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20898 3040 20904 3052
rect 20859 3012 20904 3040
rect 20349 3003 20407 3009
rect 20898 3000 20904 3012
rect 20956 3000 20962 3052
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 31294 3000 31300 3052
rect 31352 3040 31358 3052
rect 31352 3012 32812 3040
rect 31352 3000 31358 3012
rect 19886 2972 19892 2984
rect 18340 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 21082 2972 21088 2984
rect 20036 2944 21088 2972
rect 20036 2932 20042 2944
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 32674 2972 32680 2984
rect 29144 2944 32680 2972
rect 29144 2932 29150 2944
rect 32674 2932 32680 2944
rect 32732 2932 32738 2984
rect 21450 2904 21456 2916
rect 17880 2876 21456 2904
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 22830 2904 22836 2916
rect 21560 2876 22836 2904
rect 7282 2836 7288 2848
rect 7243 2808 7288 2836
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 21560 2836 21588 2876
rect 22830 2864 22836 2876
rect 22888 2864 22894 2916
rect 23014 2864 23020 2916
rect 23072 2904 23078 2916
rect 32122 2904 32128 2916
rect 23072 2876 32128 2904
rect 23072 2864 23078 2876
rect 32122 2864 32128 2876
rect 32180 2864 32186 2916
rect 17460 2808 21588 2836
rect 17460 2796 17466 2808
rect 23198 2796 23204 2848
rect 23256 2836 23262 2848
rect 25682 2836 25688 2848
rect 23256 2808 25688 2836
rect 23256 2796 23262 2808
rect 25682 2796 25688 2808
rect 25740 2796 25746 2848
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 32214 2836 32220 2848
rect 25832 2808 32220 2836
rect 25832 2796 25838 2808
rect 32214 2796 32220 2808
rect 32272 2796 32278 2848
rect 32784 2836 32812 3012
rect 32876 2972 32904 3080
rect 32950 3068 32956 3120
rect 33008 3108 33014 3120
rect 33229 3111 33287 3117
rect 33229 3108 33241 3111
rect 33008 3080 33241 3108
rect 33008 3068 33014 3080
rect 33229 3077 33241 3080
rect 33275 3077 33287 3111
rect 33229 3071 33287 3077
rect 33410 3068 33416 3120
rect 33468 3108 33474 3120
rect 39684 3108 39712 3148
rect 41414 3136 41420 3148
rect 41472 3136 41478 3188
rect 41509 3179 41567 3185
rect 41509 3145 41521 3179
rect 41555 3176 41567 3179
rect 43806 3176 43812 3188
rect 41555 3148 43812 3176
rect 41555 3145 41567 3148
rect 41509 3139 41567 3145
rect 43806 3136 43812 3148
rect 43864 3136 43870 3188
rect 48038 3176 48044 3188
rect 44284 3148 48044 3176
rect 41046 3108 41052 3120
rect 33468 3080 39712 3108
rect 39776 3080 41052 3108
rect 33468 3068 33474 3080
rect 33042 3040 33048 3052
rect 33003 3012 33048 3040
rect 33042 3000 33048 3012
rect 33100 3000 33106 3052
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 36136 3012 36369 3040
rect 36136 3000 36142 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 39117 3043 39175 3049
rect 39117 3009 39129 3043
rect 39163 3040 39175 3043
rect 39666 3040 39672 3052
rect 39163 3012 39672 3040
rect 39163 3009 39175 3012
rect 39117 3003 39175 3009
rect 39666 3000 39672 3012
rect 39724 3000 39730 3052
rect 33318 2972 33324 2984
rect 32876 2944 33324 2972
rect 33318 2932 33324 2944
rect 33376 2932 33382 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 35894 2932 35900 2984
rect 35952 2972 35958 2984
rect 38933 2975 38991 2981
rect 38933 2972 38945 2975
rect 35952 2944 38945 2972
rect 35952 2932 35958 2944
rect 38933 2941 38945 2944
rect 38979 2972 38991 2975
rect 39776 2972 39804 3080
rect 41046 3068 41052 3080
rect 41104 3068 41110 3120
rect 41322 3068 41328 3120
rect 41380 3108 41386 3120
rect 44284 3117 44312 3148
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 41380 3080 42625 3108
rect 41380 3068 41386 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 42613 3071 42671 3077
rect 44269 3111 44327 3117
rect 44269 3077 44281 3111
rect 44315 3077 44327 3111
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 44269 3071 44327 3077
rect 39850 3000 39856 3052
rect 39908 3040 39914 3052
rect 40126 3040 40132 3052
rect 39908 3012 40132 3040
rect 39908 3000 39914 3012
rect 40126 3000 40132 3012
rect 40184 3040 40190 3052
rect 40313 3043 40371 3049
rect 40313 3040 40325 3043
rect 40184 3012 40325 3040
rect 40184 3000 40190 3012
rect 40313 3009 40325 3012
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 40586 3000 40592 3052
rect 40644 3040 40650 3052
rect 41417 3043 41475 3049
rect 41417 3040 41429 3043
rect 40644 3012 41429 3040
rect 40644 3000 40650 3012
rect 41417 3009 41429 3012
rect 41463 3009 41475 3043
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 41417 3003 41475 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 38979 2944 39804 2972
rect 38979 2941 38991 2944
rect 38933 2935 38991 2941
rect 39942 2932 39948 2984
rect 40000 2972 40006 2984
rect 40037 2975 40095 2981
rect 40037 2972 40049 2975
rect 40000 2944 40049 2972
rect 40000 2932 40006 2944
rect 40037 2941 40049 2944
rect 40083 2941 40095 2975
rect 40037 2935 40095 2941
rect 40218 2932 40224 2984
rect 40276 2972 40282 2984
rect 44284 2972 44312 3071
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 46750 3000 46756 3052
rect 46808 3040 46814 3052
rect 47765 3043 47823 3049
rect 47765 3040 47777 3043
rect 46808 3012 47777 3040
rect 46808 3000 46814 3012
rect 47765 3009 47777 3012
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 40276 2944 44312 2972
rect 47029 2975 47087 2981
rect 40276 2932 40282 2944
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 32858 2864 32864 2916
rect 32916 2904 32922 2916
rect 47949 2907 48007 2913
rect 47949 2904 47961 2907
rect 32916 2876 47961 2904
rect 32916 2864 32922 2876
rect 47949 2873 47961 2876
rect 47995 2873 48007 2907
rect 47949 2867 48007 2873
rect 40402 2836 40408 2848
rect 32784 2808 40408 2836
rect 40402 2796 40408 2808
rect 40460 2796 40466 2848
rect 40494 2796 40500 2848
rect 40552 2836 40558 2848
rect 45094 2836 45100 2848
rect 40552 2808 45100 2836
rect 40552 2796 40558 2808
rect 45094 2796 45100 2808
rect 45152 2796 45158 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 15194 2632 15200 2644
rect 6886 2604 15200 2632
rect 6886 2564 6914 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 18598 2632 18604 2644
rect 18559 2604 18604 2632
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 19334 2632 19340 2644
rect 19295 2604 19340 2632
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 23017 2635 23075 2641
rect 20496 2604 20852 2632
rect 20496 2592 20502 2604
rect 5276 2536 6914 2564
rect 5276 2505 5304 2536
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 20533 2567 20591 2573
rect 7156 2536 7420 2564
rect 7156 2524 7162 2536
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 7282 2496 7288 2508
rect 6595 2468 7288 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7392 2505 7420 2536
rect 20533 2533 20545 2567
rect 20579 2564 20591 2567
rect 20714 2564 20720 2576
rect 20579 2536 20720 2564
rect 20579 2533 20591 2536
rect 20533 2527 20591 2533
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 20824 2564 20852 2604
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 23382 2632 23388 2644
rect 23063 2604 23388 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 25038 2592 25044 2644
rect 25096 2632 25102 2644
rect 25501 2635 25559 2641
rect 25501 2632 25513 2635
rect 25096 2604 25513 2632
rect 25096 2592 25102 2604
rect 25501 2601 25513 2604
rect 25547 2601 25559 2635
rect 26326 2632 26332 2644
rect 26287 2604 26332 2632
rect 25501 2595 25559 2601
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 45465 2635 45523 2641
rect 45465 2632 45477 2635
rect 27448 2604 45477 2632
rect 27448 2564 27476 2604
rect 45465 2601 45477 2604
rect 45511 2601 45523 2635
rect 45465 2595 45523 2601
rect 27614 2564 27620 2576
rect 20824 2536 27476 2564
rect 27575 2536 27620 2564
rect 27614 2524 27620 2536
rect 27672 2524 27678 2576
rect 32490 2524 32496 2576
rect 32548 2564 32554 2576
rect 38381 2567 38439 2573
rect 38381 2564 38393 2567
rect 32548 2536 38393 2564
rect 32548 2524 32554 2536
rect 38381 2533 38393 2536
rect 38427 2533 38439 2567
rect 38381 2527 38439 2533
rect 39298 2524 39304 2576
rect 39356 2564 39362 2576
rect 40497 2567 40555 2573
rect 40497 2564 40509 2567
rect 39356 2536 40509 2564
rect 39356 2524 39362 2536
rect 40497 2533 40509 2536
rect 40543 2533 40555 2567
rect 47949 2567 48007 2573
rect 47949 2564 47961 2567
rect 40497 2527 40555 2533
rect 45526 2536 47961 2564
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2465 7435 2499
rect 15562 2496 15568 2508
rect 15523 2468 15568 2496
rect 7377 2459 7435 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 20254 2456 20260 2508
rect 20312 2496 20318 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 20312 2468 25053 2496
rect 20312 2456 20318 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26786 2456 26792 2508
rect 26844 2496 26850 2508
rect 28721 2499 28779 2505
rect 28721 2496 28733 2499
rect 26844 2468 28733 2496
rect 26844 2456 26850 2468
rect 28721 2465 28733 2468
rect 28767 2465 28779 2499
rect 30006 2496 30012 2508
rect 29967 2468 30012 2496
rect 28721 2459 28779 2465
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 45526 2496 45554 2536
rect 47949 2533 47961 2536
rect 47995 2533 48007 2567
rect 47949 2527 48007 2533
rect 30668 2468 45554 2496
rect 46201 2499 46259 2505
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2648 2400 2697 2428
rect 2648 2388 2654 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8536 2400 8953 2428
rect 8536 2388 8542 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19208 2400 19257 2428
rect 19208 2388 19214 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21315 2400 22017 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23566 2428 23572 2440
rect 23155 2400 23572 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 25682 2428 25688 2440
rect 25643 2400 25688 2428
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 27154 2388 27160 2440
rect 27212 2428 27218 2440
rect 27212 2400 28672 2428
rect 27212 2388 27218 2400
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1360 2332 1869 2360
rect 1360 2320 1366 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7190 2360 7196 2372
rect 6779 2332 7196 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 20349 2363 20407 2369
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 20622 2360 20628 2372
rect 20395 2332 20628 2360
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21910 2360 21916 2372
rect 21131 2332 21916 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 24544 2332 24869 2360
rect 24544 2320 24550 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26237 2363 26295 2369
rect 26237 2329 26249 2363
rect 26283 2360 26295 2363
rect 26418 2360 26424 2372
rect 26283 2332 26424 2360
rect 26283 2329 26295 2332
rect 26237 2323 26295 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27120 2332 27445 2360
rect 27120 2320 27126 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28644 2360 28672 2400
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30668 2360 30696 2468
rect 46201 2465 46213 2499
rect 46247 2496 46259 2499
rect 47026 2496 47032 2508
rect 46247 2468 47032 2496
rect 46247 2465 46259 2468
rect 46201 2459 46259 2465
rect 47026 2456 47032 2468
rect 47084 2456 47090 2508
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35802 2428 35808 2440
rect 35763 2400 35808 2428
rect 35529 2391 35587 2397
rect 35802 2388 35808 2400
rect 35860 2388 35866 2440
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41230 2428 41236 2440
rect 41095 2400 41236 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 43625 2431 43683 2437
rect 41380 2400 41473 2428
rect 41380 2388 41386 2400
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 43898 2388 43904 2440
rect 43956 2428 43962 2440
rect 43956 2400 44001 2428
rect 43956 2388 43962 2400
rect 46014 2388 46020 2440
rect 46072 2428 46078 2440
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 46072 2400 46489 2428
rect 46072 2388 46078 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 46477 2391 46535 2397
rect 28644 2332 30696 2360
rect 28537 2323 28595 2329
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39356 2332 40325 2360
rect 39356 2320 39362 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40954 2320 40960 2372
rect 41012 2360 41018 2372
rect 41340 2360 41368 2388
rect 41012 2332 41368 2360
rect 45373 2363 45431 2369
rect 41012 2320 41018 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46382 2360 46388 2372
rect 45419 2332 46388 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46382 2320 46388 2332
rect 46440 2320 46446 2372
rect 47765 2363 47823 2369
rect 47765 2329 47777 2363
rect 47811 2360 47823 2363
rect 48314 2360 48320 2372
rect 47811 2332 48320 2360
rect 47811 2329 47823 2332
rect 47765 2323 47823 2329
rect 48314 2320 48320 2332
rect 48372 2320 48378 2372
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 9122 2292 9128 2304
rect 9083 2264 9128 2292
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2292 17279 2295
rect 23474 2292 23480 2304
rect 17267 2264 23480 2292
rect 17267 2261 17279 2264
rect 17221 2255 17279 2261
rect 23474 2252 23480 2264
rect 23532 2252 23538 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 9122 1980 9128 2032
rect 9180 2020 9186 2032
rect 23934 2020 23940 2032
rect 9180 1992 23940 2020
rect 9180 1980 9186 1992
rect 23934 1980 23940 1992
rect 23992 1980 23998 2032
rect 2130 1912 2136 1964
rect 2188 1952 2194 1964
rect 24670 1952 24676 1964
rect 2188 1924 24676 1952
rect 2188 1912 2194 1924
rect 24670 1912 24676 1924
rect 24728 1912 24734 1964
rect 2866 1844 2872 1896
rect 2924 1884 2930 1896
rect 21174 1884 21180 1896
rect 2924 1856 21180 1884
rect 2924 1844 2930 1856
rect 21174 1844 21180 1856
rect 21232 1844 21238 1896
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19340 47132 19392 47184
rect 29368 47132 29420 47184
rect 47860 47132 47912 47184
rect 13820 47064 13872 47116
rect 22100 47064 22152 47116
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 43168 47107 43220 47116
rect 43168 47073 43177 47107
rect 43177 47073 43211 47107
rect 43211 47073 43220 47107
rect 43168 47064 43220 47073
rect 48320 47064 48372 47116
rect 2136 47039 2188 47048
rect 2136 47005 2145 47039
rect 2145 47005 2179 47039
rect 2179 47005 2188 47039
rect 2136 46996 2188 47005
rect 2780 46996 2832 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7104 46996 7156 47048
rect 9036 46996 9088 47048
rect 11612 47039 11664 47048
rect 11612 47005 11621 47039
rect 11621 47005 11655 47039
rect 11655 47005 11664 47039
rect 11612 46996 11664 47005
rect 12256 46996 12308 47048
rect 12900 46996 12952 47048
rect 14372 47039 14424 47048
rect 14372 47005 14381 47039
rect 14381 47005 14415 47039
rect 14415 47005 14424 47039
rect 14372 46996 14424 47005
rect 16488 46996 16540 47048
rect 18696 46996 18748 47048
rect 19432 46996 19484 47048
rect 20904 47039 20956 47048
rect 20904 47005 20913 47039
rect 20913 47005 20947 47039
rect 20947 47005 20956 47039
rect 20904 46996 20956 47005
rect 2504 46971 2556 46980
rect 2504 46937 2513 46971
rect 2513 46937 2547 46971
rect 2547 46937 2556 46971
rect 2504 46928 2556 46937
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 7840 46928 7892 46980
rect 9496 46928 9548 46980
rect 11704 46928 11756 46980
rect 12440 46928 12492 46980
rect 15844 46928 15896 46980
rect 3148 46903 3200 46912
rect 3148 46869 3157 46903
rect 3157 46869 3191 46903
rect 3191 46869 3200 46903
rect 3148 46860 3200 46869
rect 6920 46903 6972 46912
rect 6920 46869 6929 46903
rect 6929 46869 6963 46903
rect 6963 46869 6972 46903
rect 6920 46860 6972 46869
rect 15292 46860 15344 46912
rect 16488 46860 16540 46912
rect 19984 46860 20036 46912
rect 24584 46996 24636 47048
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 31116 46996 31168 47048
rect 38108 46996 38160 47048
rect 41880 47039 41932 47048
rect 41880 47005 41889 47039
rect 41889 47005 41923 47039
rect 41923 47005 41932 47039
rect 41880 46996 41932 47005
rect 42616 47039 42668 47048
rect 42616 47005 42625 47039
rect 42625 47005 42659 47039
rect 42659 47005 42668 47039
rect 42616 46996 42668 47005
rect 45192 47039 45244 47048
rect 45192 47005 45201 47039
rect 45201 47005 45235 47039
rect 45235 47005 45244 47039
rect 45192 46996 45244 47005
rect 47676 46996 47728 47048
rect 21824 46903 21876 46912
rect 21824 46869 21833 46903
rect 21833 46869 21867 46903
rect 21867 46869 21876 46903
rect 21824 46860 21876 46869
rect 28264 46860 28316 46912
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 42892 46928 42944 46980
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 46388 46860 46440 46912
rect 47124 46860 47176 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 1860 46631 1912 46640
rect 1860 46597 1869 46631
rect 1869 46597 1903 46631
rect 1903 46597 1912 46631
rect 1860 46588 1912 46597
rect 3148 46588 3200 46640
rect 19432 46563 19484 46572
rect 19432 46529 19441 46563
rect 19441 46529 19475 46563
rect 19475 46529 19484 46563
rect 19432 46520 19484 46529
rect 24584 46563 24636 46572
rect 24584 46529 24593 46563
rect 24593 46529 24627 46563
rect 24627 46529 24636 46563
rect 24584 46520 24636 46529
rect 28264 46563 28316 46572
rect 28264 46529 28273 46563
rect 28273 46529 28307 46563
rect 28307 46529 28316 46563
rect 28264 46520 28316 46529
rect 3884 46452 3936 46504
rect 3976 46452 4028 46504
rect 13820 46495 13872 46504
rect 4620 46384 4672 46436
rect 11244 46384 11296 46436
rect 2596 46316 2648 46368
rect 2872 46359 2924 46368
rect 2872 46325 2881 46359
rect 2881 46325 2915 46359
rect 2915 46325 2924 46359
rect 2872 46316 2924 46325
rect 10968 46316 11020 46368
rect 13820 46461 13829 46495
rect 13829 46461 13863 46495
rect 13863 46461 13872 46495
rect 13820 46452 13872 46461
rect 14004 46495 14056 46504
rect 14004 46461 14013 46495
rect 14013 46461 14047 46495
rect 14047 46461 14056 46495
rect 14004 46452 14056 46461
rect 14188 46452 14240 46504
rect 20168 46452 20220 46504
rect 20628 46495 20680 46504
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 32220 46384 32272 46436
rect 38384 46588 38436 46640
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 45928 46588 45980 46640
rect 41880 46520 41932 46572
rect 47952 46520 48004 46572
rect 38292 46495 38344 46504
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 33784 46316 33836 46368
rect 39948 46316 40000 46368
rect 41328 46316 41380 46368
rect 42524 46384 42576 46436
rect 46296 46452 46348 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 47768 46384 47820 46436
rect 43536 46316 43588 46368
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3884 46155 3936 46164
rect 3884 46121 3893 46155
rect 3893 46121 3927 46155
rect 3927 46121 3936 46155
rect 3884 46112 3936 46121
rect 4620 46155 4672 46164
rect 4620 46121 4629 46155
rect 4629 46121 4663 46155
rect 4663 46121 4672 46155
rect 4620 46112 4672 46121
rect 11244 46155 11296 46164
rect 11244 46121 11253 46155
rect 11253 46121 11287 46155
rect 11287 46121 11296 46155
rect 11244 46112 11296 46121
rect 13820 46112 13872 46164
rect 20168 46155 20220 46164
rect 20168 46121 20177 46155
rect 20177 46121 20211 46155
rect 20211 46121 20220 46155
rect 20168 46112 20220 46121
rect 24768 46112 24820 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 20904 45976 20956 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25504 45976 25556 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 41328 46019 41380 46028
rect 41328 45985 41337 46019
rect 41337 45985 41371 46019
rect 41371 45985 41380 46019
rect 41328 45976 41380 45985
rect 41972 46019 42024 46028
rect 41972 45985 41981 46019
rect 41981 45985 42015 46019
rect 42015 45985 42024 46019
rect 41972 45976 42024 45985
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 20076 45951 20128 45960
rect 20076 45917 20085 45951
rect 20085 45917 20119 45951
rect 20119 45917 20128 45951
rect 20076 45908 20128 45917
rect 24124 45908 24176 45960
rect 38200 45951 38252 45960
rect 38200 45917 38209 45951
rect 38209 45917 38243 45951
rect 38243 45917 38252 45951
rect 38200 45908 38252 45917
rect 38384 45908 38436 45960
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 45836 45908 45888 45960
rect 2964 45815 3016 45824
rect 2964 45781 2973 45815
rect 2973 45781 3007 45815
rect 3007 45781 3016 45815
rect 2964 45772 3016 45781
rect 20720 45840 20772 45892
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 41512 45883 41564 45892
rect 41512 45849 41521 45883
rect 41521 45849 41555 45883
rect 41555 45849 41564 45883
rect 41512 45840 41564 45849
rect 46480 45883 46532 45892
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 25320 45772 25372 45824
rect 44088 45815 44140 45824
rect 44088 45781 44097 45815
rect 44097 45781 44131 45815
rect 44131 45781 44140 45815
rect 44088 45772 44140 45781
rect 45560 45772 45612 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 14004 45568 14056 45620
rect 20904 45611 20956 45620
rect 20904 45577 20913 45611
rect 20913 45577 20947 45611
rect 20947 45577 20956 45611
rect 20904 45568 20956 45577
rect 25412 45611 25464 45620
rect 25412 45577 25421 45611
rect 25421 45577 25455 45611
rect 25455 45577 25464 45611
rect 25412 45568 25464 45577
rect 32312 45568 32364 45620
rect 41512 45611 41564 45620
rect 41512 45577 41521 45611
rect 41521 45577 41555 45611
rect 41555 45577 41564 45611
rect 41512 45568 41564 45577
rect 45100 45568 45152 45620
rect 45652 45568 45704 45620
rect 2964 45500 3016 45552
rect 20720 45500 20772 45552
rect 13728 45475 13780 45484
rect 13728 45441 13737 45475
rect 13737 45441 13771 45475
rect 13771 45441 13780 45475
rect 13728 45432 13780 45441
rect 24124 45500 24176 45552
rect 42892 45543 42944 45552
rect 42892 45509 42901 45543
rect 42901 45509 42935 45543
rect 42935 45509 42944 45543
rect 42892 45500 42944 45509
rect 44180 45500 44232 45552
rect 45376 45500 45428 45552
rect 47124 45500 47176 45552
rect 25320 45475 25372 45484
rect 25320 45441 25329 45475
rect 25329 45441 25363 45475
rect 25363 45441 25372 45475
rect 25320 45432 25372 45441
rect 32128 45475 32180 45484
rect 32128 45441 32137 45475
rect 32137 45441 32171 45475
rect 32171 45441 32180 45475
rect 32128 45432 32180 45441
rect 42800 45475 42852 45484
rect 42800 45441 42809 45475
rect 42809 45441 42843 45475
rect 42843 45441 42852 45475
rect 42800 45432 42852 45441
rect 46664 45432 46716 45484
rect 2872 45364 2924 45416
rect 3056 45407 3108 45416
rect 3056 45373 3065 45407
rect 3065 45373 3099 45407
rect 3099 45373 3108 45407
rect 3056 45364 3108 45373
rect 20076 45364 20128 45416
rect 13728 45296 13780 45348
rect 37188 45296 37240 45348
rect 44456 45364 44508 45416
rect 45100 45364 45152 45416
rect 45652 45407 45704 45416
rect 45652 45373 45661 45407
rect 45661 45373 45695 45407
rect 45695 45373 45704 45407
rect 45652 45364 45704 45373
rect 46664 45296 46716 45348
rect 43996 45271 44048 45280
rect 43996 45237 44005 45271
rect 44005 45237 44039 45271
rect 44039 45237 44048 45271
rect 43996 45228 44048 45237
rect 47216 45228 47268 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 42616 45024 42668 45076
rect 44456 45067 44508 45076
rect 44456 45033 44465 45067
rect 44465 45033 44499 45067
rect 44499 45033 44508 45067
rect 44456 45024 44508 45033
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 46480 45024 46532 45076
rect 42800 44956 42852 45008
rect 47400 44956 47452 45008
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 44916 44820 44968 44872
rect 45652 44863 45704 44872
rect 45652 44829 45661 44863
rect 45661 44829 45695 44863
rect 45695 44829 45704 44863
rect 45652 44820 45704 44829
rect 46940 44752 46992 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 46296 44523 46348 44532
rect 46296 44489 46305 44523
rect 46305 44489 46339 44523
rect 46339 44489 46348 44523
rect 46296 44480 46348 44489
rect 46940 44523 46992 44532
rect 46940 44489 46949 44523
rect 46949 44489 46983 44523
rect 46983 44489 46992 44523
rect 46940 44480 46992 44489
rect 45652 44412 45704 44464
rect 45192 44344 45244 44396
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 37188 44276 37240 44328
rect 25320 44140 25372 44192
rect 25872 44140 25924 44192
rect 47676 44183 47728 44192
rect 47676 44149 47685 44183
rect 47685 44149 47719 44183
rect 47719 44149 47728 44183
rect 47676 44140 47728 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 47676 43800 47728 43852
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1860 43299 1912 43308
rect 1860 43265 1869 43299
rect 1869 43265 1903 43299
rect 1903 43265 1912 43299
rect 1860 43256 1912 43265
rect 25504 43256 25556 43308
rect 32128 43256 32180 43308
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 47768 43299 47820 43308
rect 47768 43265 47777 43299
rect 47777 43265 47811 43299
rect 47811 43265 47820 43299
rect 47768 43256 47820 43265
rect 1952 43095 2004 43104
rect 1952 43061 1961 43095
rect 1961 43061 1995 43095
rect 1995 43061 2004 43095
rect 1952 43052 2004 43061
rect 25964 43095 26016 43104
rect 25964 43061 25973 43095
rect 25973 43061 26007 43095
rect 26007 43061 26016 43095
rect 25964 43052 26016 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 25964 42755 26016 42764
rect 25964 42721 25973 42755
rect 25973 42721 26007 42755
rect 26007 42721 26016 42755
rect 25964 42712 26016 42721
rect 33784 42712 33836 42764
rect 25228 42644 25280 42696
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 25228 42347 25280 42356
rect 25228 42313 25237 42347
rect 25237 42313 25271 42347
rect 25271 42313 25280 42347
rect 25228 42304 25280 42313
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 25320 42168 25372 42220
rect 46296 42168 46348 42220
rect 47400 42168 47452 42220
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47676 41624 47728 41676
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 46480 41216 46532 41268
rect 2136 41123 2188 41132
rect 2136 41089 2145 41123
rect 2145 41089 2179 41123
rect 2179 41089 2188 41123
rect 2136 41080 2188 41089
rect 45836 41080 45888 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 43720 40876 43772 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 47676 40715 47728 40724
rect 47676 40681 47685 40715
rect 47685 40681 47719 40715
rect 47719 40681 47728 40715
rect 47676 40672 47728 40681
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 2412 40400 2464 40452
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 46296 39788 46348 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 46940 39312 46992 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 46940 39083 46992 39092
rect 46940 39049 46949 39083
rect 46949 39049 46983 39083
rect 46983 39049 46992 39083
rect 46940 39040 46992 39049
rect 46112 38904 46164 38956
rect 47768 38947 47820 38956
rect 47768 38913 47777 38947
rect 47777 38913 47811 38947
rect 47811 38913 47820 38947
rect 47768 38904 47820 38913
rect 47768 38700 47820 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 47676 38224 47728 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 47676 37995 47728 38004
rect 47676 37961 47685 37995
rect 47685 37961 47719 37995
rect 47719 37961 47728 37995
rect 47676 37952 47728 37961
rect 25136 37884 25188 37936
rect 19432 37816 19484 37868
rect 32128 37816 32180 37868
rect 19524 37612 19576 37664
rect 25044 37748 25096 37800
rect 26240 37680 26292 37732
rect 26148 37655 26200 37664
rect 26148 37621 26157 37655
rect 26157 37621 26191 37655
rect 26191 37621 26200 37655
rect 26148 37612 26200 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 25044 37451 25096 37460
rect 25044 37417 25053 37451
rect 25053 37417 25087 37451
rect 25087 37417 25096 37451
rect 25044 37408 25096 37417
rect 46296 37408 46348 37460
rect 19524 37315 19576 37324
rect 19524 37281 19533 37315
rect 19533 37281 19567 37315
rect 19567 37281 19576 37315
rect 19524 37272 19576 37281
rect 27252 37315 27304 37324
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 27252 37281 27261 37315
rect 27261 37281 27295 37315
rect 27295 37281 27304 37315
rect 27252 37272 27304 37281
rect 21180 37136 21232 37188
rect 20260 37068 20312 37120
rect 22468 37068 22520 37120
rect 23664 37111 23716 37120
rect 23664 37077 23673 37111
rect 23673 37077 23707 37111
rect 23707 37077 23716 37111
rect 23664 37068 23716 37077
rect 45560 37272 45612 37324
rect 27068 37111 27120 37120
rect 27068 37077 27077 37111
rect 27077 37077 27111 37111
rect 27111 37077 27120 37111
rect 27068 37068 27120 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 21180 36907 21232 36916
rect 21180 36873 21189 36907
rect 21189 36873 21223 36907
rect 21223 36873 21232 36907
rect 21180 36864 21232 36873
rect 21824 36796 21876 36848
rect 20168 36728 20220 36780
rect 21088 36771 21140 36780
rect 21088 36737 21097 36771
rect 21097 36737 21131 36771
rect 21131 36737 21140 36771
rect 21088 36728 21140 36737
rect 20444 36660 20496 36712
rect 27252 36864 27304 36916
rect 23664 36796 23716 36848
rect 25228 36728 25280 36780
rect 26148 36728 26200 36780
rect 22560 36660 22612 36712
rect 22928 36703 22980 36712
rect 22928 36669 22937 36703
rect 22937 36669 22971 36703
rect 22971 36669 22980 36703
rect 22928 36660 22980 36669
rect 24860 36660 24912 36712
rect 27068 36660 27120 36712
rect 20168 36524 20220 36576
rect 24952 36524 25004 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19432 36320 19484 36372
rect 22928 36320 22980 36372
rect 25136 36320 25188 36372
rect 12440 36252 12492 36304
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 20168 36227 20220 36236
rect 20168 36193 20177 36227
rect 20177 36193 20211 36227
rect 20211 36193 20220 36227
rect 20168 36184 20220 36193
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 20260 36116 20312 36168
rect 22468 36184 22520 36236
rect 22836 36116 22888 36168
rect 23204 36159 23256 36168
rect 2228 36048 2280 36100
rect 23204 36125 23213 36159
rect 23213 36125 23247 36159
rect 23247 36125 23256 36159
rect 23204 36116 23256 36125
rect 24400 35980 24452 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 19984 35708 20036 35760
rect 23204 35708 23256 35760
rect 1400 35640 1452 35692
rect 21088 35640 21140 35692
rect 22468 35683 22520 35692
rect 22468 35649 22477 35683
rect 22477 35649 22511 35683
rect 22511 35649 22520 35683
rect 22468 35640 22520 35649
rect 15844 35572 15896 35624
rect 22744 35572 22796 35624
rect 9496 35504 9548 35556
rect 26976 35640 27028 35692
rect 29644 35640 29696 35692
rect 26240 35572 26292 35624
rect 27528 35572 27580 35624
rect 29000 35572 29052 35624
rect 7840 35436 7892 35488
rect 18144 35436 18196 35488
rect 22468 35436 22520 35488
rect 27160 35436 27212 35488
rect 28632 35436 28684 35488
rect 30012 35479 30064 35488
rect 30012 35445 30021 35479
rect 30021 35445 30055 35479
rect 30055 35445 30064 35479
rect 30012 35436 30064 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 20260 35232 20312 35284
rect 24952 35275 25004 35284
rect 24952 35241 24961 35275
rect 24961 35241 24995 35275
rect 24995 35241 25004 35275
rect 24952 35232 25004 35241
rect 26976 35232 27028 35284
rect 29644 35275 29696 35284
rect 19064 35164 19116 35216
rect 19248 35096 19300 35148
rect 21456 35096 21508 35148
rect 22560 35096 22612 35148
rect 23020 35096 23072 35148
rect 26148 35139 26200 35148
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 2320 35028 2372 35080
rect 14740 35071 14792 35080
rect 14740 35037 14749 35071
rect 14749 35037 14783 35071
rect 14783 35037 14792 35071
rect 14740 35028 14792 35037
rect 20628 35028 20680 35080
rect 21088 35028 21140 35080
rect 25228 35071 25280 35080
rect 25228 35037 25237 35071
rect 25237 35037 25271 35071
rect 25271 35037 25280 35071
rect 25228 35028 25280 35037
rect 26148 35105 26157 35139
rect 26157 35105 26191 35139
rect 26191 35105 26200 35139
rect 26148 35096 26200 35105
rect 27620 35096 27672 35148
rect 29644 35241 29653 35275
rect 29653 35241 29687 35275
rect 29687 35241 29696 35275
rect 29644 35232 29696 35241
rect 15016 35003 15068 35012
rect 15016 34969 15025 35003
rect 15025 34969 15059 35003
rect 15059 34969 15068 35003
rect 15016 34960 15068 34969
rect 16396 34960 16448 35012
rect 1492 34892 1544 34944
rect 17132 34892 17184 34944
rect 17684 34960 17736 35012
rect 20168 34960 20220 35012
rect 21824 35003 21876 35012
rect 21824 34969 21833 35003
rect 21833 34969 21867 35003
rect 21867 34969 21876 35003
rect 21824 34960 21876 34969
rect 22468 34960 22520 35012
rect 24952 35003 25004 35012
rect 24952 34969 24961 35003
rect 24961 34969 24995 35003
rect 24995 34969 25004 35003
rect 24952 34960 25004 34969
rect 25964 34960 26016 35012
rect 31760 35028 31812 35080
rect 47308 35071 47360 35080
rect 47308 35037 47317 35071
rect 47317 35037 47351 35071
rect 47351 35037 47360 35071
rect 47308 35028 47360 35037
rect 47492 35028 47544 35080
rect 27160 34960 27212 35012
rect 20352 34892 20404 34944
rect 20996 34935 21048 34944
rect 20996 34901 21005 34935
rect 21005 34901 21039 34935
rect 21039 34901 21048 34935
rect 20996 34892 21048 34901
rect 23296 34935 23348 34944
rect 23296 34901 23305 34935
rect 23305 34901 23339 34935
rect 23339 34901 23348 34935
rect 23296 34892 23348 34901
rect 25412 34935 25464 34944
rect 25412 34901 25421 34935
rect 25421 34901 25455 34935
rect 25455 34901 25464 34935
rect 25412 34892 25464 34901
rect 26148 34892 26200 34944
rect 31208 34935 31260 34944
rect 31208 34901 31217 34935
rect 31217 34901 31251 34935
rect 31251 34901 31260 34935
rect 31208 34892 31260 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 17684 34688 17736 34740
rect 15016 34620 15068 34672
rect 15844 34595 15896 34604
rect 15844 34561 15853 34595
rect 15853 34561 15887 34595
rect 15887 34561 15896 34595
rect 15844 34552 15896 34561
rect 16120 34552 16172 34604
rect 18052 34620 18104 34672
rect 18972 34595 19024 34604
rect 17132 34484 17184 34536
rect 18144 34527 18196 34536
rect 18144 34493 18153 34527
rect 18153 34493 18187 34527
rect 18187 34493 18196 34527
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 19984 34620 20036 34672
rect 20260 34620 20312 34672
rect 21824 34688 21876 34740
rect 23112 34688 23164 34740
rect 26056 34688 26108 34740
rect 28816 34688 28868 34740
rect 29000 34731 29052 34740
rect 29000 34697 29009 34731
rect 29009 34697 29043 34731
rect 29043 34697 29052 34731
rect 29000 34688 29052 34697
rect 18144 34484 18196 34493
rect 17960 34416 18012 34468
rect 16120 34348 16172 34400
rect 19064 34484 19116 34536
rect 19524 34595 19576 34604
rect 19524 34561 19533 34595
rect 19533 34561 19567 34595
rect 19567 34561 19576 34595
rect 19524 34552 19576 34561
rect 20168 34552 20220 34604
rect 20444 34552 20496 34604
rect 21824 34595 21876 34604
rect 21824 34561 21833 34595
rect 21833 34561 21867 34595
rect 21867 34561 21876 34595
rect 21824 34552 21876 34561
rect 24768 34620 24820 34672
rect 27528 34620 27580 34672
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 22928 34552 22980 34604
rect 23020 34552 23072 34604
rect 26976 34595 27028 34604
rect 26976 34561 26985 34595
rect 26985 34561 27019 34595
rect 27019 34561 27028 34595
rect 26976 34552 27028 34561
rect 28448 34595 28500 34604
rect 23296 34484 23348 34536
rect 24492 34527 24544 34536
rect 24492 34493 24501 34527
rect 24501 34493 24535 34527
rect 24535 34493 24544 34527
rect 24492 34484 24544 34493
rect 28448 34561 28457 34595
rect 28457 34561 28491 34595
rect 28491 34561 28500 34595
rect 28448 34552 28500 34561
rect 28632 34595 28684 34604
rect 28632 34561 28641 34595
rect 28641 34561 28675 34595
rect 28675 34561 28684 34595
rect 28632 34552 28684 34561
rect 28816 34595 28868 34604
rect 28816 34561 28825 34595
rect 28825 34561 28859 34595
rect 28859 34561 28868 34595
rect 28816 34552 28868 34561
rect 31208 34552 31260 34604
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 20444 34416 20496 34468
rect 25964 34459 26016 34468
rect 25964 34425 25973 34459
rect 25973 34425 26007 34459
rect 26007 34425 26016 34459
rect 25964 34416 26016 34425
rect 29736 34484 29788 34536
rect 30104 34527 30156 34536
rect 30104 34493 30113 34527
rect 30113 34493 30147 34527
rect 30147 34493 30156 34527
rect 30104 34484 30156 34493
rect 29000 34416 29052 34468
rect 19524 34348 19576 34400
rect 20168 34391 20220 34400
rect 20168 34357 20177 34391
rect 20177 34357 20211 34391
rect 20211 34357 20220 34391
rect 20168 34348 20220 34357
rect 29736 34348 29788 34400
rect 30196 34348 30248 34400
rect 47952 34391 48004 34400
rect 47952 34357 47961 34391
rect 47961 34357 47995 34391
rect 47995 34357 48004 34391
rect 47952 34348 48004 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 16396 34187 16448 34196
rect 16396 34153 16405 34187
rect 16405 34153 16439 34187
rect 16439 34153 16448 34187
rect 16396 34144 16448 34153
rect 24492 34144 24544 34196
rect 29000 34187 29052 34196
rect 24768 34076 24820 34128
rect 28448 34076 28500 34128
rect 28540 34076 28592 34128
rect 29000 34153 29009 34187
rect 29009 34153 29043 34187
rect 29043 34153 29052 34187
rect 29000 34144 29052 34153
rect 29736 34144 29788 34196
rect 30104 34144 30156 34196
rect 30656 34144 30708 34196
rect 29644 34076 29696 34128
rect 19340 34008 19392 34060
rect 21456 34008 21508 34060
rect 24952 34051 25004 34060
rect 24952 34017 24961 34051
rect 24961 34017 24995 34051
rect 24995 34017 25004 34051
rect 24952 34008 25004 34017
rect 25228 34008 25280 34060
rect 16120 33940 16172 33992
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 25412 33940 25464 33992
rect 27712 33940 27764 33992
rect 28448 33983 28500 33992
rect 28448 33949 28457 33983
rect 28457 33949 28491 33983
rect 28491 33949 28500 33983
rect 28448 33940 28500 33949
rect 20720 33872 20772 33924
rect 20996 33872 21048 33924
rect 23388 33872 23440 33924
rect 20628 33804 20680 33856
rect 21916 33847 21968 33856
rect 21916 33813 21925 33847
rect 21925 33813 21959 33847
rect 21959 33813 21968 33847
rect 21916 33804 21968 33813
rect 23756 33804 23808 33856
rect 24768 33872 24820 33924
rect 27896 33872 27948 33924
rect 29184 34008 29236 34060
rect 31024 34008 31076 34060
rect 47952 34008 48004 34060
rect 29460 33940 29512 33992
rect 29736 33981 29788 33992
rect 29736 33947 29745 33981
rect 29745 33947 29779 33981
rect 29779 33947 29788 33981
rect 29736 33940 29788 33947
rect 30104 33983 30156 33992
rect 30104 33949 30113 33983
rect 30113 33949 30147 33983
rect 30147 33949 30156 33983
rect 30932 33983 30984 33992
rect 30104 33940 30156 33949
rect 30932 33949 30941 33983
rect 30941 33949 30975 33983
rect 30975 33949 30984 33983
rect 30932 33940 30984 33949
rect 31760 33983 31812 33992
rect 31760 33949 31769 33983
rect 31769 33949 31803 33983
rect 31803 33949 31812 33983
rect 31760 33940 31812 33949
rect 29276 33872 29328 33924
rect 26976 33804 27028 33856
rect 30564 33804 30616 33856
rect 30748 33915 30800 33924
rect 30748 33881 30757 33915
rect 30757 33881 30791 33915
rect 30791 33881 30800 33915
rect 30748 33872 30800 33881
rect 47492 33872 47544 33924
rect 31668 33804 31720 33856
rect 31944 33804 31996 33856
rect 45836 33804 45888 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 18052 33643 18104 33652
rect 18052 33609 18061 33643
rect 18061 33609 18095 33643
rect 18095 33609 18104 33643
rect 18052 33600 18104 33609
rect 18972 33600 19024 33652
rect 20536 33643 20588 33652
rect 20536 33609 20545 33643
rect 20545 33609 20579 33643
rect 20579 33609 20588 33643
rect 20536 33600 20588 33609
rect 21824 33600 21876 33652
rect 23756 33643 23808 33652
rect 19524 33464 19576 33516
rect 20260 33464 20312 33516
rect 20628 33464 20680 33516
rect 20812 33464 20864 33516
rect 21824 33507 21876 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 2044 33396 2096 33448
rect 17776 33439 17828 33448
rect 17776 33405 17785 33439
rect 17785 33405 17819 33439
rect 17819 33405 17828 33439
rect 17776 33396 17828 33405
rect 19294 33388 19346 33440
rect 21824 33473 21833 33507
rect 21833 33473 21867 33507
rect 21867 33473 21876 33507
rect 21824 33464 21876 33473
rect 22192 33507 22244 33516
rect 22192 33473 22201 33507
rect 22201 33473 22235 33507
rect 22235 33473 22244 33507
rect 22192 33464 22244 33473
rect 23296 33532 23348 33584
rect 23756 33609 23765 33643
rect 23765 33609 23799 33643
rect 23799 33609 23808 33643
rect 23756 33600 23808 33609
rect 23940 33643 23992 33652
rect 23940 33609 23949 33643
rect 23949 33609 23983 33643
rect 23983 33609 23992 33643
rect 23940 33600 23992 33609
rect 23848 33507 23900 33516
rect 23848 33473 23890 33507
rect 23890 33473 23900 33507
rect 23848 33464 23900 33473
rect 23204 33396 23256 33448
rect 24768 33532 24820 33584
rect 25044 33600 25096 33652
rect 29460 33600 29512 33652
rect 28816 33532 28868 33584
rect 17684 33303 17736 33312
rect 17684 33269 17693 33303
rect 17693 33269 17727 33303
rect 17727 33269 17736 33303
rect 17684 33260 17736 33269
rect 20168 33260 20220 33312
rect 23020 33328 23072 33380
rect 23112 33260 23164 33312
rect 23388 33260 23440 33312
rect 25228 33464 25280 33516
rect 25780 33507 25832 33516
rect 25780 33473 25789 33507
rect 25789 33473 25823 33507
rect 25823 33473 25832 33507
rect 25780 33464 25832 33473
rect 26148 33464 26200 33516
rect 26976 33507 27028 33516
rect 26976 33473 26985 33507
rect 26985 33473 27019 33507
rect 27019 33473 27028 33507
rect 26976 33464 27028 33473
rect 27896 33507 27948 33516
rect 27896 33473 27905 33507
rect 27905 33473 27939 33507
rect 27939 33473 27948 33507
rect 27896 33464 27948 33473
rect 28080 33507 28132 33516
rect 28080 33473 28089 33507
rect 28089 33473 28123 33507
rect 28123 33473 28132 33507
rect 28080 33464 28132 33473
rect 28448 33464 28500 33516
rect 27712 33396 27764 33448
rect 29276 33507 29328 33516
rect 29276 33473 29285 33507
rect 29285 33473 29319 33507
rect 29319 33473 29328 33507
rect 29736 33507 29788 33516
rect 29276 33464 29328 33473
rect 29736 33473 29745 33507
rect 29745 33473 29779 33507
rect 29779 33473 29788 33507
rect 29736 33464 29788 33473
rect 30104 33532 30156 33584
rect 30196 33464 30248 33516
rect 30656 33507 30708 33516
rect 30656 33473 30665 33507
rect 30665 33473 30699 33507
rect 30699 33473 30708 33507
rect 30656 33464 30708 33473
rect 30932 33532 30984 33584
rect 47860 33507 47912 33516
rect 47860 33473 47869 33507
rect 47869 33473 47903 33507
rect 47903 33473 47912 33507
rect 47860 33464 47912 33473
rect 30472 33396 30524 33448
rect 28448 33328 28500 33380
rect 29460 33328 29512 33380
rect 30380 33328 30432 33380
rect 25136 33303 25188 33312
rect 25136 33269 25145 33303
rect 25145 33269 25179 33303
rect 25179 33269 25188 33303
rect 25136 33260 25188 33269
rect 25596 33260 25648 33312
rect 25872 33260 25924 33312
rect 27896 33260 27948 33312
rect 29552 33260 29604 33312
rect 30012 33303 30064 33312
rect 30012 33269 30021 33303
rect 30021 33269 30055 33303
rect 30055 33269 30064 33303
rect 30012 33260 30064 33269
rect 30288 33260 30340 33312
rect 30472 33260 30524 33312
rect 30932 33260 30984 33312
rect 44180 33260 44232 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17684 33056 17736 33108
rect 21456 33056 21508 33108
rect 24400 33099 24452 33108
rect 1492 32988 1544 33040
rect 15936 32988 15988 33040
rect 20628 33031 20680 33040
rect 16672 32895 16724 32904
rect 16672 32861 16681 32895
rect 16681 32861 16715 32895
rect 16715 32861 16724 32895
rect 16672 32852 16724 32861
rect 16948 32895 17000 32904
rect 16948 32861 16957 32895
rect 16957 32861 16991 32895
rect 16991 32861 17000 32895
rect 16948 32852 17000 32861
rect 17960 32920 18012 32972
rect 18236 32920 18288 32972
rect 20628 32997 20637 33031
rect 20637 32997 20671 33031
rect 20671 32997 20680 33031
rect 20628 32988 20680 32997
rect 24400 33065 24409 33099
rect 24409 33065 24443 33099
rect 24443 33065 24452 33099
rect 24400 33056 24452 33065
rect 24860 33099 24912 33108
rect 24860 33065 24869 33099
rect 24869 33065 24903 33099
rect 24903 33065 24912 33099
rect 24860 33056 24912 33065
rect 25780 33056 25832 33108
rect 25136 32988 25188 33040
rect 19524 32963 19576 32972
rect 1400 32784 1452 32836
rect 3240 32827 3292 32836
rect 3240 32793 3249 32827
rect 3249 32793 3283 32827
rect 3283 32793 3292 32827
rect 3240 32784 3292 32793
rect 16856 32827 16908 32836
rect 16856 32793 16865 32827
rect 16865 32793 16899 32827
rect 16899 32793 16908 32827
rect 18052 32852 18104 32904
rect 19524 32929 19533 32963
rect 19533 32929 19567 32963
rect 19567 32929 19576 32963
rect 19524 32920 19576 32929
rect 18604 32852 18656 32904
rect 21640 32920 21692 32972
rect 21916 32920 21968 32972
rect 16856 32784 16908 32793
rect 20536 32784 20588 32836
rect 15200 32716 15252 32768
rect 18696 32759 18748 32768
rect 18696 32725 18705 32759
rect 18705 32725 18739 32759
rect 18739 32725 18748 32759
rect 18696 32716 18748 32725
rect 21824 32852 21876 32904
rect 22284 32852 22336 32904
rect 22744 32920 22796 32972
rect 23020 32920 23072 32972
rect 29552 33056 29604 33108
rect 30288 33056 30340 33108
rect 30656 33056 30708 33108
rect 29092 32988 29144 33040
rect 23112 32895 23164 32904
rect 23112 32861 23121 32895
rect 23121 32861 23155 32895
rect 23155 32861 23164 32895
rect 23112 32852 23164 32861
rect 23296 32852 23348 32904
rect 23848 32852 23900 32904
rect 25044 32852 25096 32904
rect 25228 32852 25280 32904
rect 26148 32852 26200 32904
rect 30656 32963 30708 32972
rect 30656 32929 30665 32963
rect 30665 32929 30699 32963
rect 30699 32929 30708 32963
rect 30656 32920 30708 32929
rect 26332 32784 26384 32836
rect 28080 32852 28132 32904
rect 28448 32852 28500 32904
rect 29000 32852 29052 32904
rect 29736 32852 29788 32904
rect 27988 32827 28040 32836
rect 27988 32793 27997 32827
rect 27997 32793 28031 32827
rect 28031 32793 28040 32827
rect 27988 32784 28040 32793
rect 23572 32759 23624 32768
rect 23572 32725 23581 32759
rect 23581 32725 23615 32759
rect 23615 32725 23624 32759
rect 23572 32716 23624 32725
rect 25780 32716 25832 32768
rect 27712 32716 27764 32768
rect 28724 32784 28776 32836
rect 30932 32852 30984 32904
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 31576 32784 31628 32836
rect 31944 32784 31996 32836
rect 47676 32784 47728 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 31024 32716 31076 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 16672 32512 16724 32564
rect 18604 32512 18656 32564
rect 24860 32512 24912 32564
rect 27620 32555 27672 32564
rect 27620 32521 27629 32555
rect 27629 32521 27663 32555
rect 27663 32521 27672 32555
rect 27620 32512 27672 32521
rect 31576 32555 31628 32564
rect 31576 32521 31585 32555
rect 31585 32521 31619 32555
rect 31619 32521 31628 32555
rect 31576 32512 31628 32521
rect 47676 32555 47728 32564
rect 47676 32521 47685 32555
rect 47685 32521 47719 32555
rect 47719 32521 47728 32555
rect 47676 32512 47728 32521
rect 2044 32487 2096 32496
rect 2044 32453 2053 32487
rect 2053 32453 2087 32487
rect 2087 32453 2096 32487
rect 2044 32444 2096 32453
rect 15936 32419 15988 32428
rect 1768 32308 1820 32360
rect 3240 32351 3292 32360
rect 3240 32317 3249 32351
rect 3249 32317 3283 32351
rect 3283 32317 3292 32351
rect 3240 32308 3292 32317
rect 15936 32385 15945 32419
rect 15945 32385 15979 32419
rect 15979 32385 15988 32419
rect 15936 32376 15988 32385
rect 14372 32240 14424 32292
rect 15660 32172 15712 32224
rect 16120 32240 16172 32292
rect 16672 32419 16724 32428
rect 16672 32385 16681 32419
rect 16681 32385 16715 32419
rect 16715 32385 16724 32419
rect 16672 32376 16724 32385
rect 16856 32240 16908 32292
rect 17408 32444 17460 32496
rect 23756 32444 23808 32496
rect 25872 32444 25924 32496
rect 26148 32444 26200 32496
rect 17316 32376 17368 32428
rect 18052 32419 18104 32428
rect 18052 32385 18061 32419
rect 18061 32385 18095 32419
rect 18095 32385 18104 32419
rect 18052 32376 18104 32385
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 19064 32419 19116 32428
rect 19064 32385 19073 32419
rect 19073 32385 19107 32419
rect 19107 32385 19116 32419
rect 19064 32376 19116 32385
rect 18604 32240 18656 32292
rect 18420 32215 18472 32224
rect 18420 32181 18429 32215
rect 18429 32181 18463 32215
rect 18463 32181 18472 32215
rect 18420 32172 18472 32181
rect 19340 32308 19392 32360
rect 19524 32376 19576 32428
rect 23572 32376 23624 32428
rect 20260 32308 20312 32360
rect 23480 32308 23532 32360
rect 24768 32376 24820 32428
rect 25780 32419 25832 32428
rect 25780 32385 25789 32419
rect 25789 32385 25823 32419
rect 25823 32385 25832 32419
rect 25780 32376 25832 32385
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 28264 32444 28316 32496
rect 30564 32444 30616 32496
rect 25044 32240 25096 32292
rect 27620 32376 27672 32428
rect 28632 32419 28684 32428
rect 28632 32385 28641 32419
rect 28641 32385 28675 32419
rect 28675 32385 28684 32419
rect 28632 32376 28684 32385
rect 29092 32376 29144 32428
rect 30840 32376 30892 32428
rect 31024 32419 31076 32428
rect 31024 32385 31034 32419
rect 31034 32385 31068 32419
rect 31068 32385 31076 32419
rect 31024 32376 31076 32385
rect 30472 32308 30524 32360
rect 31300 32419 31352 32428
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 47492 32444 47544 32496
rect 46296 32376 46348 32428
rect 44180 32308 44232 32360
rect 46664 32308 46716 32360
rect 20168 32172 20220 32224
rect 25872 32215 25924 32224
rect 25872 32181 25881 32215
rect 25881 32181 25915 32215
rect 25915 32181 25924 32215
rect 25872 32172 25924 32181
rect 28540 32172 28592 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1400 32011 1452 32020
rect 1400 31977 1409 32011
rect 1409 31977 1443 32011
rect 1443 31977 1452 32011
rect 1400 31968 1452 31977
rect 17776 31968 17828 32020
rect 16856 31900 16908 31952
rect 14740 31832 14792 31884
rect 15200 31875 15252 31884
rect 15200 31841 15209 31875
rect 15209 31841 15243 31875
rect 15243 31841 15252 31875
rect 15200 31832 15252 31841
rect 15936 31832 15988 31884
rect 17960 31943 18012 31952
rect 17960 31909 17969 31943
rect 17969 31909 18003 31943
rect 18003 31909 18012 31943
rect 19340 31968 19392 32020
rect 20352 31968 20404 32020
rect 20720 31968 20772 32020
rect 21732 31968 21784 32020
rect 28632 32011 28684 32020
rect 17960 31900 18012 31909
rect 18696 31900 18748 31952
rect 19984 31900 20036 31952
rect 20260 31900 20312 31952
rect 20996 31900 21048 31952
rect 28632 31977 28641 32011
rect 28641 31977 28675 32011
rect 28675 31977 28684 32011
rect 28632 31968 28684 31977
rect 30840 32011 30892 32020
rect 30840 31977 30849 32011
rect 30849 31977 30883 32011
rect 30883 31977 30892 32011
rect 30840 31968 30892 31977
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 2044 31764 2096 31816
rect 2964 31764 3016 31816
rect 15660 31696 15712 31748
rect 18052 31764 18104 31816
rect 19064 31764 19116 31816
rect 20904 31832 20956 31884
rect 21732 31832 21784 31884
rect 19524 31807 19576 31816
rect 19524 31773 19533 31807
rect 19533 31773 19567 31807
rect 19567 31773 19576 31807
rect 19524 31764 19576 31773
rect 20628 31807 20680 31816
rect 20628 31773 20637 31807
rect 20637 31773 20671 31807
rect 20671 31773 20680 31807
rect 20628 31764 20680 31773
rect 20812 31807 20864 31816
rect 20812 31773 20819 31807
rect 20819 31773 20864 31807
rect 20812 31764 20864 31773
rect 21088 31807 21140 31816
rect 21088 31773 21102 31807
rect 21102 31773 21136 31807
rect 21136 31773 21140 31807
rect 21088 31764 21140 31773
rect 18328 31696 18380 31748
rect 19340 31696 19392 31748
rect 20904 31739 20956 31748
rect 20904 31705 20913 31739
rect 20913 31705 20947 31739
rect 20947 31705 20956 31739
rect 20904 31696 20956 31705
rect 20996 31739 21048 31748
rect 20996 31705 21005 31739
rect 21005 31705 21039 31739
rect 21039 31705 21048 31739
rect 20996 31696 21048 31705
rect 2872 31671 2924 31680
rect 2872 31637 2881 31671
rect 2881 31637 2915 31671
rect 2915 31637 2924 31671
rect 2872 31628 2924 31637
rect 11704 31628 11756 31680
rect 16580 31628 16632 31680
rect 19984 31628 20036 31680
rect 20168 31628 20220 31680
rect 23848 31832 23900 31884
rect 27528 31900 27580 31952
rect 30932 31900 30984 31952
rect 27620 31832 27672 31884
rect 30472 31832 30524 31884
rect 47308 31875 47360 31884
rect 47308 31841 47317 31875
rect 47317 31841 47351 31875
rect 47351 31841 47360 31875
rect 47308 31832 47360 31841
rect 47492 31832 47544 31884
rect 22560 31764 22612 31816
rect 24768 31764 24820 31816
rect 25320 31764 25372 31816
rect 27160 31807 27212 31816
rect 27160 31773 27169 31807
rect 27169 31773 27203 31807
rect 27203 31773 27212 31807
rect 27160 31764 27212 31773
rect 28172 31764 28224 31816
rect 28448 31764 28500 31816
rect 29000 31764 29052 31816
rect 30656 31764 30708 31816
rect 31024 31807 31076 31816
rect 31024 31773 31033 31807
rect 31033 31773 31067 31807
rect 31067 31773 31076 31807
rect 31024 31764 31076 31773
rect 23756 31696 23808 31748
rect 27712 31696 27764 31748
rect 28264 31696 28316 31748
rect 26240 31628 26292 31680
rect 27528 31628 27580 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 16948 31424 17000 31476
rect 22284 31467 22336 31476
rect 22284 31433 22293 31467
rect 22293 31433 22327 31467
rect 22327 31433 22336 31467
rect 22284 31424 22336 31433
rect 23204 31424 23256 31476
rect 2872 31356 2924 31408
rect 16580 31356 16632 31408
rect 2044 31331 2096 31340
rect 2044 31297 2053 31331
rect 2053 31297 2087 31331
rect 2087 31297 2096 31331
rect 2044 31288 2096 31297
rect 18236 31331 18288 31340
rect 2780 31263 2832 31272
rect 2780 31229 2789 31263
rect 2789 31229 2823 31263
rect 2823 31229 2832 31263
rect 2780 31220 2832 31229
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 18328 31331 18380 31340
rect 18328 31297 18337 31331
rect 18337 31297 18371 31331
rect 18371 31297 18380 31331
rect 20352 31331 20404 31340
rect 18328 31288 18380 31297
rect 20352 31297 20361 31331
rect 20361 31297 20395 31331
rect 20395 31297 20404 31331
rect 20352 31288 20404 31297
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 26332 31356 26384 31408
rect 28172 31424 28224 31476
rect 22836 31331 22888 31340
rect 20168 31220 20220 31272
rect 22836 31297 22845 31331
rect 22845 31297 22879 31331
rect 22879 31297 22888 31331
rect 22836 31288 22888 31297
rect 23112 31288 23164 31340
rect 23204 31331 23256 31340
rect 23204 31297 23213 31331
rect 23213 31297 23247 31331
rect 23247 31297 23256 31331
rect 23204 31288 23256 31297
rect 24768 31288 24820 31340
rect 25136 31331 25188 31340
rect 25136 31297 25145 31331
rect 25145 31297 25179 31331
rect 25179 31297 25188 31331
rect 25136 31288 25188 31297
rect 28448 31356 28500 31408
rect 27528 31331 27580 31340
rect 20536 31152 20588 31204
rect 14280 31084 14332 31136
rect 19984 31084 20036 31136
rect 23572 31152 23624 31204
rect 27528 31297 27537 31331
rect 27537 31297 27571 31331
rect 27571 31297 27580 31331
rect 27528 31288 27580 31297
rect 30564 31288 30616 31340
rect 27804 31263 27856 31272
rect 27804 31229 27813 31263
rect 27813 31229 27847 31263
rect 27847 31229 27856 31263
rect 27804 31220 27856 31229
rect 31116 31331 31168 31340
rect 31116 31297 31125 31331
rect 31125 31297 31159 31331
rect 31159 31297 31168 31331
rect 31116 31288 31168 31297
rect 26516 31152 26568 31204
rect 20904 31127 20956 31136
rect 20904 31093 20913 31127
rect 20913 31093 20947 31127
rect 20947 31093 20956 31127
rect 20904 31084 20956 31093
rect 24400 31084 24452 31136
rect 25688 31084 25740 31136
rect 27344 31084 27396 31136
rect 29000 31084 29052 31136
rect 29276 31127 29328 31136
rect 29276 31093 29285 31127
rect 29285 31093 29319 31127
rect 29319 31093 29328 31127
rect 29276 31084 29328 31093
rect 31300 31084 31352 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19340 30880 19392 30932
rect 23756 30923 23808 30932
rect 23756 30889 23765 30923
rect 23765 30889 23799 30923
rect 23799 30889 23808 30923
rect 23756 30880 23808 30889
rect 26332 30880 26384 30932
rect 26976 30880 27028 30932
rect 27804 30880 27856 30932
rect 30564 30923 30616 30932
rect 30564 30889 30573 30923
rect 30573 30889 30607 30923
rect 30607 30889 30616 30923
rect 30564 30880 30616 30889
rect 16120 30719 16172 30728
rect 16120 30685 16129 30719
rect 16129 30685 16163 30719
rect 16163 30685 16172 30719
rect 16120 30676 16172 30685
rect 17592 30719 17644 30728
rect 17592 30685 17601 30719
rect 17601 30685 17635 30719
rect 17635 30685 17644 30719
rect 17592 30676 17644 30685
rect 17776 30744 17828 30796
rect 23204 30744 23256 30796
rect 18144 30676 18196 30728
rect 20352 30676 20404 30728
rect 20720 30676 20772 30728
rect 24400 30812 24452 30864
rect 28172 30812 28224 30864
rect 26700 30676 26752 30728
rect 28356 30719 28408 30728
rect 17040 30608 17092 30660
rect 17776 30651 17828 30660
rect 17776 30617 17785 30651
rect 17785 30617 17819 30651
rect 17819 30617 17828 30651
rect 17776 30608 17828 30617
rect 18420 30608 18472 30660
rect 16580 30540 16632 30592
rect 17408 30583 17460 30592
rect 17408 30549 17417 30583
rect 17417 30549 17451 30583
rect 17451 30549 17460 30583
rect 17408 30540 17460 30549
rect 20812 30608 20864 30660
rect 23388 30651 23440 30660
rect 21180 30540 21232 30592
rect 23388 30617 23397 30651
rect 23397 30617 23431 30651
rect 23431 30617 23440 30651
rect 23388 30608 23440 30617
rect 23572 30651 23624 30660
rect 23572 30617 23581 30651
rect 23581 30617 23615 30651
rect 23615 30617 23624 30651
rect 23572 30608 23624 30617
rect 24768 30651 24820 30660
rect 24768 30617 24777 30651
rect 24777 30617 24811 30651
rect 24811 30617 24820 30651
rect 24768 30608 24820 30617
rect 26792 30608 26844 30660
rect 28356 30685 28365 30719
rect 28365 30685 28399 30719
rect 28399 30685 28408 30719
rect 28356 30676 28408 30685
rect 28540 30719 28592 30728
rect 28540 30685 28547 30719
rect 28547 30685 28592 30719
rect 28540 30676 28592 30685
rect 30472 30744 30524 30796
rect 30012 30719 30064 30728
rect 30012 30685 30021 30719
rect 30021 30685 30055 30719
rect 30055 30685 30064 30719
rect 30012 30676 30064 30685
rect 30932 30744 30984 30796
rect 31300 30787 31352 30796
rect 31300 30753 31309 30787
rect 31309 30753 31343 30787
rect 31343 30753 31352 30787
rect 31300 30744 31352 30753
rect 28264 30608 28316 30660
rect 27252 30540 27304 30592
rect 29276 30608 29328 30660
rect 32312 30608 32364 30660
rect 31300 30540 31352 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17592 30336 17644 30388
rect 17776 30336 17828 30388
rect 16120 30200 16172 30252
rect 16764 30200 16816 30252
rect 18144 30243 18196 30252
rect 18144 30209 18153 30243
rect 18153 30209 18187 30243
rect 18187 30209 18196 30243
rect 18144 30200 18196 30209
rect 18420 30268 18472 30320
rect 18328 30243 18380 30252
rect 18328 30209 18337 30243
rect 18337 30209 18371 30243
rect 18371 30209 18380 30243
rect 20536 30336 20588 30388
rect 24584 30336 24636 30388
rect 28172 30336 28224 30388
rect 28356 30336 28408 30388
rect 30012 30336 30064 30388
rect 22284 30268 22336 30320
rect 23020 30268 23072 30320
rect 18328 30200 18380 30209
rect 20904 30243 20956 30252
rect 17776 30132 17828 30184
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 20812 30132 20864 30184
rect 17316 30107 17368 30116
rect 17316 30073 17325 30107
rect 17325 30073 17359 30107
rect 17359 30073 17368 30107
rect 17316 30064 17368 30073
rect 21180 30243 21232 30252
rect 21180 30209 21189 30243
rect 21189 30209 21223 30243
rect 21223 30209 21232 30243
rect 21180 30200 21232 30209
rect 23664 30200 23716 30252
rect 24400 30243 24452 30252
rect 24400 30209 24409 30243
rect 24409 30209 24443 30243
rect 24443 30209 24452 30243
rect 24400 30200 24452 30209
rect 24676 30243 24728 30252
rect 24676 30209 24685 30243
rect 24685 30209 24719 30243
rect 24719 30209 24728 30243
rect 24676 30200 24728 30209
rect 25228 30200 25280 30252
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 32312 30311 32364 30320
rect 32312 30277 32321 30311
rect 32321 30277 32355 30311
rect 32355 30277 32364 30311
rect 32312 30268 32364 30277
rect 27252 30200 27304 30252
rect 28908 30200 28960 30252
rect 23572 30132 23624 30184
rect 21180 30064 21232 30116
rect 25688 30175 25740 30184
rect 25688 30141 25697 30175
rect 25697 30141 25731 30175
rect 25731 30141 25740 30175
rect 25688 30132 25740 30141
rect 27436 30132 27488 30184
rect 28816 30132 28868 30184
rect 15936 29996 15988 30048
rect 17868 30039 17920 30048
rect 17868 30005 17877 30039
rect 17877 30005 17911 30039
rect 17911 30005 17920 30039
rect 17868 29996 17920 30005
rect 18328 29996 18380 30048
rect 19156 30039 19208 30048
rect 19156 30005 19165 30039
rect 19165 30005 19199 30039
rect 19199 30005 19208 30039
rect 19156 29996 19208 30005
rect 19340 29996 19392 30048
rect 20260 29996 20312 30048
rect 20996 29996 21048 30048
rect 25228 29996 25280 30048
rect 25412 30039 25464 30048
rect 25412 30005 25421 30039
rect 25421 30005 25455 30039
rect 25455 30005 25464 30039
rect 25412 29996 25464 30005
rect 26976 30064 27028 30116
rect 31300 30200 31352 30252
rect 33324 30200 33376 30252
rect 30840 30132 30892 30184
rect 47952 30064 48004 30116
rect 28264 29996 28316 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 16764 29835 16816 29844
rect 16764 29801 16773 29835
rect 16773 29801 16807 29835
rect 16807 29801 16816 29835
rect 16764 29792 16816 29801
rect 22192 29792 22244 29844
rect 25412 29792 25464 29844
rect 28448 29792 28500 29844
rect 29644 29792 29696 29844
rect 31852 29792 31904 29844
rect 21548 29724 21600 29776
rect 16028 29656 16080 29708
rect 17408 29656 17460 29708
rect 17776 29699 17828 29708
rect 17776 29665 17785 29699
rect 17785 29665 17819 29699
rect 17819 29665 17828 29699
rect 17776 29656 17828 29665
rect 20720 29656 20772 29708
rect 22008 29656 22060 29708
rect 17868 29588 17920 29640
rect 19984 29588 20036 29640
rect 22468 29631 22520 29640
rect 15292 29563 15344 29572
rect 15292 29529 15301 29563
rect 15301 29529 15335 29563
rect 15335 29529 15344 29563
rect 15292 29520 15344 29529
rect 15936 29520 15988 29572
rect 17316 29520 17368 29572
rect 17224 29495 17276 29504
rect 17224 29461 17233 29495
rect 17233 29461 17267 29495
rect 17267 29461 17276 29495
rect 17224 29452 17276 29461
rect 17500 29452 17552 29504
rect 17684 29452 17736 29504
rect 20996 29520 21048 29572
rect 22468 29597 22477 29631
rect 22477 29597 22511 29631
rect 22511 29597 22520 29631
rect 22468 29588 22520 29597
rect 23204 29588 23256 29640
rect 23664 29724 23716 29776
rect 24860 29724 24912 29776
rect 26700 29724 26752 29776
rect 27436 29724 27488 29776
rect 26240 29656 26292 29708
rect 26976 29656 27028 29708
rect 30564 29724 30616 29776
rect 23480 29588 23532 29640
rect 24676 29631 24728 29640
rect 24676 29597 24685 29631
rect 24685 29597 24719 29631
rect 24719 29597 24728 29631
rect 24676 29588 24728 29597
rect 27068 29588 27120 29640
rect 30840 29656 30892 29708
rect 31116 29588 31168 29640
rect 22100 29520 22152 29572
rect 23388 29520 23440 29572
rect 23572 29520 23624 29572
rect 25136 29520 25188 29572
rect 26976 29520 27028 29572
rect 27620 29563 27672 29572
rect 27620 29529 27629 29563
rect 27629 29529 27663 29563
rect 27663 29529 27672 29563
rect 27620 29520 27672 29529
rect 29828 29520 29880 29572
rect 30840 29520 30892 29572
rect 31392 29588 31444 29640
rect 45376 29656 45428 29708
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 21548 29452 21600 29504
rect 21824 29495 21876 29504
rect 21824 29461 21833 29495
rect 21833 29461 21867 29495
rect 21867 29461 21876 29495
rect 21824 29452 21876 29461
rect 23664 29452 23716 29504
rect 25228 29452 25280 29504
rect 29184 29452 29236 29504
rect 30288 29452 30340 29504
rect 30656 29495 30708 29504
rect 30656 29461 30665 29495
rect 30665 29461 30699 29495
rect 30699 29461 30708 29495
rect 30656 29452 30708 29461
rect 31208 29452 31260 29504
rect 31576 29452 31628 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2412 29248 2464 29300
rect 17224 29180 17276 29232
rect 16028 29112 16080 29164
rect 19340 29180 19392 29232
rect 20076 29180 20128 29232
rect 20720 29248 20772 29300
rect 22192 29248 22244 29300
rect 23388 29291 23440 29300
rect 23388 29257 23397 29291
rect 23397 29257 23431 29291
rect 23431 29257 23440 29291
rect 23388 29248 23440 29257
rect 23480 29248 23532 29300
rect 25044 29248 25096 29300
rect 26148 29248 26200 29300
rect 27160 29291 27212 29300
rect 27160 29257 27169 29291
rect 27169 29257 27203 29291
rect 27203 29257 27212 29291
rect 27160 29248 27212 29257
rect 26332 29180 26384 29232
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 20260 29044 20312 29096
rect 21548 29044 21600 29096
rect 22284 29112 22336 29164
rect 23020 29155 23072 29164
rect 22192 29087 22244 29096
rect 22192 29053 22201 29087
rect 22201 29053 22235 29087
rect 22235 29053 22244 29087
rect 22192 29044 22244 29053
rect 15292 28976 15344 29028
rect 21088 28976 21140 29028
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23204 29155 23256 29164
rect 23204 29121 23213 29155
rect 23213 29121 23247 29155
rect 23247 29121 23256 29155
rect 23204 29112 23256 29121
rect 24860 29112 24912 29164
rect 25596 29112 25648 29164
rect 30656 29180 30708 29232
rect 31576 29248 31628 29300
rect 32312 29248 32364 29300
rect 28816 29112 28868 29164
rect 30748 29112 30800 29164
rect 31208 29155 31260 29164
rect 31208 29121 31217 29155
rect 31217 29121 31251 29155
rect 31251 29121 31260 29155
rect 31208 29112 31260 29121
rect 23480 28976 23532 29028
rect 24584 28976 24636 29028
rect 25136 28976 25188 29028
rect 27620 28976 27672 29028
rect 28264 29019 28316 29028
rect 28264 28985 28273 29019
rect 28273 28985 28307 29019
rect 28307 28985 28316 29019
rect 28264 28976 28316 28985
rect 33416 29180 33468 29232
rect 32588 29087 32640 29096
rect 32588 29053 32597 29087
rect 32597 29053 32631 29087
rect 32631 29053 32640 29087
rect 32588 29044 32640 29053
rect 32864 29087 32916 29096
rect 32864 29053 32873 29087
rect 32873 29053 32907 29087
rect 32907 29053 32916 29087
rect 32864 29044 32916 29053
rect 19156 28908 19208 28960
rect 26884 28908 26936 28960
rect 29552 28908 29604 28960
rect 30012 28908 30064 28960
rect 30748 28908 30800 28960
rect 32036 28976 32088 29028
rect 31852 28908 31904 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 17684 28704 17736 28756
rect 22284 28704 22336 28756
rect 25320 28704 25372 28756
rect 26976 28704 27028 28756
rect 29644 28704 29696 28756
rect 31116 28747 31168 28756
rect 31116 28713 31125 28747
rect 31125 28713 31159 28747
rect 31159 28713 31168 28747
rect 31116 28704 31168 28713
rect 32864 28704 32916 28756
rect 33416 28747 33468 28756
rect 33416 28713 33425 28747
rect 33425 28713 33459 28747
rect 33459 28713 33468 28747
rect 33416 28704 33468 28713
rect 17040 28679 17092 28688
rect 17040 28645 17049 28679
rect 17049 28645 17083 28679
rect 17083 28645 17092 28679
rect 17040 28636 17092 28645
rect 44088 28704 44140 28756
rect 16028 28568 16080 28620
rect 21088 28568 21140 28620
rect 19340 28500 19392 28552
rect 22468 28568 22520 28620
rect 22744 28568 22796 28620
rect 23664 28568 23716 28620
rect 23572 28543 23624 28552
rect 23572 28509 23581 28543
rect 23581 28509 23615 28543
rect 23615 28509 23624 28543
rect 23572 28500 23624 28509
rect 24584 28500 24636 28552
rect 24860 28500 24912 28552
rect 16580 28432 16632 28484
rect 20812 28432 20864 28484
rect 22008 28475 22060 28484
rect 22008 28441 22017 28475
rect 22017 28441 22051 28475
rect 22051 28441 22060 28475
rect 22008 28432 22060 28441
rect 22560 28432 22612 28484
rect 26700 28568 26752 28620
rect 31392 28568 31444 28620
rect 32312 28611 32364 28620
rect 32312 28577 32321 28611
rect 32321 28577 32355 28611
rect 32355 28577 32364 28611
rect 32312 28568 32364 28577
rect 43996 28568 44048 28620
rect 25412 28500 25464 28552
rect 27068 28500 27120 28552
rect 27160 28500 27212 28552
rect 27988 28500 28040 28552
rect 28724 28500 28776 28552
rect 29092 28500 29144 28552
rect 29644 28543 29696 28552
rect 29644 28509 29653 28543
rect 29653 28509 29687 28543
rect 29687 28509 29696 28543
rect 29644 28500 29696 28509
rect 30012 28500 30064 28552
rect 30104 28500 30156 28552
rect 32036 28543 32088 28552
rect 32036 28509 32045 28543
rect 32045 28509 32079 28543
rect 32079 28509 32088 28543
rect 32036 28500 32088 28509
rect 23020 28364 23072 28416
rect 23204 28364 23256 28416
rect 25136 28364 25188 28416
rect 26056 28432 26108 28484
rect 26332 28364 26384 28416
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 29920 28407 29972 28416
rect 29920 28373 29929 28407
rect 29929 28373 29963 28407
rect 29963 28373 29972 28407
rect 29920 28364 29972 28373
rect 31208 28432 31260 28484
rect 32496 28500 32548 28552
rect 33324 28543 33376 28552
rect 33324 28509 33333 28543
rect 33333 28509 33367 28543
rect 33367 28509 33376 28543
rect 33324 28500 33376 28509
rect 32312 28364 32364 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 20076 28160 20128 28212
rect 20812 28203 20864 28212
rect 20812 28169 20821 28203
rect 20821 28169 20855 28203
rect 20855 28169 20864 28203
rect 20812 28160 20864 28169
rect 13452 28092 13504 28144
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 14188 28092 14240 28144
rect 14464 28092 14516 28144
rect 18052 28092 18104 28144
rect 22284 28135 22336 28144
rect 22284 28101 22293 28135
rect 22293 28101 22327 28135
rect 22327 28101 22336 28135
rect 22284 28092 22336 28101
rect 22744 28092 22796 28144
rect 25780 28160 25832 28212
rect 24584 28092 24636 28144
rect 25136 28092 25188 28144
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 8576 27999 8628 28008
rect 8576 27965 8585 27999
rect 8585 27965 8619 27999
rect 8619 27965 8628 27999
rect 8576 27956 8628 27965
rect 17960 28024 18012 28076
rect 19892 28067 19944 28076
rect 19892 28033 19901 28067
rect 19901 28033 19935 28067
rect 19935 28033 19944 28067
rect 19892 28024 19944 28033
rect 20812 28024 20864 28076
rect 22192 28067 22244 28076
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 22928 28024 22980 28076
rect 25228 28067 25280 28076
rect 25228 28033 25237 28067
rect 25237 28033 25271 28067
rect 25271 28033 25280 28067
rect 25228 28024 25280 28033
rect 26516 28092 26568 28144
rect 30196 28160 30248 28212
rect 23204 27999 23256 28008
rect 3976 27888 4028 27940
rect 23204 27965 23213 27999
rect 23213 27965 23247 27999
rect 23247 27965 23256 27999
rect 23204 27956 23256 27965
rect 24492 27956 24544 28008
rect 14556 27888 14608 27940
rect 15108 27888 15160 27940
rect 22836 27888 22888 27940
rect 15016 27863 15068 27872
rect 15016 27829 15025 27863
rect 15025 27829 15059 27863
rect 15059 27829 15068 27863
rect 15016 27820 15068 27829
rect 20720 27820 20772 27872
rect 22560 27820 22612 27872
rect 24676 27888 24728 27940
rect 26332 28067 26384 28076
rect 26332 28033 26341 28067
rect 26341 28033 26375 28067
rect 26375 28033 26384 28067
rect 26332 28024 26384 28033
rect 27712 28024 27764 28076
rect 28356 28024 28408 28076
rect 29092 28067 29144 28076
rect 29092 28033 29101 28067
rect 29101 28033 29135 28067
rect 29135 28033 29144 28067
rect 29092 28024 29144 28033
rect 29552 28067 29604 28076
rect 29552 28033 29561 28067
rect 29561 28033 29595 28067
rect 29595 28033 29604 28067
rect 29552 28024 29604 28033
rect 30288 28092 30340 28144
rect 30380 28067 30432 28076
rect 30380 28033 30389 28067
rect 30389 28033 30423 28067
rect 30423 28033 30432 28067
rect 30380 28024 30432 28033
rect 30932 28092 30984 28144
rect 28724 27956 28776 28008
rect 30196 27956 30248 28008
rect 31392 28067 31444 28076
rect 31392 28033 31401 28067
rect 31401 28033 31435 28067
rect 31435 28033 31444 28067
rect 31392 28024 31444 28033
rect 32772 28067 32824 28076
rect 32772 28033 32781 28067
rect 32781 28033 32815 28067
rect 32815 28033 32824 28067
rect 32772 28024 32824 28033
rect 36360 28067 36412 28076
rect 36360 28033 36369 28067
rect 36369 28033 36403 28067
rect 36403 28033 36412 28067
rect 36360 28024 36412 28033
rect 30932 27956 30984 28008
rect 37280 27999 37332 28008
rect 37280 27965 37289 27999
rect 37289 27965 37323 27999
rect 37323 27965 37332 27999
rect 37280 27956 37332 27965
rect 46848 27956 46900 28008
rect 26884 27888 26936 27940
rect 32496 27888 32548 27940
rect 32680 27888 32732 27940
rect 25044 27820 25096 27872
rect 25596 27820 25648 27872
rect 26148 27863 26200 27872
rect 26148 27829 26157 27863
rect 26157 27829 26191 27863
rect 26191 27829 26200 27863
rect 26148 27820 26200 27829
rect 28172 27820 28224 27872
rect 30932 27820 30984 27872
rect 31208 27863 31260 27872
rect 31208 27829 31217 27863
rect 31217 27829 31251 27863
rect 31251 27829 31260 27863
rect 31208 27820 31260 27829
rect 31300 27820 31352 27872
rect 33140 27820 33192 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8576 27616 8628 27668
rect 15016 27616 15068 27668
rect 15108 27616 15160 27668
rect 23572 27616 23624 27668
rect 26148 27616 26200 27668
rect 30380 27659 30432 27668
rect 30380 27625 30389 27659
rect 30389 27625 30423 27659
rect 30423 27625 30432 27659
rect 30380 27616 30432 27625
rect 37280 27659 37332 27668
rect 37280 27625 37289 27659
rect 37289 27625 37323 27659
rect 37323 27625 37332 27659
rect 37280 27616 37332 27625
rect 8392 27480 8444 27532
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 14648 27455 14700 27464
rect 9128 27387 9180 27396
rect 9128 27353 9137 27387
rect 9137 27353 9171 27387
rect 9171 27353 9180 27387
rect 9128 27344 9180 27353
rect 13360 27387 13412 27396
rect 13360 27353 13369 27387
rect 13369 27353 13403 27387
rect 13403 27353 13412 27387
rect 13360 27344 13412 27353
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 16212 27412 16264 27464
rect 20352 27548 20404 27600
rect 22192 27548 22244 27600
rect 25412 27548 25464 27600
rect 28264 27548 28316 27600
rect 20720 27480 20772 27532
rect 23480 27480 23532 27532
rect 24584 27480 24636 27532
rect 27712 27480 27764 27532
rect 20996 27455 21048 27464
rect 15200 27344 15252 27396
rect 16672 27344 16724 27396
rect 17132 27344 17184 27396
rect 18696 27387 18748 27396
rect 18696 27353 18705 27387
rect 18705 27353 18739 27387
rect 18739 27353 18748 27387
rect 18696 27344 18748 27353
rect 20076 27344 20128 27396
rect 9680 27276 9732 27328
rect 12716 27276 12768 27328
rect 13452 27319 13504 27328
rect 13452 27285 13461 27319
rect 13461 27285 13495 27319
rect 13495 27285 13504 27319
rect 13452 27276 13504 27285
rect 13544 27276 13596 27328
rect 13728 27276 13780 27328
rect 18880 27276 18932 27328
rect 20996 27421 21005 27455
rect 21005 27421 21039 27455
rect 21039 27421 21048 27455
rect 20996 27412 21048 27421
rect 21916 27455 21968 27464
rect 20812 27387 20864 27396
rect 20812 27353 20821 27387
rect 20821 27353 20855 27387
rect 20855 27353 20864 27387
rect 20812 27344 20864 27353
rect 21180 27344 21232 27396
rect 21916 27421 21925 27455
rect 21925 27421 21959 27455
rect 21959 27421 21968 27455
rect 21916 27412 21968 27421
rect 22928 27455 22980 27464
rect 22928 27421 22937 27455
rect 22937 27421 22971 27455
rect 22971 27421 22980 27455
rect 22928 27412 22980 27421
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 22100 27344 22152 27396
rect 25320 27412 25372 27464
rect 24400 27387 24452 27396
rect 24400 27353 24409 27387
rect 24409 27353 24443 27387
rect 24443 27353 24452 27387
rect 24400 27344 24452 27353
rect 25044 27344 25096 27396
rect 27068 27344 27120 27396
rect 28172 27455 28224 27464
rect 28172 27421 28181 27455
rect 28181 27421 28215 27455
rect 28215 27421 28224 27455
rect 32128 27480 32180 27532
rect 32588 27480 32640 27532
rect 28172 27412 28224 27421
rect 29644 27412 29696 27464
rect 29920 27344 29972 27396
rect 30012 27387 30064 27396
rect 30012 27353 30021 27387
rect 30021 27353 30055 27387
rect 30055 27353 30064 27387
rect 30012 27344 30064 27353
rect 31300 27344 31352 27396
rect 32496 27387 32548 27396
rect 32496 27353 32505 27387
rect 32505 27353 32539 27387
rect 32539 27353 32548 27387
rect 32496 27344 32548 27353
rect 33140 27344 33192 27396
rect 28172 27276 28224 27328
rect 30196 27276 30248 27328
rect 32404 27276 32456 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9128 27072 9180 27124
rect 14188 27072 14240 27124
rect 14464 27115 14516 27124
rect 14464 27081 14473 27115
rect 14473 27081 14507 27115
rect 14507 27081 14516 27115
rect 14464 27072 14516 27081
rect 14648 27072 14700 27124
rect 17132 27115 17184 27124
rect 17132 27081 17141 27115
rect 17141 27081 17175 27115
rect 17175 27081 17184 27115
rect 17132 27072 17184 27081
rect 18696 27072 18748 27124
rect 46572 27072 46624 27124
rect 12440 27004 12492 27056
rect 13728 27004 13780 27056
rect 14372 27004 14424 27056
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 10232 26936 10284 26988
rect 11520 26911 11572 26920
rect 11520 26877 11529 26911
rect 11529 26877 11563 26911
rect 11563 26877 11572 26911
rect 11520 26868 11572 26877
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 13728 26868 13780 26920
rect 14740 26936 14792 26988
rect 15292 27004 15344 27056
rect 18880 27047 18932 27056
rect 18880 27013 18889 27047
rect 18889 27013 18923 27047
rect 18923 27013 18932 27047
rect 18880 27004 18932 27013
rect 19892 27004 19944 27056
rect 21916 27004 21968 27056
rect 23020 27004 23072 27056
rect 27068 27047 27120 27056
rect 27068 27013 27077 27047
rect 27077 27013 27111 27047
rect 27111 27013 27120 27047
rect 27068 27004 27120 27013
rect 28172 27047 28224 27056
rect 28172 27013 28181 27047
rect 28181 27013 28215 27047
rect 28215 27013 28224 27047
rect 28172 27004 28224 27013
rect 29644 27004 29696 27056
rect 32496 27004 32548 27056
rect 15384 26936 15436 26988
rect 16948 26936 17000 26988
rect 13360 26800 13412 26852
rect 8944 26732 8996 26784
rect 13176 26732 13228 26784
rect 13728 26732 13780 26784
rect 21548 26868 21600 26920
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 23480 26936 23532 26988
rect 26976 26979 27028 26988
rect 26976 26945 26985 26979
rect 26985 26945 27019 26979
rect 27019 26945 27028 26979
rect 26976 26936 27028 26945
rect 30932 26936 30984 26988
rect 32312 26979 32364 26988
rect 32312 26945 32321 26979
rect 32321 26945 32355 26979
rect 32355 26945 32364 26979
rect 32312 26936 32364 26945
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32680 26979 32732 26988
rect 32404 26936 32456 26945
rect 32680 26945 32689 26979
rect 32689 26945 32723 26979
rect 32723 26945 32732 26979
rect 32680 26936 32732 26945
rect 22836 26868 22888 26920
rect 25320 26868 25372 26920
rect 27896 26911 27948 26920
rect 27896 26877 27905 26911
rect 27905 26877 27939 26911
rect 27939 26877 27948 26911
rect 27896 26868 27948 26877
rect 29736 26868 29788 26920
rect 32588 26868 32640 26920
rect 21640 26800 21692 26852
rect 21824 26800 21876 26852
rect 25044 26800 25096 26852
rect 19340 26732 19392 26784
rect 21180 26732 21232 26784
rect 22928 26775 22980 26784
rect 22928 26741 22937 26775
rect 22937 26741 22971 26775
rect 22971 26741 22980 26775
rect 22928 26732 22980 26741
rect 24400 26732 24452 26784
rect 30288 26732 30340 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2596 26528 2648 26580
rect 11796 26528 11848 26580
rect 27436 26528 27488 26580
rect 29644 26571 29696 26580
rect 8944 26435 8996 26444
rect 8944 26401 8953 26435
rect 8953 26401 8987 26435
rect 8987 26401 8996 26435
rect 8944 26392 8996 26401
rect 11612 26392 11664 26444
rect 13360 26392 13412 26444
rect 14096 26392 14148 26444
rect 16212 26460 16264 26512
rect 16672 26503 16724 26512
rect 16672 26469 16681 26503
rect 16681 26469 16715 26503
rect 16715 26469 16724 26503
rect 16672 26460 16724 26469
rect 19892 26503 19944 26512
rect 19892 26469 19901 26503
rect 19901 26469 19935 26503
rect 19935 26469 19944 26503
rect 19892 26460 19944 26469
rect 21456 26460 21508 26512
rect 21824 26460 21876 26512
rect 29644 26537 29653 26571
rect 29653 26537 29687 26571
rect 29687 26537 29696 26571
rect 29644 26528 29696 26537
rect 30472 26528 30524 26580
rect 31116 26571 31168 26580
rect 31116 26537 31125 26571
rect 31125 26537 31159 26571
rect 31159 26537 31168 26571
rect 31116 26528 31168 26537
rect 22560 26435 22612 26444
rect 12624 26324 12676 26376
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 15752 26324 15804 26376
rect 16580 26367 16632 26376
rect 16580 26333 16589 26367
rect 16589 26333 16623 26367
rect 16623 26333 16632 26367
rect 16580 26324 16632 26333
rect 19984 26324 20036 26376
rect 9220 26299 9272 26308
rect 9220 26265 9229 26299
rect 9229 26265 9263 26299
rect 9263 26265 9272 26299
rect 9220 26256 9272 26265
rect 9956 26256 10008 26308
rect 14648 26299 14700 26308
rect 14648 26265 14657 26299
rect 14657 26265 14691 26299
rect 14691 26265 14700 26299
rect 14648 26256 14700 26265
rect 21548 26324 21600 26376
rect 21824 26324 21876 26376
rect 22560 26401 22569 26435
rect 22569 26401 22603 26435
rect 22603 26401 22612 26435
rect 22560 26392 22612 26401
rect 22836 26435 22888 26444
rect 22836 26401 22845 26435
rect 22845 26401 22879 26435
rect 22879 26401 22888 26435
rect 22836 26392 22888 26401
rect 24492 26392 24544 26444
rect 25044 26324 25096 26376
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 27068 26324 27120 26376
rect 28080 26392 28132 26444
rect 27344 26367 27396 26376
rect 27344 26333 27353 26367
rect 27353 26333 27387 26367
rect 27387 26333 27396 26367
rect 27344 26324 27396 26333
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 8484 26188 8536 26240
rect 11796 26188 11848 26240
rect 12532 26188 12584 26240
rect 14096 26188 14148 26240
rect 23020 26256 23072 26308
rect 27252 26256 27304 26308
rect 28264 26299 28316 26308
rect 28264 26265 28273 26299
rect 28273 26265 28307 26299
rect 28307 26265 28316 26299
rect 28264 26256 28316 26265
rect 29460 26392 29512 26444
rect 29552 26367 29604 26376
rect 29552 26333 29561 26367
rect 29561 26333 29595 26367
rect 29595 26333 29604 26367
rect 29552 26324 29604 26333
rect 30564 26324 30616 26376
rect 31760 26367 31812 26376
rect 31760 26333 31769 26367
rect 31769 26333 31803 26367
rect 31803 26333 31812 26367
rect 31760 26324 31812 26333
rect 32312 26460 32364 26512
rect 40408 26392 40460 26444
rect 32036 26333 32045 26354
rect 32045 26333 32079 26354
rect 32079 26333 32088 26354
rect 32036 26302 32088 26333
rect 32680 26324 32732 26376
rect 22100 26188 22152 26240
rect 25412 26188 25464 26240
rect 25964 26188 26016 26240
rect 32496 26231 32548 26240
rect 32496 26197 32505 26231
rect 32505 26197 32539 26231
rect 32539 26197 32548 26231
rect 32496 26188 32548 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9220 25984 9272 26036
rect 9956 25984 10008 26036
rect 11612 26027 11664 26036
rect 11612 25993 11621 26027
rect 11621 25993 11655 26027
rect 11655 25993 11664 26027
rect 11612 25984 11664 25993
rect 11796 25984 11848 26036
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 14188 25984 14240 26036
rect 11704 25959 11756 25968
rect 11704 25925 11713 25959
rect 11713 25925 11747 25959
rect 11747 25925 11756 25959
rect 11704 25916 11756 25925
rect 8484 25891 8536 25900
rect 8484 25857 8493 25891
rect 8493 25857 8527 25891
rect 8527 25857 8536 25891
rect 8484 25848 8536 25857
rect 10048 25848 10100 25900
rect 10600 25848 10652 25900
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 14648 25984 14700 26036
rect 15752 25984 15804 26036
rect 31760 25984 31812 26036
rect 12532 25891 12584 25900
rect 11796 25848 11848 25857
rect 8576 25823 8628 25832
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 12624 25823 12676 25832
rect 12624 25789 12633 25823
rect 12633 25789 12667 25823
rect 12667 25789 12676 25823
rect 12992 25823 13044 25832
rect 12624 25780 12676 25789
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 13176 25848 13228 25900
rect 13176 25712 13228 25764
rect 13820 25780 13872 25832
rect 14924 25891 14976 25900
rect 14924 25857 14933 25891
rect 14933 25857 14967 25891
rect 14967 25857 14976 25891
rect 14924 25848 14976 25857
rect 15660 25848 15712 25900
rect 16580 25848 16632 25900
rect 19984 25848 20036 25900
rect 21088 25891 21140 25900
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 24860 25891 24912 25900
rect 16856 25823 16908 25832
rect 16856 25789 16865 25823
rect 16865 25789 16899 25823
rect 16899 25789 16908 25823
rect 16856 25780 16908 25789
rect 18880 25780 18932 25832
rect 19340 25780 19392 25832
rect 22100 25823 22152 25832
rect 22100 25789 22109 25823
rect 22109 25789 22143 25823
rect 22143 25789 22152 25823
rect 22100 25780 22152 25789
rect 22560 25780 22612 25832
rect 14096 25712 14148 25764
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 25596 25916 25648 25968
rect 25136 25848 25188 25900
rect 25044 25823 25096 25832
rect 25044 25789 25053 25823
rect 25053 25789 25087 25823
rect 25087 25789 25096 25823
rect 25412 25848 25464 25900
rect 30564 25916 30616 25968
rect 32496 25959 32548 25968
rect 26976 25891 27028 25900
rect 26976 25857 26985 25891
rect 26985 25857 27019 25891
rect 27019 25857 27028 25891
rect 26976 25848 27028 25857
rect 28816 25848 28868 25900
rect 29828 25848 29880 25900
rect 30840 25891 30892 25900
rect 30840 25857 30849 25891
rect 30849 25857 30883 25891
rect 30883 25857 30892 25891
rect 30840 25848 30892 25857
rect 32496 25925 32505 25959
rect 32505 25925 32539 25959
rect 32539 25925 32548 25959
rect 32496 25916 32548 25925
rect 33232 25916 33284 25968
rect 25044 25780 25096 25789
rect 32128 25780 32180 25832
rect 21088 25644 21140 25696
rect 25228 25644 25280 25696
rect 25596 25644 25648 25696
rect 25964 25687 26016 25696
rect 25964 25653 25973 25687
rect 25973 25653 26007 25687
rect 26007 25653 26016 25687
rect 25964 25644 26016 25653
rect 26884 25644 26936 25696
rect 27344 25644 27396 25696
rect 31484 25712 31536 25764
rect 31392 25644 31444 25696
rect 32036 25644 32088 25696
rect 46296 25644 46348 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 11520 25440 11572 25492
rect 12440 25483 12492 25492
rect 12440 25449 12449 25483
rect 12449 25449 12483 25483
rect 12483 25449 12492 25483
rect 14372 25483 14424 25492
rect 12440 25440 12492 25449
rect 14372 25449 14381 25483
rect 14381 25449 14415 25483
rect 14415 25449 14424 25483
rect 14372 25440 14424 25449
rect 16856 25483 16908 25492
rect 16856 25449 16865 25483
rect 16865 25449 16899 25483
rect 16899 25449 16908 25483
rect 16856 25440 16908 25449
rect 22100 25483 22152 25492
rect 22100 25449 22109 25483
rect 22109 25449 22143 25483
rect 22143 25449 22152 25483
rect 22100 25440 22152 25449
rect 25228 25440 25280 25492
rect 30840 25483 30892 25492
rect 10600 25372 10652 25424
rect 12532 25372 12584 25424
rect 12992 25372 13044 25424
rect 27068 25415 27120 25424
rect 27068 25381 27077 25415
rect 27077 25381 27111 25415
rect 27111 25381 27120 25415
rect 27068 25372 27120 25381
rect 9680 25304 9732 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 8576 25236 8628 25288
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 9588 25236 9640 25288
rect 10048 25236 10100 25288
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 11704 25304 11756 25356
rect 12716 25304 12768 25356
rect 14924 25304 14976 25356
rect 16580 25304 16632 25356
rect 11336 25279 11388 25288
rect 11336 25245 11345 25279
rect 11345 25245 11379 25279
rect 11379 25245 11388 25279
rect 12348 25279 12400 25288
rect 11336 25236 11388 25245
rect 12348 25245 12357 25279
rect 12357 25245 12391 25279
rect 12391 25245 12400 25279
rect 12348 25236 12400 25245
rect 14372 25279 14424 25288
rect 14372 25245 14381 25279
rect 14381 25245 14415 25279
rect 14415 25245 14424 25279
rect 14372 25236 14424 25245
rect 15384 25236 15436 25288
rect 16856 25236 16908 25288
rect 17960 25236 18012 25288
rect 18328 25279 18380 25288
rect 18328 25245 18337 25279
rect 18337 25245 18371 25279
rect 18371 25245 18380 25279
rect 18328 25236 18380 25245
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 21180 25304 21232 25356
rect 25596 25347 25648 25356
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 21548 25279 21600 25288
rect 21548 25245 21558 25279
rect 21558 25245 21592 25279
rect 21592 25245 21600 25279
rect 21548 25236 21600 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 25596 25313 25605 25347
rect 25605 25313 25639 25347
rect 25639 25313 25648 25347
rect 25596 25304 25648 25313
rect 30012 25372 30064 25424
rect 30840 25449 30849 25483
rect 30849 25449 30883 25483
rect 30883 25449 30892 25483
rect 30840 25440 30892 25449
rect 31392 25483 31444 25492
rect 31392 25449 31401 25483
rect 31401 25449 31435 25483
rect 31435 25449 31444 25483
rect 31392 25440 31444 25449
rect 31484 25440 31536 25492
rect 32772 25440 32824 25492
rect 33232 25483 33284 25492
rect 33232 25449 33241 25483
rect 33241 25449 33275 25483
rect 33275 25449 33284 25483
rect 33232 25440 33284 25449
rect 31852 25372 31904 25424
rect 31484 25304 31536 25356
rect 21732 25236 21784 25245
rect 24676 25279 24728 25288
rect 24676 25245 24685 25279
rect 24685 25245 24719 25279
rect 24719 25245 24728 25279
rect 24676 25236 24728 25245
rect 25136 25236 25188 25288
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 29460 25236 29512 25288
rect 17868 25168 17920 25220
rect 24860 25168 24912 25220
rect 26884 25168 26936 25220
rect 27620 25168 27672 25220
rect 29644 25236 29696 25288
rect 32036 25304 32088 25356
rect 46296 25347 46348 25356
rect 46296 25313 46305 25347
rect 46305 25313 46339 25347
rect 46339 25313 46348 25347
rect 46296 25304 46348 25313
rect 30288 25168 30340 25220
rect 9220 25100 9272 25152
rect 9956 25100 10008 25152
rect 18052 25100 18104 25152
rect 19340 25143 19392 25152
rect 19340 25109 19349 25143
rect 19349 25109 19383 25143
rect 19383 25109 19392 25143
rect 19340 25100 19392 25109
rect 24400 25100 24452 25152
rect 29920 25143 29972 25152
rect 29920 25109 29929 25143
rect 29929 25109 29963 25143
rect 29963 25109 29972 25143
rect 31852 25279 31904 25288
rect 31852 25245 31861 25279
rect 31861 25245 31895 25279
rect 31895 25245 31904 25279
rect 33140 25279 33192 25288
rect 31852 25236 31904 25245
rect 33140 25245 33149 25279
rect 33149 25245 33183 25279
rect 33183 25245 33192 25279
rect 33140 25236 33192 25245
rect 47676 25168 47728 25220
rect 48136 25211 48188 25220
rect 48136 25177 48145 25211
rect 48145 25177 48179 25211
rect 48179 25177 48188 25211
rect 48136 25168 48188 25177
rect 29920 25100 29972 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 24032 24939 24084 24948
rect 24032 24905 24041 24939
rect 24041 24905 24075 24939
rect 24075 24905 24084 24939
rect 24032 24896 24084 24905
rect 8484 24828 8536 24880
rect 14372 24871 14424 24880
rect 14372 24837 14381 24871
rect 14381 24837 14415 24871
rect 14415 24837 14424 24871
rect 14372 24828 14424 24837
rect 18052 24828 18104 24880
rect 19340 24828 19392 24880
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 11336 24760 11388 24812
rect 12532 24760 12584 24812
rect 12808 24803 12860 24812
rect 12808 24769 12817 24803
rect 12817 24769 12851 24803
rect 12851 24769 12860 24803
rect 12808 24760 12860 24769
rect 14096 24760 14148 24812
rect 25964 24896 26016 24948
rect 26976 24896 27028 24948
rect 24400 24871 24452 24880
rect 24400 24837 24409 24871
rect 24409 24837 24443 24871
rect 24443 24837 24452 24871
rect 24400 24828 24452 24837
rect 24860 24828 24912 24880
rect 25136 24828 25188 24880
rect 8208 24692 8260 24744
rect 16764 24735 16816 24744
rect 4804 24624 4856 24676
rect 16764 24701 16773 24735
rect 16773 24701 16807 24735
rect 16807 24701 16816 24735
rect 16764 24692 16816 24701
rect 17776 24692 17828 24744
rect 18972 24735 19024 24744
rect 18972 24701 18981 24735
rect 18981 24701 19015 24735
rect 19015 24701 19024 24735
rect 18972 24692 19024 24701
rect 20628 24692 20680 24744
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 24676 24803 24728 24812
rect 24676 24769 24685 24803
rect 24685 24769 24719 24803
rect 24719 24769 24728 24803
rect 24676 24760 24728 24769
rect 25228 24760 25280 24812
rect 26240 24760 26292 24812
rect 27344 24828 27396 24880
rect 26700 24760 26752 24812
rect 27620 24760 27672 24812
rect 29552 24828 29604 24880
rect 29736 24803 29788 24812
rect 25964 24692 26016 24744
rect 28632 24692 28684 24744
rect 29736 24769 29745 24803
rect 29745 24769 29779 24803
rect 29779 24769 29788 24803
rect 29736 24760 29788 24769
rect 30012 24760 30064 24812
rect 30104 24803 30156 24812
rect 30104 24769 30113 24803
rect 30113 24769 30147 24803
rect 30147 24769 30156 24803
rect 30104 24760 30156 24769
rect 33140 24760 33192 24812
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 3700 24556 3752 24608
rect 8576 24556 8628 24608
rect 8944 24556 8996 24608
rect 12624 24556 12676 24608
rect 15200 24556 15252 24608
rect 15844 24556 15896 24608
rect 18144 24556 18196 24608
rect 18512 24599 18564 24608
rect 18512 24565 18521 24599
rect 18521 24565 18555 24599
rect 18555 24565 18564 24599
rect 18512 24556 18564 24565
rect 24768 24624 24820 24676
rect 46756 24760 46808 24812
rect 45928 24692 45980 24744
rect 46112 24692 46164 24744
rect 47492 24760 47544 24812
rect 47676 24803 47728 24812
rect 47676 24769 47685 24803
rect 47685 24769 47719 24803
rect 47719 24769 47728 24803
rect 47676 24760 47728 24769
rect 20536 24556 20588 24608
rect 22836 24599 22888 24608
rect 22836 24565 22845 24599
rect 22845 24565 22879 24599
rect 22879 24565 22888 24599
rect 22836 24556 22888 24565
rect 24676 24556 24728 24608
rect 25228 24556 25280 24608
rect 28264 24556 28316 24608
rect 30012 24599 30064 24608
rect 30012 24565 30021 24599
rect 30021 24565 30055 24599
rect 30055 24565 30064 24599
rect 30012 24556 30064 24565
rect 30656 24599 30708 24608
rect 30656 24565 30665 24599
rect 30665 24565 30699 24599
rect 30699 24565 30708 24599
rect 30656 24556 30708 24565
rect 31024 24599 31076 24608
rect 31024 24565 31033 24599
rect 31033 24565 31067 24599
rect 31067 24565 31076 24599
rect 31024 24556 31076 24565
rect 32404 24556 32456 24608
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8208 24395 8260 24404
rect 8208 24361 8217 24395
rect 8217 24361 8251 24395
rect 8251 24361 8260 24395
rect 8208 24352 8260 24361
rect 9680 24352 9732 24404
rect 11704 24395 11756 24404
rect 11704 24361 11713 24395
rect 11713 24361 11747 24395
rect 11747 24361 11756 24395
rect 11704 24352 11756 24361
rect 18972 24352 19024 24404
rect 20628 24395 20680 24404
rect 20628 24361 20637 24395
rect 20637 24361 20671 24395
rect 20671 24361 20680 24395
rect 20628 24352 20680 24361
rect 14740 24284 14792 24336
rect 25044 24352 25096 24404
rect 25136 24352 25188 24404
rect 29460 24352 29512 24404
rect 30196 24352 30248 24404
rect 31024 24352 31076 24404
rect 31852 24352 31904 24404
rect 28816 24284 28868 24336
rect 30932 24284 30984 24336
rect 8944 24259 8996 24268
rect 8944 24225 8953 24259
rect 8953 24225 8987 24259
rect 8987 24225 8996 24259
rect 8944 24216 8996 24225
rect 9220 24259 9272 24268
rect 9220 24225 9229 24259
rect 9229 24225 9263 24259
rect 9263 24225 9272 24259
rect 9220 24216 9272 24225
rect 9588 24216 9640 24268
rect 12072 24216 12124 24268
rect 12624 24259 12676 24268
rect 12624 24225 12633 24259
rect 12633 24225 12667 24259
rect 12667 24225 12676 24259
rect 12624 24216 12676 24225
rect 15200 24216 15252 24268
rect 17408 24259 17460 24268
rect 17408 24225 17417 24259
rect 17417 24225 17451 24259
rect 17451 24225 17460 24259
rect 17408 24216 17460 24225
rect 17592 24216 17644 24268
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 10784 24148 10836 24200
rect 11704 24148 11756 24200
rect 9956 24080 10008 24132
rect 14832 24148 14884 24200
rect 14924 24148 14976 24200
rect 18144 24191 18196 24200
rect 18144 24157 18153 24191
rect 18153 24157 18187 24191
rect 18187 24157 18196 24191
rect 18144 24148 18196 24157
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 19340 24191 19392 24200
rect 19340 24157 19349 24191
rect 19349 24157 19383 24191
rect 19383 24157 19392 24191
rect 19340 24148 19392 24157
rect 15752 24123 15804 24132
rect 15752 24089 15761 24123
rect 15761 24089 15795 24123
rect 15795 24089 15804 24123
rect 15752 24080 15804 24089
rect 17960 24080 18012 24132
rect 20536 24148 20588 24200
rect 25320 24216 25372 24268
rect 27252 24259 27304 24268
rect 27252 24225 27261 24259
rect 27261 24225 27295 24259
rect 27295 24225 27304 24259
rect 27252 24216 27304 24225
rect 29920 24216 29972 24268
rect 31116 24259 31168 24268
rect 31116 24225 31125 24259
rect 31125 24225 31159 24259
rect 31159 24225 31168 24259
rect 31116 24216 31168 24225
rect 32128 24216 32180 24268
rect 26976 24191 27028 24200
rect 11244 24012 11296 24064
rect 11796 24012 11848 24064
rect 13452 24012 13504 24064
rect 19064 24012 19116 24064
rect 26976 24157 26985 24191
rect 26985 24157 27019 24191
rect 27019 24157 27028 24191
rect 26976 24148 27028 24157
rect 30104 24148 30156 24200
rect 40040 24352 40092 24404
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 46296 24191 46348 24200
rect 24676 24123 24728 24132
rect 24676 24089 24685 24123
rect 24685 24089 24719 24123
rect 24719 24089 24728 24123
rect 24676 24080 24728 24089
rect 26332 24080 26384 24132
rect 27988 24080 28040 24132
rect 22836 24012 22888 24064
rect 26700 24012 26752 24064
rect 27344 24012 27396 24064
rect 27896 24012 27948 24064
rect 30656 24080 30708 24132
rect 32404 24080 32456 24132
rect 46296 24157 46305 24191
rect 46305 24157 46339 24191
rect 46339 24157 46348 24191
rect 46296 24148 46348 24157
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 14740 23808 14792 23860
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 15660 23808 15712 23860
rect 16764 23808 16816 23860
rect 17776 23808 17828 23860
rect 18328 23808 18380 23860
rect 19064 23851 19116 23860
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 9588 23672 9640 23724
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 10784 23647 10836 23656
rect 10784 23613 10793 23647
rect 10793 23613 10827 23647
rect 10827 23613 10836 23647
rect 10784 23604 10836 23613
rect 9772 23468 9824 23520
rect 10048 23511 10100 23520
rect 10048 23477 10057 23511
rect 10057 23477 10091 23511
rect 10091 23477 10100 23511
rect 10048 23468 10100 23477
rect 11244 23536 11296 23588
rect 11704 23783 11756 23792
rect 11704 23749 11713 23783
rect 11713 23749 11747 23783
rect 11747 23749 11756 23783
rect 11704 23740 11756 23749
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 12532 23740 12584 23792
rect 13452 23783 13504 23792
rect 13452 23749 13461 23783
rect 13461 23749 13495 23783
rect 13495 23749 13504 23783
rect 13452 23740 13504 23749
rect 14004 23740 14056 23792
rect 19064 23817 19073 23851
rect 19073 23817 19107 23851
rect 19107 23817 19116 23851
rect 19064 23808 19116 23817
rect 19340 23808 19392 23860
rect 20812 23808 20864 23860
rect 26332 23851 26384 23860
rect 26332 23817 26341 23851
rect 26341 23817 26375 23851
rect 26375 23817 26384 23851
rect 26332 23808 26384 23817
rect 26976 23808 27028 23860
rect 14832 23672 14884 23724
rect 16948 23672 17000 23724
rect 17592 23672 17644 23724
rect 17868 23672 17920 23724
rect 17960 23715 18012 23724
rect 17960 23681 17969 23715
rect 17969 23681 18003 23715
rect 18003 23681 18012 23715
rect 17960 23672 18012 23681
rect 19340 23672 19392 23724
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 27896 23740 27948 23792
rect 12624 23604 12676 23656
rect 12808 23604 12860 23656
rect 13176 23647 13228 23656
rect 13176 23613 13185 23647
rect 13185 23613 13219 23647
rect 13219 23613 13228 23647
rect 13176 23604 13228 23613
rect 14096 23604 14148 23656
rect 20536 23672 20588 23724
rect 25044 23672 25096 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 11796 23468 11848 23520
rect 12072 23511 12124 23520
rect 12072 23477 12081 23511
rect 12081 23477 12115 23511
rect 12115 23477 12124 23511
rect 12072 23468 12124 23477
rect 16856 23536 16908 23588
rect 12716 23468 12768 23520
rect 18144 23468 18196 23520
rect 20352 23468 20404 23520
rect 20812 23468 20864 23520
rect 25044 23468 25096 23520
rect 26884 23672 26936 23724
rect 31116 23808 31168 23860
rect 29000 23740 29052 23792
rect 29920 23740 29972 23792
rect 29736 23672 29788 23724
rect 30656 23715 30708 23724
rect 30656 23681 30665 23715
rect 30665 23681 30699 23715
rect 30699 23681 30708 23715
rect 30932 23715 30984 23724
rect 30656 23672 30708 23681
rect 29460 23604 29512 23656
rect 29644 23604 29696 23656
rect 30932 23681 30941 23715
rect 30941 23681 30975 23715
rect 30975 23681 30984 23715
rect 30932 23672 30984 23681
rect 31392 23715 31444 23724
rect 31392 23681 31401 23715
rect 31401 23681 31435 23715
rect 31435 23681 31444 23715
rect 31392 23672 31444 23681
rect 47768 23808 47820 23860
rect 46296 23672 46348 23724
rect 46204 23647 46256 23656
rect 46204 23613 46213 23647
rect 46213 23613 46247 23647
rect 46247 23613 46256 23647
rect 46204 23604 46256 23613
rect 30012 23468 30064 23520
rect 30196 23468 30248 23520
rect 30380 23511 30432 23520
rect 30380 23477 30389 23511
rect 30389 23477 30423 23511
rect 30423 23477 30432 23511
rect 30380 23468 30432 23477
rect 45284 23536 45336 23588
rect 45468 23536 45520 23588
rect 31484 23511 31536 23520
rect 31484 23477 31493 23511
rect 31493 23477 31527 23511
rect 31527 23477 31536 23511
rect 31484 23468 31536 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 9956 23264 10008 23316
rect 12348 23264 12400 23316
rect 13176 23264 13228 23316
rect 15752 23307 15804 23316
rect 15752 23273 15761 23307
rect 15761 23273 15795 23307
rect 15795 23273 15804 23307
rect 15752 23264 15804 23273
rect 19616 23264 19668 23316
rect 22468 23264 22520 23316
rect 27988 23307 28040 23316
rect 27988 23273 27997 23307
rect 27997 23273 28031 23307
rect 28031 23273 28040 23307
rect 27988 23264 28040 23273
rect 29000 23264 29052 23316
rect 29460 23264 29512 23316
rect 31392 23264 31444 23316
rect 15660 23196 15712 23248
rect 31484 23196 31536 23248
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 9496 23103 9548 23112
rect 9496 23069 9505 23103
rect 9505 23069 9539 23103
rect 9539 23069 9548 23103
rect 9496 23060 9548 23069
rect 13084 23060 13136 23112
rect 14832 23060 14884 23112
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 16948 23103 17000 23112
rect 16948 23069 16957 23103
rect 16957 23069 16991 23103
rect 16991 23069 17000 23103
rect 16948 23060 17000 23069
rect 19984 23128 20036 23180
rect 19340 23060 19392 23112
rect 20536 23060 20588 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 22100 23060 22152 23112
rect 10048 22992 10100 23044
rect 18144 22992 18196 23044
rect 20996 23035 21048 23044
rect 20996 23001 21005 23035
rect 21005 23001 21039 23035
rect 21039 23001 21048 23035
rect 20996 22992 21048 23001
rect 24216 23128 24268 23180
rect 25412 23128 25464 23180
rect 23296 23060 23348 23112
rect 25044 23103 25096 23112
rect 25044 23069 25053 23103
rect 25053 23069 25087 23103
rect 25087 23069 25096 23103
rect 25044 23060 25096 23069
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 29552 22992 29604 23044
rect 11244 22967 11296 22976
rect 11244 22933 11253 22967
rect 11253 22933 11287 22967
rect 11287 22933 11296 22967
rect 11244 22924 11296 22933
rect 12348 22924 12400 22976
rect 13912 22924 13964 22976
rect 16672 22924 16724 22976
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 19248 22924 19300 22976
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 27160 22967 27212 22976
rect 27160 22933 27169 22967
rect 27169 22933 27203 22967
rect 27203 22933 27212 22967
rect 27160 22924 27212 22933
rect 30380 23128 30432 23180
rect 46756 23128 46808 23180
rect 46848 23171 46900 23180
rect 46848 23137 46857 23171
rect 46857 23137 46891 23171
rect 46891 23137 46900 23171
rect 46848 23128 46900 23137
rect 30288 23060 30340 23112
rect 30656 23103 30708 23112
rect 30656 23069 30665 23103
rect 30665 23069 30699 23103
rect 30699 23069 30708 23103
rect 30656 23060 30708 23069
rect 42800 23060 42852 23112
rect 45560 23060 45612 23112
rect 31208 22992 31260 23044
rect 47676 22992 47728 23044
rect 36360 22924 36412 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9496 22720 9548 22772
rect 14004 22763 14056 22772
rect 14004 22729 14013 22763
rect 14013 22729 14047 22763
rect 14047 22729 14056 22763
rect 14004 22720 14056 22729
rect 19064 22720 19116 22772
rect 17684 22652 17736 22704
rect 19984 22652 20036 22704
rect 20720 22720 20772 22772
rect 20996 22720 21048 22772
rect 47676 22763 47728 22772
rect 9680 22627 9732 22636
rect 9680 22593 9689 22627
rect 9689 22593 9723 22627
rect 9723 22593 9732 22627
rect 9680 22584 9732 22593
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 15844 22584 15896 22636
rect 16672 22627 16724 22636
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 19248 22584 19300 22636
rect 20352 22652 20404 22704
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 27160 22695 27212 22704
rect 27160 22661 27169 22695
rect 27169 22661 27203 22695
rect 27203 22661 27212 22695
rect 27160 22652 27212 22661
rect 47676 22729 47685 22763
rect 47685 22729 47719 22763
rect 47719 22729 47728 22763
rect 47676 22720 47728 22729
rect 37372 22652 37424 22704
rect 45376 22695 45428 22704
rect 45376 22661 45385 22695
rect 45385 22661 45419 22695
rect 45419 22661 45428 22695
rect 45376 22652 45428 22661
rect 12808 22448 12860 22500
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 22468 22584 22520 22636
rect 25044 22584 25096 22636
rect 43444 22627 43496 22636
rect 43444 22593 43453 22627
rect 43453 22593 43487 22627
rect 43487 22593 43496 22627
rect 43444 22584 43496 22593
rect 43720 22627 43772 22636
rect 43720 22593 43729 22627
rect 43729 22593 43763 22627
rect 43763 22593 43772 22627
rect 43720 22584 43772 22593
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 23204 22559 23256 22568
rect 23204 22525 23213 22559
rect 23213 22525 23247 22559
rect 23247 22525 23256 22559
rect 23204 22516 23256 22525
rect 25504 22516 25556 22568
rect 25964 22516 26016 22568
rect 26976 22559 27028 22568
rect 26976 22525 26985 22559
rect 26985 22525 27019 22559
rect 27019 22525 27028 22559
rect 26976 22516 27028 22525
rect 26608 22448 26660 22500
rect 44548 22516 44600 22568
rect 45560 22516 45612 22568
rect 46572 22559 46624 22568
rect 46572 22525 46581 22559
rect 46581 22525 46615 22559
rect 46615 22525 46624 22559
rect 46572 22516 46624 22525
rect 12992 22423 13044 22432
rect 12992 22389 13001 22423
rect 13001 22389 13035 22423
rect 13035 22389 13044 22423
rect 12992 22380 13044 22389
rect 15016 22380 15068 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 23204 22219 23256 22228
rect 23204 22185 23213 22219
rect 23213 22185 23247 22219
rect 23247 22185 23256 22219
rect 23204 22176 23256 22185
rect 2504 22040 2556 22092
rect 11244 22040 11296 22092
rect 15016 22083 15068 22092
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 15016 22040 15068 22049
rect 12624 21972 12676 22024
rect 14648 21972 14700 22024
rect 11060 21947 11112 21956
rect 11060 21913 11069 21947
rect 11069 21913 11103 21947
rect 11103 21913 11112 21947
rect 11060 21904 11112 21913
rect 12716 21947 12768 21956
rect 12716 21913 12725 21947
rect 12725 21913 12759 21947
rect 12759 21913 12768 21947
rect 12716 21904 12768 21913
rect 45284 22083 45336 22092
rect 45284 22049 45293 22083
rect 45293 22049 45327 22083
rect 45327 22049 45336 22083
rect 45284 22040 45336 22049
rect 45744 22040 45796 22092
rect 46848 22083 46900 22092
rect 46848 22049 46857 22083
rect 46857 22049 46891 22083
rect 46891 22049 46900 22083
rect 46848 22040 46900 22049
rect 16488 21972 16540 22024
rect 19064 21972 19116 22024
rect 20812 21972 20864 22024
rect 23296 21972 23348 22024
rect 23848 21972 23900 22024
rect 24584 21972 24636 22024
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 44180 22015 44232 22024
rect 19432 21947 19484 21956
rect 19432 21913 19441 21947
rect 19441 21913 19475 21947
rect 19475 21913 19484 21947
rect 19432 21904 19484 21913
rect 21272 21904 21324 21956
rect 44180 21981 44189 22015
rect 44189 21981 44223 22015
rect 44223 21981 44232 22015
rect 44180 21972 44232 21981
rect 44916 21972 44968 22024
rect 45376 21972 45428 22024
rect 26976 21904 27028 21956
rect 29000 21904 29052 21956
rect 40684 21904 40736 21956
rect 46020 21972 46072 22024
rect 47676 21904 47728 21956
rect 21364 21836 21416 21888
rect 25044 21836 25096 21888
rect 43720 21836 43772 21888
rect 44456 21879 44508 21888
rect 44456 21845 44465 21879
rect 44465 21845 44499 21879
rect 44499 21845 44508 21879
rect 44456 21836 44508 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11060 21632 11112 21684
rect 11980 21564 12032 21616
rect 12992 21564 13044 21616
rect 13912 21564 13964 21616
rect 9036 21428 9088 21480
rect 3608 21360 3660 21412
rect 9680 21428 9732 21480
rect 11060 21496 11112 21548
rect 11704 21496 11756 21548
rect 12808 21496 12860 21548
rect 15660 21496 15712 21548
rect 18144 21564 18196 21616
rect 20260 21632 20312 21684
rect 20628 21632 20680 21684
rect 22100 21632 22152 21684
rect 25044 21564 25096 21616
rect 40684 21564 40736 21616
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 14648 21428 14700 21480
rect 18420 21471 18472 21480
rect 12900 21360 12952 21412
rect 18420 21437 18429 21471
rect 18429 21437 18463 21471
rect 18463 21437 18472 21471
rect 18420 21428 18472 21437
rect 21548 21496 21600 21548
rect 23480 21496 23532 21548
rect 25596 21496 25648 21548
rect 44180 21632 44232 21684
rect 47676 21675 47728 21684
rect 47676 21641 47685 21675
rect 47685 21641 47719 21675
rect 47719 21641 47728 21675
rect 47676 21632 47728 21641
rect 43720 21496 43772 21548
rect 44456 21539 44508 21548
rect 44456 21505 44465 21539
rect 44465 21505 44499 21539
rect 44499 21505 44508 21539
rect 44456 21496 44508 21505
rect 44548 21539 44600 21548
rect 44548 21505 44557 21539
rect 44557 21505 44591 21539
rect 44591 21505 44600 21539
rect 44548 21496 44600 21505
rect 44916 21496 44968 21548
rect 45376 21496 45428 21548
rect 47584 21539 47636 21548
rect 47584 21505 47593 21539
rect 47593 21505 47627 21539
rect 47627 21505 47636 21539
rect 47584 21496 47636 21505
rect 20720 21428 20772 21480
rect 24032 21471 24084 21480
rect 24032 21437 24041 21471
rect 24041 21437 24075 21471
rect 24075 21437 24084 21471
rect 24032 21428 24084 21437
rect 10232 21335 10284 21344
rect 10232 21301 10241 21335
rect 10241 21301 10275 21335
rect 10275 21301 10284 21335
rect 10232 21292 10284 21301
rect 11612 21335 11664 21344
rect 11612 21301 11621 21335
rect 11621 21301 11655 21335
rect 11655 21301 11664 21335
rect 11612 21292 11664 21301
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 13084 21292 13136 21344
rect 19340 21292 19392 21344
rect 20536 21292 20588 21344
rect 23112 21360 23164 21412
rect 26976 21360 27028 21412
rect 46020 21360 46072 21412
rect 23296 21335 23348 21344
rect 23296 21301 23305 21335
rect 23305 21301 23339 21335
rect 23339 21301 23348 21335
rect 23296 21292 23348 21301
rect 24768 21292 24820 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 11980 21131 12032 21140
rect 3516 21020 3568 21072
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 12992 21088 13044 21140
rect 19432 21088 19484 21140
rect 24032 21088 24084 21140
rect 43720 21131 43772 21140
rect 43720 21097 43729 21131
rect 43729 21097 43763 21131
rect 43763 21097 43772 21131
rect 43720 21088 43772 21097
rect 44180 21088 44232 21140
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10232 20952 10284 20961
rect 12164 20952 12216 21004
rect 23112 21063 23164 21072
rect 20076 20952 20128 21004
rect 20352 20952 20404 21004
rect 21364 20995 21416 21004
rect 21364 20961 21373 20995
rect 21373 20961 21407 20995
rect 21407 20961 21416 20995
rect 21364 20952 21416 20961
rect 23112 21029 23121 21063
rect 23121 21029 23155 21063
rect 23155 21029 23164 21063
rect 23112 21020 23164 21029
rect 22928 20952 22980 21004
rect 26608 20995 26660 21004
rect 26608 20961 26617 20995
rect 26617 20961 26651 20995
rect 26651 20961 26660 20995
rect 26608 20952 26660 20961
rect 8484 20884 8536 20936
rect 9680 20884 9732 20936
rect 11612 20884 11664 20936
rect 12900 20884 12952 20936
rect 14096 20927 14148 20936
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 17776 20884 17828 20936
rect 20260 20884 20312 20936
rect 20720 20884 20772 20936
rect 23296 20884 23348 20936
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 29368 20952 29420 21004
rect 13636 20816 13688 20868
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 22100 20816 22152 20868
rect 25136 20816 25188 20868
rect 26332 20859 26384 20868
rect 26332 20825 26341 20859
rect 26341 20825 26375 20859
rect 26375 20825 26384 20859
rect 26332 20816 26384 20825
rect 31392 20859 31444 20868
rect 31392 20825 31401 20859
rect 31401 20825 31435 20859
rect 31435 20825 31444 20859
rect 31392 20816 31444 20825
rect 43904 20884 43956 20936
rect 44364 20884 44416 20936
rect 47216 20952 47268 21004
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 46296 20927 46348 20936
rect 46296 20893 46305 20927
rect 46305 20893 46339 20927
rect 46339 20893 46348 20927
rect 46296 20884 46348 20893
rect 44732 20816 44784 20868
rect 47676 20816 47728 20868
rect 28356 20748 28408 20800
rect 44456 20791 44508 20800
rect 44456 20757 44465 20791
rect 44465 20757 44499 20791
rect 44499 20757 44508 20791
rect 44456 20748 44508 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 3792 20544 3844 20596
rect 11980 20476 12032 20528
rect 7840 20408 7892 20460
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 13728 20544 13780 20596
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 15292 20544 15344 20596
rect 18420 20544 18472 20596
rect 20352 20544 20404 20596
rect 22100 20587 22152 20596
rect 22100 20553 22109 20587
rect 22109 20553 22143 20587
rect 22143 20553 22152 20587
rect 22100 20544 22152 20553
rect 26332 20544 26384 20596
rect 12164 20476 12216 20528
rect 13636 20476 13688 20528
rect 16856 20519 16908 20528
rect 16856 20485 16865 20519
rect 16865 20485 16899 20519
rect 16899 20485 16908 20519
rect 16856 20476 16908 20485
rect 20812 20476 20864 20528
rect 25044 20476 25096 20528
rect 25780 20476 25832 20528
rect 27804 20519 27856 20528
rect 11796 20408 11848 20417
rect 11888 20340 11940 20392
rect 11244 20272 11296 20324
rect 11704 20272 11756 20324
rect 4988 20204 5040 20256
rect 12164 20204 12216 20256
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 14832 20408 14884 20460
rect 20720 20408 20772 20460
rect 21088 20408 21140 20460
rect 21548 20408 21600 20460
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 24768 20451 24820 20460
rect 23480 20408 23532 20417
rect 24768 20417 24777 20451
rect 24777 20417 24811 20451
rect 24811 20417 24820 20451
rect 24768 20408 24820 20417
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 26608 20408 26660 20460
rect 27804 20485 27813 20519
rect 27813 20485 27847 20519
rect 27847 20485 27856 20519
rect 27804 20476 27856 20485
rect 29552 20408 29604 20460
rect 40684 20544 40736 20596
rect 42800 20408 42852 20460
rect 16580 20340 16632 20392
rect 17776 20340 17828 20392
rect 23664 20340 23716 20392
rect 24952 20383 25004 20392
rect 24952 20349 24961 20383
rect 24961 20349 24995 20383
rect 24995 20349 25004 20383
rect 24952 20340 25004 20349
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 29000 20383 29052 20392
rect 29000 20349 29009 20383
rect 29009 20349 29043 20383
rect 29043 20349 29052 20383
rect 29000 20340 29052 20349
rect 31392 20340 31444 20392
rect 39304 20383 39356 20392
rect 19248 20272 19300 20324
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 17132 20204 17184 20256
rect 22928 20272 22980 20324
rect 39304 20349 39313 20383
rect 39313 20349 39347 20383
rect 39347 20349 39356 20383
rect 39304 20340 39356 20349
rect 45928 20544 45980 20596
rect 47676 20587 47728 20596
rect 47676 20553 47685 20587
rect 47685 20553 47719 20587
rect 47719 20553 47728 20587
rect 47676 20544 47728 20553
rect 45468 20476 45520 20528
rect 45744 20476 45796 20528
rect 46940 20408 46992 20460
rect 19984 20204 20036 20256
rect 20536 20204 20588 20256
rect 23020 20204 23072 20256
rect 28264 20204 28316 20256
rect 30472 20247 30524 20256
rect 30472 20213 30481 20247
rect 30481 20213 30515 20247
rect 30515 20213 30524 20247
rect 30472 20204 30524 20213
rect 44180 20340 44232 20392
rect 44364 20340 44416 20392
rect 46572 20340 46624 20392
rect 47952 20340 48004 20392
rect 44456 20272 44508 20324
rect 43812 20204 43864 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 11980 20000 12032 20052
rect 15292 20000 15344 20052
rect 1768 19932 1820 19984
rect 17132 20000 17184 20052
rect 26608 20043 26660 20052
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 1768 19796 1820 19848
rect 10876 19796 10928 19848
rect 11888 19839 11940 19848
rect 11888 19805 11894 19839
rect 11894 19805 11928 19839
rect 11928 19805 11940 19839
rect 11888 19796 11940 19805
rect 11980 19796 12032 19848
rect 12164 19864 12216 19916
rect 20536 19864 20588 19916
rect 9680 19728 9732 19780
rect 3976 19660 4028 19712
rect 12164 19728 12216 19780
rect 14832 19796 14884 19848
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 16672 19796 16724 19848
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 21548 19839 21600 19848
rect 15568 19771 15620 19780
rect 15568 19737 15577 19771
rect 15577 19737 15611 19771
rect 15611 19737 15620 19771
rect 15568 19728 15620 19737
rect 19432 19728 19484 19780
rect 20168 19728 20220 19780
rect 11796 19660 11848 19712
rect 11980 19660 12032 19712
rect 12256 19660 12308 19712
rect 13820 19660 13872 19712
rect 15752 19660 15804 19712
rect 16580 19660 16632 19712
rect 17868 19703 17920 19712
rect 17868 19669 17877 19703
rect 17877 19669 17911 19703
rect 17911 19669 17920 19703
rect 17868 19660 17920 19669
rect 18052 19660 18104 19712
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 26608 20009 26617 20043
rect 26617 20009 26651 20043
rect 26651 20009 26660 20043
rect 26608 20000 26660 20009
rect 31392 19932 31444 19984
rect 44180 19932 44232 19984
rect 24768 19796 24820 19848
rect 26424 19839 26476 19848
rect 26424 19805 26433 19839
rect 26433 19805 26467 19839
rect 26467 19805 26476 19839
rect 27436 19839 27488 19848
rect 26424 19796 26476 19805
rect 27436 19805 27445 19839
rect 27445 19805 27479 19839
rect 27479 19805 27488 19839
rect 27436 19796 27488 19805
rect 27804 19864 27856 19916
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 44364 19907 44416 19916
rect 44364 19873 44373 19907
rect 44373 19873 44407 19907
rect 44407 19873 44416 19907
rect 44364 19864 44416 19873
rect 44456 19864 44508 19916
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 43812 19839 43864 19848
rect 25320 19728 25372 19780
rect 25412 19728 25464 19780
rect 27804 19728 27856 19780
rect 43812 19805 43821 19839
rect 43821 19805 43855 19839
rect 43855 19805 43864 19839
rect 43812 19796 43864 19805
rect 44824 19796 44876 19848
rect 45376 19864 45428 19916
rect 48044 19864 48096 19916
rect 31944 19728 31996 19780
rect 32128 19771 32180 19780
rect 32128 19737 32137 19771
rect 32137 19737 32171 19771
rect 32171 19737 32180 19771
rect 32128 19728 32180 19737
rect 40776 19771 40828 19780
rect 40776 19737 40785 19771
rect 40785 19737 40819 19771
rect 40819 19737 40828 19771
rect 40776 19728 40828 19737
rect 42432 19771 42484 19780
rect 42432 19737 42441 19771
rect 42441 19737 42475 19771
rect 42475 19737 42484 19771
rect 42432 19728 42484 19737
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 21548 19660 21600 19712
rect 26148 19660 26200 19712
rect 28356 19703 28408 19712
rect 28356 19669 28365 19703
rect 28365 19669 28399 19703
rect 28399 19669 28408 19703
rect 28356 19660 28408 19669
rect 40592 19660 40644 19712
rect 48044 19728 48096 19780
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 11888 19499 11940 19508
rect 11888 19465 11897 19499
rect 11897 19465 11931 19499
rect 11931 19465 11940 19499
rect 11888 19456 11940 19465
rect 16672 19456 16724 19508
rect 11244 19388 11296 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 11060 19320 11112 19372
rect 11888 19320 11940 19372
rect 12348 19363 12400 19372
rect 12348 19329 12357 19363
rect 12357 19329 12391 19363
rect 12391 19329 12400 19363
rect 12348 19320 12400 19329
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 12164 19252 12216 19304
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 15936 19320 15988 19372
rect 19248 19456 19300 19508
rect 17868 19431 17920 19440
rect 17868 19397 17877 19431
rect 17877 19397 17911 19431
rect 17911 19397 17920 19431
rect 17868 19388 17920 19397
rect 16028 19252 16080 19304
rect 20996 19456 21048 19508
rect 21088 19456 21140 19508
rect 27620 19456 27672 19508
rect 28080 19499 28132 19508
rect 28080 19465 28089 19499
rect 28089 19465 28123 19499
rect 28123 19465 28132 19499
rect 28080 19456 28132 19465
rect 31944 19456 31996 19508
rect 40592 19456 40644 19508
rect 40776 19499 40828 19508
rect 40776 19465 40785 19499
rect 40785 19465 40819 19499
rect 40819 19465 40828 19499
rect 40776 19456 40828 19465
rect 44088 19456 44140 19508
rect 45836 19456 45888 19508
rect 46480 19456 46532 19508
rect 20352 19388 20404 19440
rect 21824 19431 21876 19440
rect 20812 19320 20864 19372
rect 21824 19397 21833 19431
rect 21833 19397 21867 19431
rect 21867 19397 21876 19431
rect 21824 19388 21876 19397
rect 23020 19431 23072 19440
rect 23020 19397 23029 19431
rect 23029 19397 23063 19431
rect 23063 19397 23072 19431
rect 23020 19388 23072 19397
rect 25228 19363 25280 19372
rect 18052 19252 18104 19304
rect 20536 19295 20588 19304
rect 3424 19184 3476 19236
rect 11796 19116 11848 19168
rect 12900 19116 12952 19168
rect 15568 19184 15620 19236
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 25228 19329 25237 19363
rect 25237 19329 25271 19363
rect 25271 19329 25280 19363
rect 25228 19320 25280 19329
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 26424 19320 26476 19372
rect 21824 19252 21876 19304
rect 22928 19295 22980 19304
rect 22928 19261 22937 19295
rect 22937 19261 22971 19295
rect 22971 19261 22980 19295
rect 22928 19252 22980 19261
rect 23756 19295 23808 19304
rect 23756 19261 23765 19295
rect 23765 19261 23799 19295
rect 23799 19261 23808 19295
rect 23756 19252 23808 19261
rect 24860 19252 24912 19304
rect 28448 19320 28500 19372
rect 28724 19320 28776 19372
rect 43260 19388 43312 19440
rect 40684 19363 40736 19372
rect 40684 19329 40693 19363
rect 40693 19329 40727 19363
rect 40727 19329 40736 19363
rect 47584 19388 47636 19440
rect 43904 19363 43956 19372
rect 40684 19320 40736 19329
rect 43904 19329 43913 19363
rect 43913 19329 43947 19363
rect 43947 19329 43956 19363
rect 43904 19320 43956 19329
rect 44088 19363 44140 19372
rect 44088 19329 44097 19363
rect 44097 19329 44131 19363
rect 44131 19329 44140 19363
rect 44088 19320 44140 19329
rect 44180 19320 44232 19372
rect 45008 19363 45060 19372
rect 45008 19329 45017 19363
rect 45017 19329 45051 19363
rect 45051 19329 45060 19363
rect 45008 19320 45060 19329
rect 27988 19252 28040 19304
rect 28816 19252 28868 19304
rect 44272 19252 44324 19304
rect 45560 19295 45612 19304
rect 45560 19261 45569 19295
rect 45569 19261 45603 19295
rect 45603 19261 45612 19295
rect 45560 19252 45612 19261
rect 46296 19252 46348 19304
rect 20720 19184 20772 19236
rect 44180 19184 44232 19236
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 21088 19116 21140 19168
rect 46296 19116 46348 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 11888 18912 11940 18964
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 13636 18912 13688 18964
rect 15292 18912 15344 18964
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 21824 18912 21876 18964
rect 27988 18955 28040 18964
rect 27988 18921 27997 18955
rect 27997 18921 28031 18955
rect 28031 18921 28040 18955
rect 27988 18912 28040 18921
rect 31944 18955 31996 18964
rect 31944 18921 31953 18955
rect 31953 18921 31987 18955
rect 31987 18921 31996 18955
rect 31944 18912 31996 18921
rect 44272 18955 44324 18964
rect 44272 18921 44281 18955
rect 44281 18921 44315 18955
rect 44315 18921 44324 18955
rect 44272 18912 44324 18921
rect 11980 18776 12032 18828
rect 16028 18844 16080 18896
rect 19984 18844 20036 18896
rect 24860 18844 24912 18896
rect 27804 18887 27856 18896
rect 27804 18853 27813 18887
rect 27813 18853 27847 18887
rect 27847 18853 27856 18887
rect 27804 18844 27856 18853
rect 2320 18708 2372 18760
rect 7564 18708 7616 18760
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 12256 18708 12308 18760
rect 11796 18683 11848 18692
rect 11796 18649 11805 18683
rect 11805 18649 11839 18683
rect 11839 18649 11848 18683
rect 11796 18640 11848 18649
rect 14832 18708 14884 18760
rect 15752 18708 15804 18760
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 23756 18776 23808 18828
rect 25228 18776 25280 18828
rect 28448 18819 28500 18828
rect 28448 18785 28457 18819
rect 28457 18785 28491 18819
rect 28491 18785 28500 18819
rect 28448 18776 28500 18785
rect 19432 18708 19484 18760
rect 19984 18708 20036 18760
rect 24492 18751 24544 18760
rect 13912 18640 13964 18692
rect 14556 18640 14608 18692
rect 18236 18683 18288 18692
rect 18236 18649 18245 18683
rect 18245 18649 18279 18683
rect 18279 18649 18288 18683
rect 20812 18683 20864 18692
rect 18236 18640 18288 18649
rect 20812 18649 20821 18683
rect 20821 18649 20855 18683
rect 20855 18649 20864 18683
rect 20812 18640 20864 18649
rect 21548 18640 21600 18692
rect 24492 18717 24501 18751
rect 24501 18717 24535 18751
rect 24535 18717 24544 18751
rect 24492 18708 24544 18717
rect 24676 18708 24728 18760
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 27620 18708 27672 18760
rect 28724 18708 28776 18760
rect 46296 18819 46348 18828
rect 46296 18785 46305 18819
rect 46305 18785 46339 18819
rect 46339 18785 46348 18819
rect 46296 18776 46348 18785
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 43260 18751 43312 18760
rect 43260 18717 43269 18751
rect 43269 18717 43303 18751
rect 43303 18717 43312 18751
rect 43260 18708 43312 18717
rect 44180 18751 44232 18760
rect 25228 18683 25280 18692
rect 25228 18649 25237 18683
rect 25237 18649 25271 18683
rect 25271 18649 25280 18683
rect 25228 18640 25280 18649
rect 27804 18640 27856 18692
rect 28816 18640 28868 18692
rect 44180 18717 44189 18751
rect 44189 18717 44223 18751
rect 44223 18717 44232 18751
rect 44180 18708 44232 18717
rect 44916 18708 44968 18760
rect 45192 18751 45244 18760
rect 45192 18717 45201 18751
rect 45201 18717 45235 18751
rect 45235 18717 45244 18751
rect 45192 18708 45244 18717
rect 45100 18640 45152 18692
rect 47676 18640 47728 18692
rect 11244 18572 11296 18624
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13820 18572 13872 18624
rect 14740 18572 14792 18624
rect 15476 18572 15528 18624
rect 20628 18572 20680 18624
rect 26240 18572 26292 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7564 18300 7616 18352
rect 12532 18300 12584 18352
rect 12900 18343 12952 18352
rect 12900 18309 12909 18343
rect 12909 18309 12943 18343
rect 12943 18309 12952 18343
rect 12900 18300 12952 18309
rect 13452 18300 13504 18352
rect 19984 18368 20036 18420
rect 20812 18368 20864 18420
rect 20076 18300 20128 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 11888 18275 11940 18284
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 15936 18275 15988 18284
rect 11980 18232 12032 18241
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 4896 18096 4948 18148
rect 11796 18164 11848 18216
rect 12624 18207 12676 18216
rect 12348 18096 12400 18148
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 18052 18232 18104 18284
rect 19432 18232 19484 18284
rect 20996 18300 21048 18352
rect 27896 18368 27948 18420
rect 47676 18411 47728 18420
rect 27620 18343 27672 18352
rect 20720 18232 20772 18284
rect 21824 18232 21876 18284
rect 25780 18275 25832 18284
rect 25780 18241 25789 18275
rect 25789 18241 25823 18275
rect 25823 18241 25832 18275
rect 25780 18232 25832 18241
rect 27620 18309 27629 18343
rect 27629 18309 27663 18343
rect 27663 18309 27672 18343
rect 27620 18300 27672 18309
rect 27436 18275 27488 18284
rect 27436 18241 27445 18275
rect 27445 18241 27479 18275
rect 27479 18241 27488 18275
rect 28080 18275 28132 18284
rect 27436 18232 27488 18241
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 18604 18164 18656 18216
rect 20168 18164 20220 18216
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 25136 18207 25188 18216
rect 25136 18173 25145 18207
rect 25145 18173 25179 18207
rect 25179 18173 25188 18207
rect 25136 18164 25188 18173
rect 26332 18164 26384 18216
rect 28264 18207 28316 18216
rect 28264 18173 28273 18207
rect 28273 18173 28307 18207
rect 28307 18173 28316 18207
rect 28264 18164 28316 18173
rect 29920 18207 29972 18216
rect 29920 18173 29929 18207
rect 29929 18173 29963 18207
rect 29963 18173 29972 18207
rect 29920 18164 29972 18173
rect 25412 18096 25464 18148
rect 44180 18275 44232 18284
rect 44180 18241 44189 18275
rect 44189 18241 44223 18275
rect 44223 18241 44232 18275
rect 44180 18232 44232 18241
rect 45008 18300 45060 18352
rect 44916 18275 44968 18284
rect 44916 18241 44925 18275
rect 44925 18241 44959 18275
rect 44959 18241 44968 18275
rect 44916 18232 44968 18241
rect 45928 18275 45980 18284
rect 45928 18241 45937 18275
rect 45937 18241 45971 18275
rect 45971 18241 45980 18275
rect 45928 18232 45980 18241
rect 44456 18164 44508 18216
rect 46848 18232 46900 18284
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 47400 18232 47452 18284
rect 44824 18096 44876 18148
rect 21456 18028 21508 18080
rect 25596 18028 25648 18080
rect 25872 18071 25924 18080
rect 25872 18037 25881 18071
rect 25881 18037 25915 18071
rect 25915 18037 25924 18071
rect 25872 18028 25924 18037
rect 45100 18028 45152 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 12624 17867 12676 17876
rect 2136 17756 2188 17808
rect 8760 17756 8812 17808
rect 12624 17833 12633 17867
rect 12633 17833 12667 17867
rect 12667 17833 12676 17867
rect 12624 17824 12676 17833
rect 15936 17824 15988 17876
rect 18236 17824 18288 17876
rect 23480 17867 23532 17876
rect 23480 17833 23489 17867
rect 23489 17833 23523 17867
rect 23523 17833 23532 17867
rect 23480 17824 23532 17833
rect 28264 17824 28316 17876
rect 44456 17867 44508 17876
rect 44456 17833 44465 17867
rect 44465 17833 44499 17867
rect 44499 17833 44508 17867
rect 44456 17824 44508 17833
rect 44916 17824 44968 17876
rect 3976 17688 4028 17740
rect 9036 17731 9088 17740
rect 9036 17697 9045 17731
rect 9045 17697 9079 17731
rect 9079 17697 9088 17731
rect 9036 17688 9088 17697
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 8484 17620 8536 17672
rect 8576 17620 8628 17672
rect 1952 17484 2004 17536
rect 14464 17688 14516 17740
rect 44640 17756 44692 17808
rect 47400 17756 47452 17808
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 12348 17620 12400 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 10508 17552 10560 17604
rect 11244 17552 11296 17604
rect 11888 17484 11940 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 17592 17620 17644 17672
rect 19340 17620 19392 17672
rect 25872 17731 25924 17740
rect 25872 17697 25878 17731
rect 25878 17697 25912 17731
rect 25912 17697 25924 17731
rect 26148 17731 26200 17740
rect 25872 17688 25924 17697
rect 26148 17697 26157 17731
rect 26157 17697 26191 17731
rect 26191 17697 26200 17731
rect 26148 17688 26200 17697
rect 20996 17620 21048 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 19248 17484 19300 17536
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 19984 17484 20036 17536
rect 22100 17552 22152 17604
rect 23296 17620 23348 17672
rect 23664 17620 23716 17672
rect 44088 17663 44140 17672
rect 26240 17552 26292 17604
rect 23020 17484 23072 17536
rect 25780 17484 25832 17536
rect 44088 17629 44097 17663
rect 44097 17629 44131 17663
rect 44131 17629 44140 17663
rect 44088 17620 44140 17629
rect 44272 17663 44324 17672
rect 44272 17629 44281 17663
rect 44281 17629 44315 17663
rect 44315 17629 44324 17663
rect 44272 17620 44324 17629
rect 45100 17620 45152 17672
rect 46296 17663 46348 17672
rect 46296 17629 46305 17663
rect 46305 17629 46339 17663
rect 46339 17629 46348 17663
rect 46296 17620 46348 17629
rect 45192 17595 45244 17604
rect 45192 17561 45201 17595
rect 45201 17561 45235 17595
rect 45235 17561 45244 17595
rect 45192 17552 45244 17561
rect 47676 17552 47728 17604
rect 48136 17595 48188 17604
rect 48136 17561 48145 17595
rect 48145 17561 48179 17595
rect 48179 17561 48188 17595
rect 48136 17552 48188 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 20 17280 72 17332
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 9956 17280 10008 17332
rect 10692 17280 10744 17332
rect 2044 17076 2096 17128
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 12440 17212 12492 17264
rect 20996 17212 21048 17264
rect 22100 17280 22152 17332
rect 22652 17280 22704 17332
rect 26148 17280 26200 17332
rect 45928 17280 45980 17332
rect 47676 17323 47728 17332
rect 47676 17289 47685 17323
rect 47685 17289 47719 17323
rect 47719 17289 47728 17323
rect 47676 17280 47728 17289
rect 23020 17255 23072 17264
rect 23020 17221 23029 17255
rect 23029 17221 23063 17255
rect 23063 17221 23072 17255
rect 23020 17212 23072 17221
rect 43536 17212 43588 17264
rect 44088 17212 44140 17264
rect 12348 17144 12400 17196
rect 14280 17144 14332 17196
rect 15476 17144 15528 17196
rect 16856 17144 16908 17196
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 22284 17144 22336 17196
rect 26240 17144 26292 17196
rect 44272 17187 44324 17196
rect 44272 17153 44281 17187
rect 44281 17153 44315 17187
rect 44315 17153 44324 17187
rect 44272 17144 44324 17153
rect 46296 17144 46348 17196
rect 47400 17144 47452 17196
rect 8116 17119 8168 17128
rect 8116 17085 8125 17119
rect 8125 17085 8159 17119
rect 8159 17085 8168 17119
rect 8116 17076 8168 17085
rect 9036 17076 9088 17128
rect 11980 17076 12032 17128
rect 12532 17076 12584 17128
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 20260 17076 20312 17128
rect 8484 17008 8536 17060
rect 15936 17008 15988 17060
rect 3976 16940 4028 16992
rect 12716 16940 12768 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14648 16940 14700 16992
rect 15660 16940 15712 16992
rect 17040 16940 17092 16992
rect 19340 16940 19392 16992
rect 23572 17076 23624 17128
rect 27252 17076 27304 17128
rect 29000 17076 29052 17128
rect 46572 17076 46624 17128
rect 46664 17008 46716 17060
rect 22100 16940 22152 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 8116 16736 8168 16788
rect 13636 16736 13688 16788
rect 17776 16736 17828 16788
rect 18144 16736 18196 16788
rect 19248 16668 19300 16720
rect 47492 16668 47544 16720
rect 8208 16600 8260 16652
rect 14464 16600 14516 16652
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 14924 16643 14976 16652
rect 14924 16609 14933 16643
rect 14933 16609 14967 16643
rect 14967 16609 14976 16643
rect 14924 16600 14976 16609
rect 16396 16643 16448 16652
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 29000 16600 29052 16652
rect 47768 16600 47820 16652
rect 11980 16575 12032 16584
rect 11336 16507 11388 16516
rect 11336 16473 11345 16507
rect 11345 16473 11379 16507
rect 11379 16473 11388 16507
rect 11336 16464 11388 16473
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 13268 16532 13320 16584
rect 18420 16532 18472 16584
rect 19984 16532 20036 16584
rect 21732 16532 21784 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 23388 16532 23440 16584
rect 27344 16575 27396 16584
rect 27344 16541 27353 16575
rect 27353 16541 27387 16575
rect 27387 16541 27396 16575
rect 27344 16532 27396 16541
rect 12348 16464 12400 16516
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 15660 16464 15712 16516
rect 18696 16507 18748 16516
rect 18696 16473 18705 16507
rect 18705 16473 18739 16507
rect 18739 16473 18748 16507
rect 18696 16464 18748 16473
rect 20168 16464 20220 16516
rect 21456 16464 21508 16516
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 15108 16396 15160 16448
rect 26056 16464 26108 16516
rect 40684 16464 40736 16516
rect 46756 16464 46808 16516
rect 48136 16507 48188 16516
rect 48136 16473 48145 16507
rect 48145 16473 48179 16507
rect 48179 16473 48188 16507
rect 48136 16464 48188 16473
rect 21824 16396 21876 16448
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 27620 16396 27672 16448
rect 28540 16396 28592 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 13268 16235 13320 16244
rect 13268 16201 13277 16235
rect 13277 16201 13311 16235
rect 13311 16201 13320 16235
rect 13268 16192 13320 16201
rect 11796 16167 11848 16176
rect 11796 16133 11805 16167
rect 11805 16133 11839 16167
rect 11839 16133 11848 16167
rect 11796 16124 11848 16133
rect 11336 16056 11388 16108
rect 15476 16192 15528 16244
rect 18696 16192 18748 16244
rect 46388 16192 46440 16244
rect 46756 16235 46808 16244
rect 46756 16201 46765 16235
rect 46765 16201 46799 16235
rect 46799 16201 46808 16235
rect 46756 16192 46808 16201
rect 15936 16124 15988 16176
rect 22100 16167 22152 16176
rect 22100 16133 22109 16167
rect 22109 16133 22143 16167
rect 22143 16133 22152 16167
rect 22100 16124 22152 16133
rect 22744 16124 22796 16176
rect 23388 16124 23440 16176
rect 14372 16099 14424 16108
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 16856 16056 16908 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 21824 16099 21876 16108
rect 21824 16065 21833 16099
rect 21833 16065 21867 16099
rect 21867 16065 21876 16099
rect 21824 16056 21876 16065
rect 27620 16124 27672 16176
rect 38200 16124 38252 16176
rect 13176 15988 13228 16040
rect 14096 15988 14148 16040
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15108 15988 15160 16040
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 20352 16031 20404 16040
rect 2964 15852 3016 15904
rect 20352 15997 20361 16031
rect 20361 15997 20395 16031
rect 20395 15997 20404 16031
rect 20352 15988 20404 15997
rect 21456 15988 21508 16040
rect 40684 16056 40736 16108
rect 47768 16099 47820 16108
rect 47768 16065 47777 16099
rect 47777 16065 47811 16099
rect 47811 16065 47820 16099
rect 47768 16056 47820 16065
rect 21088 15852 21140 15904
rect 22192 15852 22244 15904
rect 23572 15895 23624 15904
rect 23572 15861 23581 15895
rect 23581 15861 23615 15895
rect 23615 15861 23624 15895
rect 23572 15852 23624 15861
rect 24032 15852 24084 15904
rect 25504 15895 25556 15904
rect 25504 15861 25513 15895
rect 25513 15861 25547 15895
rect 25547 15861 25556 15895
rect 25504 15852 25556 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13360 15691 13412 15700
rect 13360 15657 13369 15691
rect 13369 15657 13403 15691
rect 13403 15657 13412 15691
rect 13360 15648 13412 15657
rect 15384 15648 15436 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 20352 15648 20404 15700
rect 46940 15648 46992 15700
rect 12256 15580 12308 15632
rect 15200 15580 15252 15632
rect 19524 15580 19576 15632
rect 14096 15555 14148 15564
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 16396 15512 16448 15564
rect 1768 15444 1820 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 13268 15308 13320 15360
rect 15476 15444 15528 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 20720 15512 20772 15564
rect 21732 15512 21784 15564
rect 21916 15512 21968 15564
rect 25504 15555 25556 15564
rect 25504 15521 25513 15555
rect 25513 15521 25547 15555
rect 25547 15521 25556 15555
rect 25504 15512 25556 15521
rect 27160 15555 27212 15564
rect 27160 15521 27169 15555
rect 27169 15521 27203 15555
rect 27203 15521 27212 15555
rect 27160 15512 27212 15521
rect 45560 15512 45612 15564
rect 21088 15487 21140 15496
rect 18420 15376 18472 15428
rect 14004 15308 14056 15360
rect 15384 15308 15436 15360
rect 16856 15308 16908 15360
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 22100 15487 22152 15496
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22100 15444 22152 15453
rect 21364 15376 21416 15428
rect 22192 15376 22244 15428
rect 24400 15444 24452 15496
rect 22008 15308 22060 15360
rect 22468 15351 22520 15360
rect 22468 15317 22477 15351
rect 22477 15317 22511 15351
rect 22511 15317 22520 15351
rect 22468 15308 22520 15317
rect 22652 15308 22704 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 14648 15104 14700 15156
rect 21732 15104 21784 15156
rect 22192 15104 22244 15156
rect 24400 15147 24452 15156
rect 24400 15113 24409 15147
rect 24409 15113 24443 15147
rect 24443 15113 24452 15147
rect 24400 15104 24452 15113
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 13912 15036 13964 15088
rect 13820 14968 13872 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 15200 15036 15252 15088
rect 18328 15011 18380 15020
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 14004 14943 14056 14952
rect 2780 14900 2832 14909
rect 14004 14909 14013 14943
rect 14013 14909 14047 14943
rect 14047 14909 14056 14943
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21364 14968 21416 15020
rect 21916 15036 21968 15088
rect 22468 15036 22520 15088
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22284 14968 22336 15020
rect 22652 15011 22704 15020
rect 22652 14977 22661 15011
rect 22661 14977 22695 15011
rect 22695 14977 22704 15011
rect 22652 14968 22704 14977
rect 24032 14968 24084 15020
rect 14004 14900 14056 14909
rect 18696 14900 18748 14952
rect 14924 14832 14976 14884
rect 18328 14832 18380 14884
rect 23572 14900 23624 14952
rect 13268 14764 13320 14816
rect 20904 14764 20956 14816
rect 22100 14764 22152 14816
rect 24400 14764 24452 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 24952 14560 25004 14612
rect 13820 14492 13872 14544
rect 13912 14424 13964 14476
rect 17776 14424 17828 14476
rect 21088 14492 21140 14544
rect 20904 14467 20956 14476
rect 20904 14433 20913 14467
rect 20913 14433 20947 14467
rect 20947 14433 20956 14467
rect 20904 14424 20956 14433
rect 2136 14356 2188 14365
rect 17040 14356 17092 14408
rect 17316 14331 17368 14340
rect 17316 14297 17325 14331
rect 17325 14297 17359 14331
rect 17359 14297 17368 14331
rect 17316 14288 17368 14297
rect 18328 14356 18380 14408
rect 20168 14356 20220 14408
rect 18696 14288 18748 14340
rect 21640 14356 21692 14408
rect 21364 14288 21416 14340
rect 17132 14220 17184 14272
rect 19984 14220 20036 14272
rect 20076 14220 20128 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 16764 13991 16816 14000
rect 16764 13957 16773 13991
rect 16773 13957 16807 13991
rect 16807 13957 16816 13991
rect 16764 13948 16816 13957
rect 17684 13948 17736 14000
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 20168 14059 20220 14068
rect 20168 14025 20177 14059
rect 20177 14025 20211 14059
rect 20211 14025 20220 14059
rect 20168 14016 20220 14025
rect 21824 14016 21876 14068
rect 18788 13991 18840 14000
rect 18788 13957 18797 13991
rect 18797 13957 18831 13991
rect 18831 13957 18840 13991
rect 18788 13948 18840 13957
rect 20904 13948 20956 14000
rect 15752 13880 15804 13932
rect 18696 13880 18748 13932
rect 20720 13923 20772 13932
rect 17316 13812 17368 13864
rect 3792 13676 3844 13728
rect 4804 13676 4856 13728
rect 16580 13676 16632 13728
rect 17224 13676 17276 13728
rect 17868 13744 17920 13796
rect 19340 13812 19392 13864
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 20996 13880 21048 13932
rect 27344 13880 27396 13932
rect 21640 13812 21692 13864
rect 20076 13787 20128 13796
rect 20076 13753 20085 13787
rect 20085 13753 20119 13787
rect 20119 13753 20128 13787
rect 20076 13744 20128 13753
rect 20720 13676 20772 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 21640 13472 21692 13524
rect 17776 13404 17828 13456
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 19432 13404 19484 13456
rect 19340 13379 19392 13388
rect 19340 13345 19349 13379
rect 19349 13345 19383 13379
rect 19383 13345 19392 13379
rect 19340 13336 19392 13345
rect 20720 13336 20772 13388
rect 14832 13200 14884 13252
rect 16672 13243 16724 13252
rect 16672 13209 16681 13243
rect 16681 13209 16715 13243
rect 16715 13209 16724 13243
rect 16672 13200 16724 13209
rect 18236 13200 18288 13252
rect 15384 13132 15436 13184
rect 17316 13132 17368 13184
rect 19984 13200 20036 13252
rect 21916 13200 21968 13252
rect 20904 13132 20956 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 14832 12928 14884 12980
rect 16396 12928 16448 12980
rect 17224 12928 17276 12980
rect 17776 12928 17828 12980
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 16764 12860 16816 12912
rect 17316 12860 17368 12912
rect 19340 12928 19392 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 15200 12792 15252 12844
rect 15844 12792 15896 12844
rect 16580 12724 16632 12776
rect 18236 12792 18288 12844
rect 19524 12860 19576 12912
rect 20168 12860 20220 12912
rect 20720 12792 20772 12844
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 16948 12588 17000 12640
rect 30012 12656 30064 12708
rect 47768 12631 47820 12640
rect 47768 12597 47777 12631
rect 47777 12597 47811 12631
rect 47811 12597 47820 12631
rect 47768 12588 47820 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 16672 12384 16724 12436
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 20168 12384 20220 12436
rect 15200 12180 15252 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17224 12180 17276 12232
rect 17868 12180 17920 12232
rect 20996 12248 21048 12300
rect 47768 12248 47820 12300
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 18236 12112 18288 12164
rect 20628 12180 20680 12232
rect 47676 12112 47728 12164
rect 15200 12044 15252 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 47676 11883 47728 11892
rect 47676 11849 47685 11883
rect 47685 11849 47719 11883
rect 47719 11849 47728 11883
rect 47676 11840 47728 11849
rect 15568 11772 15620 11824
rect 16948 11815 17000 11824
rect 16948 11781 16973 11815
rect 16973 11781 17000 11815
rect 16948 11772 17000 11781
rect 16580 11704 16632 11756
rect 25964 11704 26016 11756
rect 13820 11500 13872 11552
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 17776 11568 17828 11620
rect 17040 11500 17092 11552
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13268 11092 13320 11144
rect 15660 11296 15712 11348
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 16672 11160 16724 11212
rect 47768 11160 47820 11212
rect 14188 11024 14240 11076
rect 14096 10956 14148 11008
rect 15660 11092 15712 11144
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 19432 11024 19484 11076
rect 24860 11024 24912 11076
rect 25964 11024 26016 11076
rect 46480 11067 46532 11076
rect 46480 11033 46489 11067
rect 46489 11033 46523 11067
rect 46523 11033 46532 11067
rect 46480 11024 46532 11033
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 15568 10956 15620 11008
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 46480 10752 46532 10804
rect 2780 10684 2832 10736
rect 4896 10684 4948 10736
rect 14096 10727 14148 10736
rect 14096 10693 14105 10727
rect 14105 10693 14139 10727
rect 14139 10693 14148 10727
rect 14096 10684 14148 10693
rect 19432 10684 19484 10736
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 15200 10616 15252 10668
rect 16948 10616 17000 10668
rect 17684 10616 17736 10668
rect 23296 10616 23348 10668
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 17224 10548 17276 10600
rect 19432 10412 19484 10464
rect 46296 10455 46348 10464
rect 46296 10421 46305 10455
rect 46305 10421 46339 10455
rect 46339 10421 46348 10455
rect 46296 10412 46348 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 16672 10208 16724 10260
rect 16948 10140 17000 10192
rect 17868 10140 17920 10192
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 17224 10072 17276 10124
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 15568 9979 15620 9988
rect 15568 9945 15577 9979
rect 15577 9945 15611 9979
rect 15611 9945 15620 9979
rect 15568 9936 15620 9945
rect 17592 9936 17644 9988
rect 16580 9868 16632 9920
rect 17776 9936 17828 9988
rect 17868 9979 17920 9988
rect 17868 9945 17877 9979
rect 17877 9945 17911 9979
rect 17911 9945 17920 9979
rect 17868 9936 17920 9945
rect 47676 9936 47728 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17224 9664 17276 9716
rect 17868 9664 17920 9716
rect 19432 9664 19484 9716
rect 16580 9596 16632 9648
rect 18420 9596 18472 9648
rect 16856 9528 16908 9580
rect 19248 9528 19300 9580
rect 47676 9639 47728 9648
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 46204 9571 46256 9580
rect 46204 9537 46213 9571
rect 46213 9537 46247 9571
rect 46247 9537 46256 9571
rect 46204 9528 46256 9537
rect 47492 9528 47544 9580
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 29000 9460 29052 9512
rect 46480 9503 46532 9512
rect 46480 9469 46489 9503
rect 46489 9469 46523 9503
rect 46523 9469 46532 9503
rect 46480 9460 46532 9469
rect 15660 9392 15712 9444
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 17224 9324 17276 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 15568 9120 15620 9172
rect 19616 9120 19668 9172
rect 15200 8916 15252 8968
rect 16764 9052 16816 9104
rect 46388 9052 46440 9104
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 46480 9027 46532 9036
rect 46480 8993 46489 9027
rect 46489 8993 46523 9027
rect 46523 8993 46532 9027
rect 46480 8984 46532 8993
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 27160 8916 27212 8968
rect 28356 8916 28408 8968
rect 46296 8959 46348 8968
rect 46296 8925 46305 8959
rect 46305 8925 46339 8959
rect 46339 8925 46348 8959
rect 46296 8916 46348 8925
rect 16764 8891 16816 8900
rect 16764 8857 16773 8891
rect 16773 8857 16807 8891
rect 16807 8857 16816 8891
rect 16764 8848 16816 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 17224 8551 17276 8560
rect 3332 8304 3384 8356
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 17224 8517 17233 8551
rect 17233 8517 17267 8551
rect 17267 8517 17276 8551
rect 17224 8508 17276 8517
rect 47768 8551 47820 8560
rect 47768 8517 47777 8551
rect 47777 8517 47811 8551
rect 47811 8517 47820 8551
rect 47768 8508 47820 8517
rect 19248 8440 19300 8492
rect 17408 8372 17460 8424
rect 3148 8236 3200 8288
rect 17960 8304 18012 8356
rect 30104 8304 30156 8356
rect 17592 8236 17644 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 16764 8032 16816 8084
rect 17132 7964 17184 8016
rect 17960 7896 18012 7948
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 46020 7896 46072 7948
rect 48044 7939 48096 7948
rect 48044 7905 48053 7939
rect 48053 7905 48087 7939
rect 48087 7905 48096 7939
rect 48044 7896 48096 7905
rect 15200 7828 15252 7880
rect 16764 7828 16816 7880
rect 47492 7760 47544 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 3608 7488 3660 7540
rect 18052 7488 18104 7540
rect 1676 7420 1728 7472
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 45192 7327 45244 7336
rect 45192 7293 45201 7327
rect 45201 7293 45235 7327
rect 45235 7293 45244 7327
rect 45192 7284 45244 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 17408 6944 17460 6996
rect 3424 6808 3476 6860
rect 17960 6808 18012 6860
rect 47308 6851 47360 6860
rect 47308 6817 47317 6851
rect 47317 6817 47351 6851
rect 47351 6817 47360 6851
rect 47308 6808 47360 6817
rect 47492 6808 47544 6860
rect 16764 6740 16816 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 48136 6307 48188 6316
rect 48136 6273 48145 6307
rect 48145 6273 48179 6307
rect 48179 6273 48188 6307
rect 48136 6264 48188 6273
rect 47952 6103 48004 6112
rect 47952 6069 47961 6103
rect 47961 6069 47995 6103
rect 47995 6069 48004 6103
rect 47952 6060 48004 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 46848 5720 46900 5772
rect 21640 5652 21692 5704
rect 46572 5652 46624 5704
rect 22192 5516 22244 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 45836 5312 45888 5364
rect 46296 5312 46348 5364
rect 47952 5244 48004 5296
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 19984 5176 20036 5228
rect 20352 5176 20404 5228
rect 20996 5176 21048 5228
rect 22284 5176 22336 5228
rect 22100 5108 22152 5160
rect 46848 5176 46900 5228
rect 45192 5040 45244 5092
rect 18696 5015 18748 5024
rect 18696 4981 18705 5015
rect 18705 4981 18739 5015
rect 18739 4981 18748 5015
rect 18696 4972 18748 4981
rect 19616 5015 19668 5024
rect 19616 4981 19625 5015
rect 19625 4981 19659 5015
rect 19659 4981 19668 5015
rect 19616 4972 19668 4981
rect 20812 4972 20864 5024
rect 21548 4972 21600 5024
rect 22376 4972 22428 5024
rect 23020 4972 23072 5024
rect 27344 4972 27396 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 20352 4811 20404 4820
rect 20352 4777 20361 4811
rect 20361 4777 20395 4811
rect 20395 4777 20404 4811
rect 20352 4768 20404 4777
rect 20996 4811 21048 4820
rect 20996 4777 21005 4811
rect 21005 4777 21039 4811
rect 21039 4777 21048 4811
rect 20996 4768 21048 4777
rect 21640 4811 21692 4820
rect 21640 4777 21649 4811
rect 21649 4777 21683 4811
rect 21683 4777 21692 4811
rect 21640 4768 21692 4777
rect 22284 4811 22336 4820
rect 22284 4777 22293 4811
rect 22293 4777 22327 4811
rect 22327 4777 22336 4811
rect 22284 4768 22336 4777
rect 6920 4632 6972 4684
rect 9128 4564 9180 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 19340 4564 19392 4616
rect 19616 4564 19668 4616
rect 20812 4564 20864 4616
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 39856 4607 39908 4616
rect 15568 4496 15620 4548
rect 17132 4539 17184 4548
rect 17132 4505 17141 4539
rect 17141 4505 17175 4539
rect 17175 4505 17184 4539
rect 17132 4496 17184 4505
rect 39856 4573 39865 4607
rect 39865 4573 39899 4607
rect 39899 4573 39908 4607
rect 39856 4564 39908 4573
rect 46940 4700 46992 4752
rect 45836 4675 45888 4684
rect 45836 4641 45845 4675
rect 45845 4641 45879 4675
rect 45879 4641 45888 4675
rect 45836 4632 45888 4641
rect 47032 4675 47084 4684
rect 47032 4641 47041 4675
rect 47041 4641 47075 4675
rect 47075 4641 47084 4675
rect 47032 4632 47084 4641
rect 45192 4564 45244 4616
rect 46020 4539 46072 4548
rect 46020 4505 46029 4539
rect 46029 4505 46063 4539
rect 46063 4505 46072 4539
rect 46020 4496 46072 4505
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 20076 4428 20128 4480
rect 20812 4428 20864 4480
rect 22468 4428 22520 4480
rect 23572 4471 23624 4480
rect 23572 4437 23581 4471
rect 23581 4437 23615 4471
rect 23615 4437 23624 4471
rect 23572 4428 23624 4437
rect 39948 4471 40000 4480
rect 39948 4437 39957 4471
rect 39957 4437 39991 4471
rect 39991 4437 40000 4471
rect 39948 4428 40000 4437
rect 42800 4471 42852 4480
rect 42800 4437 42809 4471
rect 42809 4437 42843 4471
rect 42843 4437 42852 4471
rect 42800 4428 42852 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 18420 4224 18472 4276
rect 19984 4224 20036 4276
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 32956 4224 33008 4276
rect 39856 4224 39908 4276
rect 43076 4224 43128 4276
rect 45836 4224 45888 4276
rect 17500 4156 17552 4208
rect 21732 4156 21784 4208
rect 21824 4156 21876 4208
rect 22192 4156 22244 4208
rect 22376 4156 22428 4208
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 2872 4020 2924 4072
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 10140 4020 10192 4072
rect 3884 3952 3936 4004
rect 9036 3952 9088 4004
rect 17960 4088 18012 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 20076 4131 20128 4140
rect 17224 4020 17276 4072
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 22468 4088 22520 4140
rect 23848 4156 23900 4208
rect 24492 4156 24544 4208
rect 25136 4156 25188 4208
rect 22928 4088 22980 4140
rect 23388 4088 23440 4140
rect 19340 4020 19392 4072
rect 22100 4020 22152 4072
rect 25044 4088 25096 4140
rect 25412 4088 25464 4140
rect 32680 4156 32732 4208
rect 29184 4088 29236 4140
rect 33140 4131 33192 4140
rect 27620 4020 27672 4072
rect 29092 4020 29144 4072
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 30012 4020 30064 4072
rect 21824 3952 21876 4004
rect 8116 3884 8168 3936
rect 10876 3884 10928 3936
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14924 3884 14976 3936
rect 18236 3884 18288 3936
rect 18788 3884 18840 3936
rect 19248 3884 19300 3936
rect 20444 3884 20496 3936
rect 22008 3884 22060 3936
rect 24768 3884 24820 3936
rect 26976 3952 27028 4004
rect 31300 4063 31352 4072
rect 31300 4029 31309 4063
rect 31309 4029 31343 4063
rect 31343 4029 31352 4063
rect 31300 4020 31352 4029
rect 33140 4097 33149 4131
rect 33149 4097 33183 4131
rect 33183 4097 33192 4131
rect 33140 4088 33192 4097
rect 40040 4156 40092 4208
rect 46664 4199 46716 4208
rect 39212 4088 39264 4140
rect 39580 4088 39632 4140
rect 31668 4020 31720 4072
rect 40960 4088 41012 4140
rect 46664 4165 46673 4199
rect 46673 4165 46707 4199
rect 46707 4165 46716 4199
rect 46664 4156 46716 4165
rect 47768 4199 47820 4208
rect 47768 4165 47777 4199
rect 47777 4165 47811 4199
rect 47811 4165 47820 4199
rect 47768 4156 47820 4165
rect 41052 4063 41104 4072
rect 41052 4029 41061 4063
rect 41061 4029 41095 4063
rect 41095 4029 41104 4063
rect 41052 4020 41104 4029
rect 41328 4020 41380 4072
rect 41420 4020 41472 4072
rect 43076 4063 43128 4072
rect 43076 4029 43085 4063
rect 43085 4029 43119 4063
rect 43119 4029 43128 4063
rect 43076 4020 43128 4029
rect 43904 4020 43956 4072
rect 44088 4020 44140 4072
rect 45744 4088 45796 4140
rect 33140 3884 33192 3936
rect 39120 3884 39172 3936
rect 42432 3884 42484 3936
rect 42616 3927 42668 3936
rect 42616 3893 42625 3927
rect 42625 3893 42659 3927
rect 42659 3893 42668 3927
rect 42616 3884 42668 3893
rect 46480 3884 46532 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 3884 3680 3936 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 18144 3680 18196 3732
rect 19432 3680 19484 3732
rect 21272 3680 21324 3732
rect 3792 3612 3844 3664
rect 29920 3680 29972 3732
rect 39028 3680 39080 3732
rect 39212 3723 39264 3732
rect 39212 3689 39221 3723
rect 39221 3689 39255 3723
rect 39255 3689 39264 3723
rect 39212 3680 39264 3689
rect 42340 3680 42392 3732
rect 43444 3680 43496 3732
rect 44088 3680 44140 3732
rect 10876 3587 10928 3596
rect 1768 3476 1820 3528
rect 2136 3519 2188 3528
rect 2136 3485 2145 3519
rect 2145 3485 2179 3519
rect 2179 3485 2188 3519
rect 2136 3476 2188 3485
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 6460 3408 6512 3460
rect 7932 3408 7984 3460
rect 1952 3340 2004 3392
rect 7196 3340 7248 3392
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 10968 3544 11020 3596
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 13544 3476 13596 3528
rect 18696 3544 18748 3596
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 18236 3476 18288 3528
rect 15200 3408 15252 3460
rect 21916 3544 21968 3596
rect 22192 3544 22244 3596
rect 25596 3544 25648 3596
rect 27160 3587 27212 3596
rect 27160 3553 27169 3587
rect 27169 3553 27203 3587
rect 27203 3553 27212 3587
rect 27160 3544 27212 3553
rect 27344 3587 27396 3596
rect 27344 3553 27353 3587
rect 27353 3553 27387 3587
rect 27387 3553 27396 3587
rect 27620 3587 27672 3596
rect 27344 3544 27396 3553
rect 27620 3553 27629 3587
rect 27629 3553 27663 3587
rect 27663 3553 27672 3587
rect 27620 3544 27672 3553
rect 29000 3544 29052 3596
rect 30932 3544 30984 3596
rect 19340 3476 19392 3528
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 23020 3519 23072 3528
rect 20996 3408 21048 3460
rect 21088 3408 21140 3460
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 24584 3476 24636 3528
rect 33232 3587 33284 3596
rect 33232 3553 33241 3587
rect 33241 3553 33275 3587
rect 33275 3553 33284 3587
rect 42248 3612 42300 3664
rect 33232 3544 33284 3553
rect 35900 3519 35952 3528
rect 18420 3340 18472 3392
rect 18788 3340 18840 3392
rect 20904 3340 20956 3392
rect 22100 3340 22152 3392
rect 22192 3340 22244 3392
rect 22652 3408 22704 3460
rect 25228 3408 25280 3460
rect 25320 3408 25372 3460
rect 35900 3485 35909 3519
rect 35909 3485 35943 3519
rect 35943 3485 35952 3519
rect 35900 3476 35952 3485
rect 23296 3340 23348 3392
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 23848 3340 23900 3392
rect 35808 3408 35860 3460
rect 36176 3408 36228 3460
rect 29184 3340 29236 3392
rect 39856 3587 39908 3596
rect 39856 3553 39865 3587
rect 39865 3553 39899 3587
rect 39899 3553 39908 3587
rect 39856 3544 39908 3553
rect 40040 3544 40092 3596
rect 40224 3544 40276 3596
rect 40408 3544 40460 3596
rect 44732 3612 44784 3664
rect 47032 3612 47084 3664
rect 42616 3587 42668 3596
rect 42616 3553 42625 3587
rect 42625 3553 42659 3587
rect 42659 3553 42668 3587
rect 42616 3544 42668 3553
rect 42800 3587 42852 3596
rect 42800 3553 42809 3587
rect 42809 3553 42843 3587
rect 42843 3553 42852 3587
rect 42800 3544 42852 3553
rect 43168 3587 43220 3596
rect 43168 3553 43177 3587
rect 43177 3553 43211 3587
rect 43211 3553 43220 3587
rect 43168 3544 43220 3553
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 40132 3408 40184 3460
rect 41420 3408 41472 3460
rect 43444 3408 43496 3460
rect 47400 3408 47452 3460
rect 48964 3408 49016 3460
rect 43536 3340 43588 3392
rect 45376 3340 45428 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 17776 3136 17828 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 13728 3111 13780 3120
rect 13728 3077 13737 3111
rect 13737 3077 13771 3111
rect 13771 3077 13780 3111
rect 13728 3068 13780 3077
rect 17132 3068 17184 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 5908 3000 5960 3052
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 10692 3000 10744 3052
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 664 2932 716 2984
rect 7748 2932 7800 2984
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15200 2932 15252 2984
rect 8484 2864 8536 2916
rect 17684 2864 17736 2916
rect 18236 2975 18288 2984
rect 18236 2941 18245 2975
rect 18245 2941 18279 2975
rect 18279 2941 18288 2975
rect 18236 2932 18288 2941
rect 18420 3068 18472 3120
rect 19156 3068 19208 3120
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 23756 3136 23808 3188
rect 20812 3068 20864 3120
rect 20996 3111 21048 3120
rect 20996 3077 21005 3111
rect 21005 3077 21039 3111
rect 21039 3077 21048 3111
rect 20996 3068 21048 3077
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 22284 3068 22336 3120
rect 25780 3136 25832 3188
rect 28908 3136 28960 3188
rect 32772 3136 32824 3188
rect 36176 3179 36228 3188
rect 36176 3145 36185 3179
rect 36185 3145 36219 3179
rect 36219 3145 36228 3179
rect 36176 3136 36228 3145
rect 39580 3179 39632 3188
rect 39580 3145 39589 3179
rect 39589 3145 39623 3179
rect 39623 3145 39632 3179
rect 39580 3136 39632 3145
rect 24768 3111 24820 3120
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 24860 3068 24912 3120
rect 20076 3000 20128 3052
rect 20904 3043 20956 3052
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 31300 3000 31352 3052
rect 19892 2932 19944 2984
rect 19984 2932 20036 2984
rect 21088 2932 21140 2984
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 29092 2932 29144 2984
rect 32680 2932 32732 2984
rect 21456 2864 21508 2916
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 17408 2796 17460 2848
rect 22836 2864 22888 2916
rect 23020 2864 23072 2916
rect 32128 2864 32180 2916
rect 23204 2796 23256 2848
rect 25688 2796 25740 2848
rect 25780 2796 25832 2848
rect 32220 2796 32272 2848
rect 32956 3068 33008 3120
rect 33416 3068 33468 3120
rect 41420 3136 41472 3188
rect 43812 3136 43864 3188
rect 33048 3043 33100 3052
rect 33048 3009 33057 3043
rect 33057 3009 33091 3043
rect 33091 3009 33100 3043
rect 33048 3000 33100 3009
rect 36084 3000 36136 3052
rect 39672 3000 39724 3052
rect 33324 2932 33376 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 35900 2932 35952 2984
rect 41052 3068 41104 3120
rect 41328 3068 41380 3120
rect 48044 3136 48096 3188
rect 45376 3111 45428 3120
rect 39856 3000 39908 3052
rect 40132 3000 40184 3052
rect 40592 3000 40644 3052
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 39948 2932 40000 2984
rect 40224 2932 40276 2984
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 46756 3000 46808 3052
rect 47676 2932 47728 2984
rect 32864 2864 32916 2916
rect 40408 2796 40460 2848
rect 40500 2796 40552 2848
rect 45100 2796 45152 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 15200 2592 15252 2644
rect 18604 2635 18656 2644
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 18604 2592 18656 2601
rect 19340 2635 19392 2644
rect 19340 2601 19349 2635
rect 19349 2601 19383 2635
rect 19383 2601 19392 2635
rect 19340 2592 19392 2601
rect 20444 2592 20496 2644
rect 7104 2524 7156 2576
rect 7288 2456 7340 2508
rect 20720 2524 20772 2576
rect 23388 2592 23440 2644
rect 25044 2592 25096 2644
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 27620 2567 27672 2576
rect 27620 2533 27629 2567
rect 27629 2533 27663 2567
rect 27663 2533 27672 2567
rect 27620 2524 27672 2533
rect 32496 2524 32548 2576
rect 39304 2524 39356 2576
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 20260 2456 20312 2508
rect 26792 2456 26844 2508
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 2596 2388 2648 2440
rect 5172 2388 5224 2440
rect 8484 2388 8536 2440
rect 15476 2388 15528 2440
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 19156 2388 19208 2440
rect 23572 2388 23624 2440
rect 25688 2431 25740 2440
rect 25688 2397 25697 2431
rect 25697 2397 25731 2431
rect 25731 2397 25740 2431
rect 25688 2388 25740 2397
rect 27160 2388 27212 2440
rect 1308 2320 1360 2372
rect 7196 2320 7248 2372
rect 16120 2320 16172 2372
rect 20628 2320 20680 2372
rect 21916 2320 21968 2372
rect 24492 2320 24544 2372
rect 26424 2320 26476 2372
rect 27068 2320 27120 2372
rect 28356 2320 28408 2372
rect 29644 2388 29696 2440
rect 47032 2456 47084 2508
rect 35440 2388 35492 2440
rect 35808 2431 35860 2440
rect 35808 2397 35817 2431
rect 35817 2397 35851 2431
rect 35851 2397 35860 2431
rect 35808 2388 35860 2397
rect 41236 2388 41288 2440
rect 41328 2431 41380 2440
rect 41328 2397 41337 2431
rect 41337 2397 41371 2431
rect 41371 2397 41380 2431
rect 41328 2388 41380 2397
rect 43812 2388 43864 2440
rect 43904 2431 43956 2440
rect 43904 2397 43913 2431
rect 43913 2397 43947 2431
rect 43947 2397 43956 2431
rect 43904 2388 43956 2397
rect 46020 2388 46072 2440
rect 38016 2320 38068 2372
rect 39304 2320 39356 2372
rect 40960 2320 41012 2372
rect 46388 2320 46440 2372
rect 48320 2320 48372 2372
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 23480 2252 23532 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 9128 1980 9180 2032
rect 23940 1980 23992 2032
rect 2136 1912 2188 1964
rect 24676 1912 24728 1964
rect 2872 1844 2924 1896
rect 21180 1844 21232 1896
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49314 2034 50000
rect 1922 49286 2176 49314
rect 1922 49200 2034 49286
rect 32 17338 60 49200
rect 1858 47696 1914 47705
rect 1858 47631 1914 47640
rect 1872 46646 1900 47631
rect 2148 47054 2176 49286
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 2608 47138 2636 49200
rect 2608 47110 2820 47138
rect 2792 47054 2820 47110
rect 3252 47054 3280 49200
rect 2136 47048 2188 47054
rect 2136 46990 2188 46996
rect 2780 47048 2832 47054
rect 2780 46990 2832 46996
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3422 47016 3478 47025
rect 2504 46980 2556 46986
rect 3422 46951 3478 46960
rect 2504 46922 2556 46928
rect 1860 46640 1912 46646
rect 1860 46582 1912 46588
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1872 42945 1900 43250
rect 1952 43104 2004 43110
rect 1952 43046 2004 43052
rect 1858 42936 1914 42945
rect 1858 42871 1914 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1584 41540 1636 41546
rect 1858 41511 1914 41520
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 35698 1440 36110
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1596 35086 1624 35391
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 34886
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1400 32836 1452 32842
rect 1400 32778 1452 32784
rect 1412 32026 1440 32778
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 1596 31822 1624 32671
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 20 17332 72 17338
rect 20 17274 72 17280
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1688 7478 1716 25162
rect 1780 19990 1808 32302
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1964 20505 1992 43046
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 2044 33448 2096 33454
rect 2044 33390 2096 33396
rect 2056 32502 2084 33390
rect 2044 32496 2096 32502
rect 2044 32438 2096 32444
rect 2044 31816 2096 31822
rect 2044 31758 2096 31764
rect 2056 31346 2084 31758
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1950 20496 2006 20505
rect 1950 20431 2006 20440
rect 1768 19984 1820 19990
rect 1768 19926 1820 19932
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1872 17785 1900 18226
rect 2148 17814 2176 41074
rect 2412 40452 2464 40458
rect 2412 40394 2464 40400
rect 2228 36100 2280 36106
rect 2228 36042 2280 36048
rect 2240 35290 2268 36042
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2320 35080 2372 35086
rect 2320 35022 2372 35028
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2332 18766 2360 35022
rect 2424 29306 2452 40394
rect 2412 29300 2464 29306
rect 2412 29242 2464 29248
rect 2516 22098 2544 46922
rect 3148 46912 3200 46918
rect 3148 46854 3200 46860
rect 3160 46646 3188 46854
rect 3148 46640 3200 46646
rect 3148 46582 3200 46588
rect 2596 46368 2648 46374
rect 2596 46310 2648 46316
rect 2872 46368 2924 46374
rect 2872 46310 2924 46316
rect 3054 46336 3110 46345
rect 2608 26586 2636 46310
rect 2884 45422 2912 46310
rect 3054 46271 3110 46280
rect 2964 45824 3016 45830
rect 2964 45766 3016 45772
rect 2976 45558 3004 45766
rect 2964 45552 3016 45558
rect 2964 45494 3016 45500
rect 3068 45422 3096 46271
rect 2872 45416 2924 45422
rect 2872 45358 2924 45364
rect 3056 45416 3108 45422
rect 3056 45358 3108 45364
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36242 2820 36751
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 3240 32836 3292 32842
rect 3240 32778 3292 32784
rect 3252 32366 3280 32778
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2792 31278 2820 31991
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2872 31680 2924 31686
rect 2872 31622 2924 31628
rect 2884 31414 2912 31622
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2596 26580 2648 26586
rect 2596 26522 2648 26528
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2136 17808 2188 17814
rect 1858 17776 1914 17785
rect 2136 17750 2188 17756
rect 1858 17711 1914 17720
rect 2148 17678 2176 17750
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17270 1992 17478
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2056 16794 2084 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2792 16425 2820 17070
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2976 15910 3004 31758
rect 3252 19961 3280 32302
rect 3238 19952 3294 19961
rect 3238 19887 3294 19896
rect 3436 19242 3464 46951
rect 3896 46594 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 5828 47054 5856 49200
rect 7116 47054 7144 49200
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 3896 46566 4016 46594
rect 3988 46510 4016 46566
rect 3884 46504 3936 46510
rect 3884 46446 3936 46452
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3896 46170 3924 46446
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3514 44976 3570 44985
rect 3514 44911 3570 44920
rect 3528 21078 3556 44911
rect 3698 43616 3754 43625
rect 3698 43551 3754 43560
rect 3606 39536 3662 39545
rect 3606 39471 3662 39480
rect 3620 21418 3648 39471
rect 3712 24614 3740 43551
rect 3790 31376 3846 31385
rect 3790 31311 3846 31320
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3608 21412 3660 21418
rect 3608 21354 3660 21360
rect 3516 21072 3568 21078
rect 3516 21014 3568 21020
rect 3804 20602 3832 31311
rect 3974 28656 4030 28665
rect 3974 28591 4030 28600
rect 3988 27946 4016 28591
rect 3976 27940 4028 27946
rect 3976 27882 4028 27888
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3988 19718 4016 19751
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3988 17746 4016 18391
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3974 17096 4030 17105
rect 3974 17031 4030 17040
rect 3988 16998 4016 17031
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 2778 15056 2834 15065
rect 1768 15020 1820 15026
rect 2778 14991 2834 15000
rect 1768 14962 1820 14968
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 2148 3534 2176 14350
rect 3792 13728 3844 13734
rect 3790 13696 3792 13705
rect 3844 13696 3846 13705
rect 3790 13631 3846 13640
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2792 10305 2820 10678
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7585 3188 8230
rect 3146 7576 3202 7585
rect 3146 7511 3202 7520
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2884 3738 2912 4014
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1780 3058 1808 3470
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3126 1992 3334
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 800 1348 2314
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1970 2176 2246
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 2608 800 2636 2382
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 1902 2912 2246
rect 2872 1896 2924 1902
rect 2872 1838 2924 1844
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2976 785 3004 4014
rect 3344 1465 3372 8298
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3422 6896 3478 6905
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3424 6802 3476 6808
rect 3620 3505 3648 7482
rect 4080 6914 4108 46922
rect 4620 46436 4672 46442
rect 4620 46378 4672 46384
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46170 4660 46378
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4816 13734 4844 24618
rect 5000 20262 5028 46922
rect 6920 46912 6972 46918
rect 6920 46854 6972 46860
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4908 10742 4936 18090
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3988 6886 4108 6914
rect 3988 4049 4016 6886
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6932 4690 6960 46854
rect 7852 35494 7880 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 8312 45526 8432 45554
rect 8312 35894 8340 45526
rect 8312 35866 8432 35894
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 8404 27538 8432 35866
rect 9508 35562 9536 46922
rect 10980 46374 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 12912 47054 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49450 15558 50000
rect 15304 49422 15558 49450
rect 13740 47122 13860 47138
rect 13740 47116 13872 47122
rect 13740 47110 13820 47116
rect 13820 47058 13872 47064
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 11704 46980 11756 46986
rect 11704 46922 11756 46928
rect 12440 46980 12492 46986
rect 12440 46922 12492 46928
rect 11244 46436 11296 46442
rect 11244 46378 11296 46384
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 11256 46170 11284 46378
rect 11244 46164 11296 46170
rect 11244 46106 11296 46112
rect 9496 35556 9548 35562
rect 9496 35498 9548 35504
rect 11716 31686 11744 46922
rect 12452 36310 12480 46922
rect 14200 46510 14228 49200
rect 14372 47048 14424 47054
rect 14372 46990 14424 46996
rect 13820 46504 13872 46510
rect 13820 46446 13872 46452
rect 14004 46504 14056 46510
rect 14004 46446 14056 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 13832 46170 13860 46446
rect 13820 46164 13872 46170
rect 13820 46106 13872 46112
rect 14016 45626 14044 46446
rect 14004 45620 14056 45626
rect 14004 45562 14056 45568
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 13740 45354 13768 45426
rect 13728 45348 13780 45354
rect 13728 45290 13780 45296
rect 12440 36304 12492 36310
rect 12440 36246 12492 36252
rect 13740 31754 13768 45290
rect 14384 32298 14412 46990
rect 15304 46918 15332 49422
rect 15446 49200 15558 49422
rect 16090 49314 16202 50000
rect 16090 49286 16528 49314
rect 16090 49200 16202 49286
rect 16500 47054 16528 49286
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26712 49286 27150 49314
rect 16488 47048 16540 47054
rect 16488 46990 16540 46996
rect 15844 46980 15896 46986
rect 15844 46922 15896 46928
rect 15292 46912 15344 46918
rect 15292 46854 15344 46860
rect 15856 35630 15884 46922
rect 16488 46912 16540 46918
rect 16488 46854 16540 46860
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 14740 35080 14792 35086
rect 14740 35022 14792 35028
rect 14372 32292 14424 32298
rect 14372 32234 14424 32240
rect 14752 31890 14780 35022
rect 15016 35012 15068 35018
rect 15016 34954 15068 34960
rect 15028 34678 15056 34954
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 15856 34610 15884 35566
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 15844 34604 15896 34610
rect 15844 34546 15896 34552
rect 16120 34604 16172 34610
rect 16120 34546 16172 34552
rect 15200 32768 15252 32774
rect 15200 32710 15252 32716
rect 15212 31890 15240 32710
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15672 31754 15700 32166
rect 13648 31726 13768 31754
rect 15660 31748 15712 31754
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 8588 27674 8616 27950
rect 8576 27668 8628 27674
rect 8576 27610 8628 27616
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8220 26994 8248 27406
rect 9128 27396 9180 27402
rect 9128 27338 9180 27344
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 9140 27130 9168 27338
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8220 26466 8248 26930
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8128 26438 8248 26466
rect 8956 26450 8984 26726
rect 8944 26444 8996 26450
rect 8128 24206 8156 26438
rect 8944 26386 8996 26392
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8496 25906 8524 26182
rect 9232 26042 9260 26250
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8496 24886 8524 25842
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8588 25294 8616 25774
rect 9692 25362 9720 27270
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 9956 26308 10008 26314
rect 9956 26250 10008 26256
rect 9968 26042 9996 26250
rect 9956 26036 10008 26042
rect 9956 25978 10008 25984
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9220 25152 9272 25158
rect 9220 25094 9272 25100
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8220 24410 8248 24686
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8208 24404 8260 24410
rect 8208 24346 8260 24352
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8496 20482 8524 20878
rect 7852 20466 8524 20482
rect 7840 20460 8524 20466
rect 7892 20454 8524 20460
rect 7840 20402 7892 20408
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18358 7604 18702
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 8496 17678 8524 20454
rect 8588 20398 8616 24550
rect 8956 24274 8984 24550
rect 9232 24274 9260 25094
rect 9600 24274 9628 25230
rect 9692 24410 9720 25298
rect 10060 25294 10088 25842
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9600 23730 9628 24210
rect 9968 24138 9996 25094
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9956 23724 10008 23730
rect 10060 23712 10088 25230
rect 10244 24818 10272 26930
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 25430 10640 25842
rect 11532 25498 11560 26862
rect 11808 26586 11836 26862
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 11624 26042 11652 26386
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11808 26042 11836 26182
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11704 25968 11756 25974
rect 11704 25910 11756 25916
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 10600 25424 10652 25430
rect 10600 25366 10652 25372
rect 10612 25294 10640 25366
rect 11716 25362 11744 25910
rect 11808 25906 11836 25978
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 12452 25498 12480 26998
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25906 12572 26182
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12636 25838 12664 26318
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12532 25424 12584 25430
rect 12532 25366 12584 25372
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11348 24818 11376 25230
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11716 24410 11744 25298
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 10008 23684 10088 23712
rect 9956 23666 10008 23672
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9784 23186 9812 23462
rect 9968 23322 9996 23666
rect 10796 23662 10824 24142
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 11256 23594 11284 24006
rect 11716 23798 11744 24142
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11808 23730 11836 24006
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9508 22778 9536 23054
rect 10060 23050 10088 23462
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 11256 22982 11284 23530
rect 11808 23526 11836 23666
rect 12084 23526 12112 24210
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12360 23322 12388 25230
rect 12544 24818 12572 25366
rect 12728 25362 12756 27270
rect 13372 26858 13400 27338
rect 13464 27334 13492 28086
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13556 27334 13584 28018
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13004 25838 13032 26318
rect 13188 25906 13216 26726
rect 13372 26450 13400 26794
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13004 25430 13032 25774
rect 13188 25770 13216 25842
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12544 23798 12572 24754
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12636 24274 12664 24550
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12360 22982 12388 23258
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9692 21486 9720 22578
rect 11256 22098 11284 22918
rect 12636 22642 12664 23598
rect 12728 23526 12756 25298
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12820 23662 12848 24754
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23798 13492 24006
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 12636 22030 12664 22578
rect 12728 22522 12756 23462
rect 13188 23322 13216 23598
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12728 22506 12848 22522
rect 12728 22500 12860 22506
rect 12728 22494 12808 22500
rect 12808 22442 12860 22448
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 11072 21690 11100 21898
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9048 21146 9076 21422
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9692 20942 9720 21422
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 21010 10272 21286
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 9692 19786 9720 20742
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 10888 19514 10916 19790
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 11072 19378 11100 21490
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11624 20942 11652 21286
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11716 20330 11744 21490
rect 11992 21146 12020 21558
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11992 20534 12020 21082
rect 12176 21010 12204 21286
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 11980 20528 12032 20534
rect 12164 20528 12216 20534
rect 12032 20476 12164 20482
rect 11980 20470 12216 20476
rect 11796 20460 11848 20466
rect 11992 20454 12204 20470
rect 11796 20402 11848 20408
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11256 19922 11284 20266
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11256 19446 11284 19858
rect 11808 19718 11836 20402
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11900 19854 11928 20334
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11992 19854 12020 19994
rect 12176 19922 12204 20198
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11900 19514 11928 19790
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11072 18766 11100 19314
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11808 18698 11836 19110
rect 11900 18970 11928 19314
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8588 17678 8616 18158
rect 8772 17814 8800 18158
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8128 16794 8156 17070
rect 8496 17066 8524 17614
rect 9048 17134 9076 17682
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9968 17338 9996 17614
rect 11256 17610 11284 18566
rect 11808 18222 11836 18634
rect 11900 18290 11928 18906
rect 11992 18834 12020 19654
rect 12176 19310 12204 19722
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12176 18970 12204 19246
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11992 18290 12020 18770
rect 12268 18766 12296 19654
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 10520 17490 10548 17546
rect 11900 17542 11928 18226
rect 11888 17536 11940 17542
rect 10520 17462 10640 17490
rect 11888 17478 11940 17484
rect 10612 17354 10640 17462
rect 10612 17338 10732 17354
rect 9956 17332 10008 17338
rect 10612 17332 10744 17338
rect 10612 17326 10692 17332
rect 9956 17274 10008 17280
rect 10692 17274 10744 17280
rect 11992 17134 12020 18226
rect 12360 18154 12388 19314
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17202 12388 17614
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 3974 4040 4030 4049
rect 3884 4004 3936 4010
rect 3974 3975 4030 3984
rect 3884 3946 3936 3952
rect 3896 3738 3924 3946
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3606 3496 3662 3505
rect 3606 3431 3662 3440
rect 3804 1850 3832 3606
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 3058 5948 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 3804 1822 3924 1850
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3896 800 3924 1822
rect 5184 800 5212 2382
rect 6472 800 6500 3402
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 800 7144 2518
rect 7208 2378 7236 3334
rect 7944 3058 7972 3402
rect 8128 3126 8156 3878
rect 8220 3534 8248 16594
rect 11992 16590 12020 17070
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11348 16114 11376 16458
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 12268 15638 12296 16526
rect 12360 16522 12388 17138
rect 12452 16590 12480 17206
rect 12544 17134 12572 18294
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17882 12664 18158
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12728 16998 12756 21898
rect 12820 21554 12848 22442
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 21622 13032 22374
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12912 20942 12940 21354
rect 13004 21146 13032 21422
rect 13096 21350 13124 23054
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 13648 20874 13676 31726
rect 15660 31690 15712 31696
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13740 27062 13768 27270
rect 14200 27130 14228 28086
rect 14292 28082 14320 31078
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 15304 29034 15332 29514
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14280 28076 14332 28082
rect 14332 28036 14412 28064
rect 14280 28018 14332 28024
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13740 26790 13768 26862
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13740 20602 13768 26726
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14108 26246 14136 26386
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13832 25838 13860 25978
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 14108 25770 14136 26182
rect 14200 26042 14228 27066
rect 14384 27062 14412 28036
rect 14476 27130 14504 28086
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 14096 25764 14148 25770
rect 14096 25706 14148 25712
rect 14384 25498 14412 26318
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14384 24886 14412 25230
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14004 23792 14056 23798
rect 14004 23734 14056 23740
rect 13912 22976 13964 22982
rect 13912 22918 13964 22924
rect 13924 22642 13952 22918
rect 14016 22778 14044 23734
rect 14108 23662 14136 24754
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13924 20602 13952 21558
rect 14108 20942 14136 23598
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18358 12940 19110
rect 13648 18970 13676 20470
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13832 19718 13860 20402
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18358 13492 18566
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 13648 16794 13676 18906
rect 13912 18692 13964 18698
rect 13912 18634 13964 18640
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16046 13216 16390
rect 13280 16250 13308 16526
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13372 15706 13400 16390
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 14822 13308 15302
rect 13832 15026 13860 18566
rect 13924 15094 13952 18634
rect 14108 17678 14136 20878
rect 14568 18698 14596 27882
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 15028 27674 15056 27814
rect 15120 27674 15148 27882
rect 15016 27668 15068 27674
rect 15016 27610 15068 27616
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14660 27130 14688 27406
rect 15200 27396 15252 27402
rect 15252 27356 15332 27384
rect 15200 27338 15252 27344
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 15304 27062 15332 27356
rect 15292 27056 15344 27062
rect 15292 26998 15344 27004
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14660 26042 14688 26250
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14752 25922 14780 26930
rect 14660 25894 14780 25922
rect 14924 25900 14976 25906
rect 14660 22094 14688 25894
rect 14924 25842 14976 25848
rect 14936 25362 14964 25842
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 15396 25294 15424 26930
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15764 26042 15792 26318
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14752 23866 14780 24278
rect 15212 24274 15240 24550
rect 15200 24268 15252 24274
rect 15200 24210 15252 24216
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14844 23730 14872 24142
rect 14936 23866 14964 24142
rect 15672 23866 15700 25842
rect 15856 24614 15884 34546
rect 16132 34406 16160 34546
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16132 33998 16160 34342
rect 16408 34202 16436 34954
rect 16396 34196 16448 34202
rect 16396 34138 16448 34144
rect 16120 33992 16172 33998
rect 16120 33934 16172 33940
rect 15936 33040 15988 33046
rect 15936 32982 15988 32988
rect 15948 32434 15976 32982
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15948 31890 15976 32370
rect 16132 32298 16160 33934
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 16132 30734 16160 32234
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 16132 30258 16160 30670
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29578 15976 29990
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 16040 29170 16068 29650
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 16040 28626 16068 29106
rect 16028 28620 16080 28626
rect 16028 28562 16080 28568
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16224 26518 16252 27406
rect 16212 26512 16264 26518
rect 16212 26454 16264 26460
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15752 24132 15804 24138
rect 15752 24074 15804 24080
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14844 23118 14872 23666
rect 15672 23254 15700 23802
rect 15764 23322 15792 24074
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 14660 22066 14780 22094
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14660 21486 14688 21966
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14752 18630 14780 22066
rect 14844 20466 14872 23054
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 15028 22098 15056 22374
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15672 21554 15700 23054
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14844 19854 14872 20402
rect 15304 20058 15332 20538
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14844 18766 14872 19790
rect 15304 18970 15332 19790
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15580 19242 15608 19722
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 19378 15792 19654
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17202 14320 17478
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16114 14412 16934
rect 14476 16658 14504 17682
rect 15488 17202 15516 18566
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16658 14688 16934
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14108 15570 14136 15982
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 13394 13308 14758
rect 13832 14550 13860 14962
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13924 14482 13952 15030
rect 14016 14958 14044 15302
rect 14108 15026 14136 15506
rect 14660 15162 14688 15982
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14936 14890 14964 16594
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16046 15148 16390
rect 15488 16250 15516 17138
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 16522 15700 16934
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15502 15148 15982
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15212 15094 15240 15574
rect 15396 15366 15424 15642
rect 15488 15502 15516 16186
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13280 11150 13308 13330
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12986 14136 13262
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14844 12986 14872 13194
rect 15396 13190 15424 15302
rect 15764 13938 15792 18702
rect 15856 18272 15884 22578
rect 16500 22030 16528 46854
rect 17420 45554 17448 49200
rect 18708 47054 18736 49200
rect 19340 47184 19392 47190
rect 19340 47126 19392 47132
rect 18696 47048 18748 47054
rect 18696 46990 18748 46996
rect 17420 45526 17540 45554
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 17144 34542 17172 34886
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 16684 32570 16712 32846
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16670 32464 16726 32473
rect 16670 32399 16672 32408
rect 16724 32399 16726 32408
rect 16672 32370 16724 32376
rect 16868 32298 16896 32778
rect 16856 32292 16908 32298
rect 16856 32234 16908 32240
rect 16868 31958 16896 32234
rect 16856 31952 16908 31958
rect 16856 31894 16908 31900
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16592 31414 16620 31622
rect 16960 31482 16988 32846
rect 17408 32496 17460 32502
rect 17406 32464 17408 32473
rect 17460 32464 17462 32473
rect 17316 32428 17368 32434
rect 17406 32399 17462 32408
rect 17316 32370 17368 32376
rect 16948 31476 17000 31482
rect 16948 31418 17000 31424
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 17040 30660 17092 30666
rect 17040 30602 17092 30608
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 28490 16620 30534
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16776 29850 16804 30194
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 17052 28694 17080 30602
rect 17328 30122 17356 32370
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17316 30116 17368 30122
rect 17316 30058 17368 30064
rect 17328 29578 17356 30058
rect 17420 29714 17448 30534
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17512 29594 17540 45526
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 17684 35012 17736 35018
rect 17684 34954 17736 34960
rect 17696 34746 17724 34954
rect 17684 34740 17736 34746
rect 17684 34682 17736 34688
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 17960 34468 18012 34474
rect 17960 34410 18012 34416
rect 17776 33448 17828 33454
rect 17776 33390 17828 33396
rect 17684 33312 17736 33318
rect 17684 33254 17736 33260
rect 17696 33114 17724 33254
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17788 32026 17816 33390
rect 17972 32978 18000 34410
rect 18064 33658 18092 34614
rect 18156 34542 18184 35430
rect 19064 35216 19116 35222
rect 19064 35158 19116 35164
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18144 34536 18196 34542
rect 18144 34478 18196 34484
rect 18984 33658 19012 34546
rect 19076 34542 19104 35158
rect 19260 35154 19288 37198
rect 19352 36258 19380 47126
rect 19432 47048 19484 47054
rect 19432 46990 19484 46996
rect 19444 46578 19472 46990
rect 19996 46918 20024 49200
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19432 46572 19484 46578
rect 19432 46514 19484 46520
rect 20640 46510 20668 49200
rect 20904 47048 20956 47054
rect 20904 46990 20956 46996
rect 20168 46504 20220 46510
rect 20168 46446 20220 46452
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 20180 46170 20208 46446
rect 20168 46164 20220 46170
rect 20168 46106 20220 46112
rect 20916 46034 20944 46990
rect 21284 46034 21312 49200
rect 22100 47116 22152 47122
rect 22100 47058 22152 47064
rect 21824 46912 21876 46918
rect 21824 46854 21876 46860
rect 20904 46028 20956 46034
rect 20904 45970 20956 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 20076 45960 20128 45966
rect 20076 45902 20128 45908
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 20088 45422 20116 45902
rect 20720 45892 20772 45898
rect 20720 45834 20772 45840
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 20732 45558 20760 45834
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 20720 45552 20772 45558
rect 20720 45494 20772 45500
rect 20076 45416 20128 45422
rect 20076 45358 20128 45364
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19432 37868 19484 37874
rect 19432 37810 19484 37816
rect 19444 36378 19472 37810
rect 19524 37664 19576 37670
rect 19524 37606 19576 37612
rect 19536 37330 19564 37606
rect 19524 37324 19576 37330
rect 19524 37266 19576 37272
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19352 36230 19472 36258
rect 19248 35148 19300 35154
rect 19248 35090 19300 35096
rect 19064 34536 19116 34542
rect 19064 34478 19116 34484
rect 19260 34218 19288 35090
rect 19260 34190 19380 34218
rect 19352 34066 19380 34190
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 18972 33652 19024 33658
rect 18972 33594 19024 33600
rect 19338 33552 19394 33561
rect 19306 33496 19338 33504
rect 19306 33487 19394 33496
rect 19306 33476 19380 33487
rect 19306 33446 19334 33476
rect 19294 33440 19346 33446
rect 19294 33382 19346 33388
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18064 32434 18092 32846
rect 18248 32434 18276 32914
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18616 32570 18644 32846
rect 18696 32768 18748 32774
rect 18696 32710 18748 32716
rect 18604 32564 18656 32570
rect 18604 32506 18656 32512
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18616 32298 18644 32506
rect 18604 32292 18656 32298
rect 18604 32234 18656 32240
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 17788 30802 17816 31962
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 17776 30796 17828 30802
rect 17776 30738 17828 30744
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17604 30394 17632 30670
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17788 30394 17816 30602
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17776 30388 17828 30394
rect 17776 30330 17828 30336
rect 17776 30184 17828 30190
rect 17776 30126 17828 30132
rect 17788 29714 17816 30126
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 17880 29646 17908 29990
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 17420 29566 17540 29594
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 17236 29238 17264 29446
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 17040 28688 17092 28694
rect 17040 28630 17092 28636
rect 16580 28484 16632 28490
rect 16580 28426 16632 28432
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 16684 26518 16712 27338
rect 17144 27130 17172 27338
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16672 26512 16724 26518
rect 16672 26454 16724 26460
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16592 25906 16620 26318
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16592 25362 16620 25842
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16868 25498 16896 25774
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16856 25288 16908 25294
rect 16960 25276 16988 26930
rect 16908 25248 16988 25276
rect 16856 25230 16908 25236
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16776 23866 16804 24686
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16868 23594 16896 25230
rect 17420 24274 17448 29566
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16960 23118 16988 23666
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22642 16712 22918
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16868 20534 16896 20742
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19378 15976 20198
rect 16592 19718 16620 20334
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 20058 17172 20198
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16684 19514 16712 19790
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18902 16068 19246
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 15936 18284 15988 18290
rect 15856 18244 15936 18272
rect 15936 18226 15988 18232
rect 15948 17882 15976 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15948 17066 15976 17818
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15948 15706 15976 16118
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16408 15570 16436 16594
rect 16868 16114 16896 17138
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16658 17080 16934
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12238 15240 12786
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13832 10674 13860 11494
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10742 14136 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14200 8498 14228 11018
rect 15212 10674 15240 12038
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15396 10130 15424 13126
rect 15856 12850 15884 15438
rect 16868 15366 16896 16050
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12986 16436 13262
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 16592 12782 16620 13670
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15580 11014 15608 11766
rect 16592 11762 16620 12718
rect 16684 12442 16712 13194
rect 16776 12918 16804 13942
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16672 12436 16724 12442
rect 16868 12434 16896 15302
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16672 12378 16724 12384
rect 16776 12406 16896 12434
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15672 11150 15700 11290
rect 16040 11218 16068 11494
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10810 15608 10950
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15580 9178 15608 9930
rect 15672 9450 15700 11086
rect 16684 10266 16712 11154
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9654 16620 9862
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 16592 9042 16620 9590
rect 16776 9110 16804 12406
rect 16960 12238 16988 12582
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16960 10674 16988 11766
rect 17052 11558 17080 14350
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 14074 17172 14214
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17328 13870 17356 14282
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17328 13682 17356 13806
rect 17236 12986 17264 13670
rect 17328 13654 17448 13682
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17236 12434 17264 12922
rect 17328 12918 17356 13126
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17144 12406 17264 12434
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16960 10198 16988 10610
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 15212 7886 15240 8910
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16776 8090 16804 8842
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 7970 16896 9522
rect 16960 9382 16988 10134
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17144 8022 17172 12406
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 10606 17264 12174
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10130 17264 10542
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9722 17264 10066
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 8566 17264 9318
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17328 8378 17356 12854
rect 17420 8430 17448 13654
rect 17236 8350 17356 8378
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 16776 7942 16896 7970
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 16776 7886 16804 7942
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4146 9168 4558
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7300 2514 7328 2790
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7760 800 7788 2926
rect 8496 2922 8524 4082
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8496 1306 8524 2382
rect 8404 1278 8524 1306
rect 8404 800 8432 1278
rect 9048 800 9076 3946
rect 10152 3738 10180 4014
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10888 3602 10916 3878
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10704 3058 10732 3470
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 2038 9168 2246
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 10980 800 11008 3538
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 3058 13584 3470
rect 13740 3126 13768 3878
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14200 800 14228 2926
rect 14936 1578 14964 3878
rect 15212 3466 15240 7822
rect 16776 6798 16804 7822
rect 17236 7410 17264 8350
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 7002 17448 7278
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2650 15240 2926
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15580 2514 15608 4490
rect 17144 3126 17172 4490
rect 17512 4214 17540 29446
rect 17696 28762 17724 29446
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 17972 28082 18000 31894
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 18064 28150 18092 31758
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 18340 31346 18368 31690
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18156 30258 18184 30670
rect 18248 30274 18276 31282
rect 18432 30666 18460 32166
rect 18708 31958 18736 32710
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 18696 31952 18748 31958
rect 18696 31894 18748 31900
rect 19076 31822 19104 32370
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19352 32026 19380 32302
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19352 30938 19380 31690
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 18432 30326 18460 30602
rect 18420 30320 18472 30326
rect 18248 30258 18368 30274
rect 18420 30262 18472 30268
rect 18144 30252 18196 30258
rect 18248 30252 18380 30258
rect 18248 30246 18328 30252
rect 18144 30194 18196 30200
rect 18328 30194 18380 30200
rect 18340 30054 18368 30194
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19168 28966 19196 29990
rect 19352 29238 19380 29990
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19352 28558 19380 29174
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17972 25294 18000 28018
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18708 27130 18736 27338
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18892 27062 18920 27270
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 19352 26790 19380 28494
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19352 25838 19380 26726
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23730 17632 24210
rect 17788 23866 17816 24686
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17880 23730 17908 25162
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24886 18092 25094
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 24206 18184 24550
rect 18340 24206 18368 25230
rect 18524 24614 18552 25230
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17972 23730 18000 24074
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 18156 23526 18184 24142
rect 18340 23866 18368 24142
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 23050 18184 23462
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17696 22710 17724 22918
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 18156 21622 18184 22986
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 20398 17816 20878
rect 18432 20602 18460 21422
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17788 19854 17816 20334
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17880 19446 17908 19654
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 18064 19310 18092 19654
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17604 17678 17632 18702
rect 18064 18290 18092 19246
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18248 17882 18276 18634
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17202 17632 17614
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17788 16794 17816 17070
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 14226 17816 14418
rect 17788 14198 17908 14226
rect 17880 14074 17908 14198
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17684 14000 17736 14006
rect 17682 13968 17684 13977
rect 17736 13968 17738 13977
rect 17682 13903 17738 13912
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 12986 17816 13398
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17880 12238 17908 13738
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 10674 17724 11494
rect 17788 11014 17816 11562
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17788 9994 17816 10950
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17880 9994 17908 10134
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17604 8294 17632 9930
rect 17880 9722 17908 9930
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17972 7954 18000 8298
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18064 7546 18092 7890
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7426 18184 16730
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18432 15434 18460 16526
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18340 14890 18368 14962
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14414 18368 14826
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12986 18276 13194
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18248 12170 18276 12786
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18248 11150 18276 12106
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18432 9654 18460 15370
rect 18616 12434 18644 18158
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16250 18736 16458
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14346 18736 14894
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18708 13938 18736 14282
rect 18788 14000 18840 14006
rect 18786 13968 18788 13977
rect 18840 13968 18842 13977
rect 18696 13932 18748 13938
rect 18786 13903 18842 13912
rect 18696 13874 18748 13880
rect 18616 12406 18828 12434
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18064 7398 18184 7426
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17972 6866 18000 7278
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17960 4140 18012 4146
rect 18064 4128 18092 7398
rect 18012 4100 18092 4128
rect 18144 4140 18196 4146
rect 17960 4082 18012 4088
rect 18144 4082 18196 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3738 17264 4014
rect 18156 3738 18184 4082
rect 18248 3942 18276 8978
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18432 4282 18460 4558
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 17788 3194 17816 3470
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 18248 2990 18276 3470
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 3126 18460 3334
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 17684 2916 17736 2922
rect 17684 2858 17736 2864
rect 17408 2848 17460 2854
rect 17696 2825 17724 2858
rect 17408 2790 17460 2796
rect 17682 2816 17738 2825
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 14844 1550 14964 1578
rect 14844 800 14872 1550
rect 15488 800 15516 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 800 16160 2314
rect 17420 800 17448 2790
rect 17682 2751 17738 2760
rect 18524 2446 18552 4422
rect 18616 2650 18644 5170
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18708 3602 18736 4966
rect 18800 3942 18828 12406
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 3058 18828 3334
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18892 2774 18920 25774
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 24886 19380 25094
rect 19340 24880 19392 24886
rect 19340 24822 19392 24828
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18984 24410 19012 24686
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23866 19104 24006
rect 19352 23866 19380 24142
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19076 22794 19104 23802
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19352 23118 19380 23666
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19076 22778 19196 22794
rect 19064 22772 19196 22778
rect 19116 22766 19196 22772
rect 19064 22714 19116 22720
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 19076 22030 19104 22578
rect 19168 22574 19196 22766
rect 19260 22642 19288 22918
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19444 22094 19472 36230
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19984 35760 20036 35766
rect 19984 35702 20036 35708
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19996 34678 20024 35702
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19524 34604 19576 34610
rect 19524 34546 19576 34552
rect 19536 34406 19564 34546
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19536 32978 19564 33458
rect 19524 32972 19576 32978
rect 19524 32914 19576 32920
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19524 32428 19576 32434
rect 19524 32370 19576 32376
rect 19536 31822 19564 32370
rect 19996 31958 20024 34614
rect 19984 31952 20036 31958
rect 19984 31894 20036 31900
rect 19524 31816 19576 31822
rect 19524 31758 19576 31764
rect 19984 31680 20036 31686
rect 19984 31622 20036 31628
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19996 31142 20024 31622
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19892 28076 19944 28082
rect 19892 28018 19944 28024
rect 19904 27384 19932 28018
rect 19996 27554 20024 29582
rect 20088 29322 20116 45358
rect 21180 37188 21232 37194
rect 21180 37130 21232 37136
rect 20260 37120 20312 37126
rect 20260 37062 20312 37068
rect 20168 36780 20220 36786
rect 20272 36768 20300 37062
rect 21192 36922 21220 37130
rect 21180 36916 21232 36922
rect 21180 36858 21232 36864
rect 21836 36854 21864 46854
rect 21824 36848 21876 36854
rect 21824 36790 21876 36796
rect 20220 36740 20300 36768
rect 20168 36722 20220 36728
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20180 36242 20208 36518
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 20272 36174 20300 36740
rect 21088 36780 21140 36786
rect 21088 36722 21140 36728
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20260 36168 20312 36174
rect 20260 36110 20312 36116
rect 20272 35290 20300 36110
rect 20260 35284 20312 35290
rect 20260 35226 20312 35232
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20180 34610 20208 34954
rect 20272 34678 20300 35226
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20260 34672 20312 34678
rect 20260 34614 20312 34620
rect 20168 34604 20220 34610
rect 20168 34546 20220 34552
rect 20168 34400 20220 34406
rect 20168 34342 20220 34348
rect 20180 33318 20208 34342
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20168 33312 20220 33318
rect 20168 33254 20220 33260
rect 20272 32366 20300 33458
rect 20260 32360 20312 32366
rect 20260 32302 20312 32308
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20180 31686 20208 32166
rect 20364 32026 20392 34886
rect 20456 34610 20484 36654
rect 21100 35698 21128 36722
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21100 35086 21128 35634
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 21088 35080 21140 35086
rect 21088 35022 21140 35028
rect 20444 34604 20496 34610
rect 20496 34564 20576 34592
rect 20444 34546 20496 34552
rect 20444 34468 20496 34474
rect 20444 34410 20496 34416
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20168 31680 20220 31686
rect 20168 31622 20220 31628
rect 20180 31278 20208 31622
rect 20168 31272 20220 31278
rect 20168 31214 20220 31220
rect 20272 30580 20300 31894
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20364 30734 20392 31282
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20272 30552 20392 30580
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 20088 29294 20208 29322
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 20088 28218 20116 29174
rect 20180 28914 20208 29294
rect 20272 29102 20300 29990
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20364 28937 20392 30552
rect 20350 28928 20406 28937
rect 20180 28886 20300 28914
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 19996 27526 20208 27554
rect 20076 27396 20128 27402
rect 19904 27356 20024 27384
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19892 27056 19944 27062
rect 19892 26998 19944 27004
rect 19904 26518 19932 26998
rect 19892 26512 19944 26518
rect 19892 26454 19944 26460
rect 19996 26382 20024 27356
rect 20076 27338 20128 27344
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25906 20024 26318
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19628 23322 19656 23666
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22710 20024 23122
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 20088 22094 20116 27338
rect 19352 22066 19472 22094
rect 19996 22066 20116 22094
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19352 21350 19380 22066
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19444 21146 19472 21898
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20346 20024 22066
rect 20074 21040 20130 21049
rect 20074 20975 20076 20984
rect 20128 20975 20130 20984
rect 20076 20946 20128 20952
rect 20180 20482 20208 27526
rect 20272 21690 20300 28886
rect 20350 28863 20406 28872
rect 20364 27606 20392 28863
rect 20352 27600 20404 27606
rect 20352 27542 20404 27548
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20364 22710 20392 23462
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20272 20942 20300 21490
rect 20364 21010 20392 22646
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20364 20602 20392 20946
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20180 20454 20300 20482
rect 19248 20324 19300 20330
rect 19996 20318 20116 20346
rect 19248 20266 19300 20272
rect 19260 19514 19288 20266
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19444 18970 19472 19722
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19996 18902 20024 20198
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19444 18290 19472 18702
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18426 20024 18702
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20088 18358 20116 20318
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19248 17536 19300 17542
rect 19352 17490 19380 17614
rect 19444 17542 19472 18226
rect 20180 18222 20208 19722
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 19300 17484 19380 17490
rect 19248 17478 19380 17484
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19260 17462 19380 17478
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16726 19288 17070
rect 19352 16998 19380 17462
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19444 15502 19472 17478
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19996 16590 20024 17478
rect 20272 17218 20300 20454
rect 20364 19446 20392 20538
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20088 17190 20300 17218
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19996 16114 20024 16526
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19536 15638 19564 15982
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20088 14498 20116 17190
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 15586 20208 16458
rect 20272 15706 20300 17070
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20364 15706 20392 15982
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20180 15558 20392 15586
rect 20088 14470 20300 14498
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13394 19380 13806
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 12986 19380 13330
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19444 12782 19472 13398
rect 19996 13258 20024 14214
rect 20088 13802 20116 14214
rect 20180 14074 20208 14350
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 20272 13138 20300 14470
rect 19996 13110 20300 13138
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19536 12442 19564 12854
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19996 12322 20024 13110
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20180 12442 20208 12854
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 19996 12294 20300 12322
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 10742 19472 11018
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 9722 19472 10406
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19260 8974 19288 9522
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19628 9178 19656 9454
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8498 19288 8910
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4622 19656 4966
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19352 4078 19380 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 4282 20024 5170
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20088 4146 20116 4422
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19156 3120 19208 3126
rect 19260 3097 19288 3878
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19156 3062 19208 3068
rect 19246 3088 19302 3097
rect 18708 2746 18920 2774
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18708 800 18736 2746
rect 19168 2446 19196 3062
rect 19246 3023 19302 3032
rect 19352 2650 19380 3470
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19444 2530 19472 3674
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20088 3058 20116 3470
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19892 2984 19944 2990
rect 19890 2952 19892 2961
rect 19984 2984 20036 2990
rect 19944 2952 19946 2961
rect 19984 2926 20036 2932
rect 19890 2887 19946 2896
rect 19352 2502 19472 2530
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19352 800 19380 2502
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2926
rect 20272 2514 20300 12294
rect 20364 6746 20392 15558
rect 20456 8378 20484 34410
rect 20548 33658 20576 34564
rect 20640 33862 20668 35022
rect 20996 34944 21048 34950
rect 20996 34886 21048 34892
rect 21008 33930 21036 34886
rect 21468 34066 21496 35090
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 21836 34746 21864 34954
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 21824 34604 21876 34610
rect 22112 34592 22140 47058
rect 24584 47048 24636 47054
rect 24584 46990 24636 46996
rect 24596 46578 24624 46990
rect 24584 46572 24636 46578
rect 24584 46514 24636 46520
rect 25148 46510 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25516 46034 25544 46990
rect 25792 46034 25820 49200
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 24124 45960 24176 45966
rect 24124 45902 24176 45908
rect 24136 45558 24164 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25320 45824 25372 45830
rect 25320 45766 25372 45772
rect 24124 45552 24176 45558
rect 24124 45494 24176 45500
rect 24136 41414 24164 45494
rect 25332 45490 25360 45766
rect 25424 45626 25452 45834
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 26712 45554 26740 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 28368 47054 28396 49200
rect 29368 47184 29420 47190
rect 29368 47126 29420 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28264 46912 28316 46918
rect 28264 46854 28316 46860
rect 28276 46578 28304 46854
rect 28264 46572 28316 46578
rect 28264 46514 28316 46520
rect 26436 45526 26740 45554
rect 25320 45484 25372 45490
rect 25320 45426 25372 45432
rect 25332 44198 25360 45426
rect 25320 44192 25372 44198
rect 25320 44134 25372 44140
rect 25872 44192 25924 44198
rect 25872 44134 25924 44140
rect 25504 43308 25556 43314
rect 25504 43250 25556 43256
rect 25228 42696 25280 42702
rect 25228 42638 25280 42644
rect 25240 42362 25268 42638
rect 25228 42356 25280 42362
rect 25228 42298 25280 42304
rect 25320 42220 25372 42226
rect 25320 42162 25372 42168
rect 24136 41386 24256 41414
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 22480 36242 22508 37062
rect 22560 36712 22612 36718
rect 22560 36654 22612 36660
rect 22468 36236 22520 36242
rect 22468 36178 22520 36184
rect 22480 35698 22508 36178
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22468 35488 22520 35494
rect 22468 35430 22520 35436
rect 22480 35018 22508 35430
rect 22572 35154 22600 36654
rect 22756 35630 22784 37198
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 23676 36854 23704 37062
rect 23664 36848 23716 36854
rect 23664 36790 23716 36796
rect 22928 36712 22980 36718
rect 22928 36654 22980 36660
rect 22940 36378 22968 36654
rect 22928 36372 22980 36378
rect 22928 36314 22980 36320
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 22744 35624 22796 35630
rect 22744 35566 22796 35572
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22468 35012 22520 35018
rect 22468 34954 22520 34960
rect 22192 34604 22244 34610
rect 22112 34564 22192 34592
rect 21824 34546 21876 34552
rect 22192 34546 22244 34552
rect 21456 34060 21508 34066
rect 21456 34002 21508 34008
rect 20720 33924 20772 33930
rect 20720 33866 20772 33872
rect 20996 33924 21048 33930
rect 20996 33866 21048 33872
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20548 32842 20576 33594
rect 20640 33522 20668 33798
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20536 32836 20588 32842
rect 20536 32778 20588 32784
rect 20640 31822 20668 32982
rect 20732 32026 20760 33866
rect 20812 33516 20864 33522
rect 20812 33458 20864 33464
rect 20720 32020 20772 32026
rect 20720 31962 20772 31968
rect 20824 31822 20852 33458
rect 21468 33114 21496 34002
rect 21836 33658 21864 34546
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21824 33652 21876 33658
rect 21824 33594 21876 33600
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 21456 33108 21508 33114
rect 21456 33050 21508 33056
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 20996 31952 21048 31958
rect 20996 31894 21048 31900
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20916 31754 20944 31826
rect 21008 31754 21036 31894
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 20904 31748 20956 31754
rect 20904 31690 20956 31696
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20548 31210 20576 31282
rect 20536 31204 20588 31210
rect 20536 31146 20588 31152
rect 20548 30394 20576 31146
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20732 29714 20760 30670
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 20824 30190 20852 30602
rect 20916 30258 20944 31078
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 21008 30054 21036 31690
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20732 29306 20760 29650
rect 21008 29578 21036 29990
rect 20996 29572 21048 29578
rect 20996 29514 21048 29520
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 21100 29186 21128 31758
rect 21180 30592 21232 30598
rect 21180 30534 21232 30540
rect 21192 30258 21220 30534
rect 21180 30252 21232 30258
rect 21180 30194 21232 30200
rect 21180 30116 21232 30122
rect 21180 30058 21232 30064
rect 20916 29158 21128 29186
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20824 28218 20852 28426
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27538 20760 27814
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20824 27402 20852 28018
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24206 20576 24550
rect 20640 24410 20668 24686
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20548 23730 20576 24142
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20548 23118 20576 23666
rect 20824 23526 20852 23802
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22778 20760 23054
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20824 22642 20852 23462
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20824 22030 20852 22578
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 20262 20576 21286
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 19310 20576 19858
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20640 18630 20668 21626
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20732 20942 20760 21422
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20466 20760 20878
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20824 19378 20852 20470
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20732 18290 20760 19178
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20824 18426 20852 18634
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20916 17626 20944 29158
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 21100 28626 21128 28970
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 21192 28200 21220 30058
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21560 29510 21588 29718
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21548 29096 21600 29102
rect 21546 29064 21548 29073
rect 21600 29064 21602 29073
rect 21546 28999 21602 29008
rect 21008 28172 21220 28200
rect 21008 27470 21036 28172
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21192 26790 21220 27338
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 21100 25702 21128 25842
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 21008 22778 21036 22986
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 21008 19514 21036 19654
rect 21100 19514 21128 20402
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21100 19174 21128 19450
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21008 18358 21036 19110
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 20824 17598 20944 17626
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20732 13938 20760 15506
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20732 13394 20760 13670
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20732 12434 20760 12786
rect 20640 12406 20760 12434
rect 20640 12238 20668 12406
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20456 8350 20668 8378
rect 20364 6718 20484 6746
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20364 4826 20392 5170
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20456 3942 20484 6718
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20640 2774 20668 8350
rect 20824 7562 20852 17598
rect 21008 17270 21036 17614
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15502 21128 15846
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 15026 21128 15438
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14482 20944 14758
rect 21100 14550 21128 14962
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 14006 20944 14418
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20916 12986 20944 13126
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21008 12306 21036 13874
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20456 2746 20668 2774
rect 20732 7534 20852 7562
rect 20456 2650 20484 2746
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20732 2582 20760 7534
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20824 4622 20852 4966
rect 21008 4826 21036 5170
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 3126 20852 4422
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 20916 3058 20944 3334
rect 21008 3126 21036 3402
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21100 2990 21128 3402
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20640 800 20668 2314
rect 21192 1902 21220 25298
rect 21468 25294 21496 26454
rect 21560 26382 21588 26862
rect 21652 26858 21680 32914
rect 21836 32910 21864 33458
rect 21928 32978 21956 33798
rect 22190 33552 22246 33561
rect 22190 33487 22192 33496
rect 22244 33487 22246 33496
rect 22192 33458 22244 33464
rect 21916 32972 21968 32978
rect 21916 32914 21968 32920
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 21744 31890 21772 31962
rect 21732 31884 21784 31890
rect 21732 31826 21784 31832
rect 21640 26852 21692 26858
rect 21640 26794 21692 26800
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21560 25294 21588 26318
rect 21744 25294 21772 31826
rect 22204 29850 22232 33458
rect 22744 32972 22796 32978
rect 22744 32914 22796 32920
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22296 31482 22324 32846
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 22296 30326 22324 31418
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21836 29170 21864 29446
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 22020 28490 22048 29650
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21928 27062 21956 27406
rect 22112 27402 22140 29514
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22204 29102 22232 29242
rect 22284 29164 22336 29170
rect 22480 29152 22508 29582
rect 22336 29124 22508 29152
rect 22284 29106 22336 29112
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22296 28150 22324 28698
rect 22480 28626 22508 29124
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22572 28490 22600 31758
rect 22756 31362 22784 32914
rect 22848 31754 22876 36110
rect 23216 35766 23244 36110
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 23032 34610 23060 35090
rect 23296 34944 23348 34950
rect 23296 34886 23348 34892
rect 23112 34740 23164 34746
rect 23112 34682 23164 34688
rect 22928 34604 22980 34610
rect 22928 34546 22980 34552
rect 23020 34604 23072 34610
rect 23020 34546 23072 34552
rect 22940 34490 22968 34546
rect 23124 34490 23152 34682
rect 23308 34542 23336 34886
rect 22940 34462 23152 34490
rect 23296 34536 23348 34542
rect 23296 34478 23348 34484
rect 23308 33590 23336 34478
rect 23388 33924 23440 33930
rect 23388 33866 23440 33872
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23204 33448 23256 33454
rect 23204 33390 23256 33396
rect 23020 33380 23072 33386
rect 23020 33322 23072 33328
rect 23032 32978 23060 33322
rect 23112 33312 23164 33318
rect 23112 33254 23164 33260
rect 23020 32972 23072 32978
rect 23020 32914 23072 32920
rect 23124 32910 23152 33254
rect 23112 32904 23164 32910
rect 23112 32846 23164 32852
rect 22848 31726 23060 31754
rect 23032 31657 23060 31726
rect 23018 31648 23074 31657
rect 23018 31583 23074 31592
rect 22756 31346 22876 31362
rect 22756 31340 22888 31346
rect 22756 31334 22836 31340
rect 22836 31282 22888 31288
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22204 27606 22232 28018
rect 22192 27600 22244 27606
rect 22192 27542 22244 27548
rect 22100 27396 22152 27402
rect 22100 27338 22152 27344
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 22112 26994 22140 27338
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21836 26518 21864 26794
rect 21824 26512 21876 26518
rect 21824 26454 21876 26460
rect 21836 26382 21864 26454
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 22112 26246 22140 26930
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22112 25498 22140 25774
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21284 3738 21312 21898
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21376 21010 21404 21830
rect 22112 21690 22140 23054
rect 22296 22094 22324 28086
rect 22572 28082 22600 28426
rect 22756 28150 22784 28562
rect 22744 28144 22796 28150
rect 22744 28086 22796 28092
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22848 27946 22876 31282
rect 23032 30326 23060 31583
rect 23216 31482 23244 33390
rect 23308 32910 23336 33526
rect 23400 33318 23428 33866
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23768 33658 23796 33798
rect 23756 33652 23808 33658
rect 23756 33594 23808 33600
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23860 32910 23888 33458
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23584 32434 23612 32710
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23480 32360 23532 32366
rect 23480 32302 23532 32308
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 23216 31346 23244 31418
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23124 31226 23152 31282
rect 23124 31198 23244 31226
rect 23216 30802 23244 31198
rect 23204 30796 23256 30802
rect 23204 30738 23256 30744
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 23216 29646 23244 30738
rect 23492 30682 23520 32302
rect 23768 31754 23796 32438
rect 23860 31890 23888 32846
rect 23848 31884 23900 31890
rect 23848 31826 23900 31832
rect 23756 31748 23808 31754
rect 23756 31690 23808 31696
rect 23572 31204 23624 31210
rect 23572 31146 23624 31152
rect 23400 30666 23520 30682
rect 23584 30666 23612 31146
rect 23768 30938 23796 31690
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23388 30660 23520 30666
rect 23440 30654 23520 30660
rect 23388 30602 23440 30608
rect 23492 29646 23520 30654
rect 23572 30660 23624 30666
rect 23572 30602 23624 30608
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23216 29170 23244 29582
rect 23584 29578 23612 30126
rect 23676 29782 23704 30194
rect 23664 29776 23716 29782
rect 23664 29718 23716 29724
rect 23388 29572 23440 29578
rect 23388 29514 23440 29520
rect 23572 29572 23624 29578
rect 23572 29514 23624 29520
rect 23400 29306 23428 29514
rect 23676 29510 23704 29718
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23032 28422 23060 29106
rect 23492 29034 23520 29242
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23676 28626 23704 29446
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22836 27940 22888 27946
rect 22836 27882 22888 27888
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22572 26450 22600 27814
rect 22940 27470 22968 28018
rect 23216 28014 23244 28358
rect 23204 28008 23256 28014
rect 23204 27950 23256 27956
rect 23584 27674 23612 28494
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22848 26450 22876 26862
rect 22940 26790 22968 27406
rect 23032 27062 23060 27406
rect 23020 27056 23072 27062
rect 23020 26998 23072 27004
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22572 25838 22600 26386
rect 23032 26314 23060 26998
rect 23492 26994 23520 27474
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22848 24070 22876 24550
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22480 23322 22508 23598
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22642 22508 22918
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23216 22234 23244 22510
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 22204 22066 22324 22094
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 21560 20466 21588 21490
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22112 20602 22140 20810
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21560 19854 21588 20402
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21560 18698 21588 19654
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21836 19310 21864 19382
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21836 18970 21864 19246
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21836 18290 21864 18906
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17678 21496 18022
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17338 22140 17546
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21468 16046 21496 16458
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 21376 15026 21404 15370
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21376 14346 21404 14962
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21468 3618 21496 15982
rect 21744 15570 21772 16526
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21836 16114 21864 16390
rect 22112 16182 22140 16934
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 22204 15910 22232 22066
rect 23308 22030 23336 23054
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23124 21078 23152 21354
rect 23308 21350 23336 21966
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22940 20330 22968 20946
rect 23308 20942 23336 21286
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23492 20466 23520 21490
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 22928 20324 22980 20330
rect 22928 20266 22980 20272
rect 22940 19310 22968 20266
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19446 23060 20198
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21744 15162 21772 15506
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21928 15094 21956 15506
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22020 15026 22048 15302
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22112 14822 22140 15438
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22204 15162 22232 15370
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22296 15026 22324 17138
rect 22664 16590 22692 17274
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16182 22784 16390
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22480 15094 22508 15302
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22664 15026 22692 15302
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 13870 21680 14350
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21652 13530 21680 13806
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21836 12850 21864 14010
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21928 12986 21956 13194
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21560 4622 21588 4966
rect 21652 4826 21680 5646
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21732 4208 21784 4214
rect 21730 4176 21732 4185
rect 21824 4208 21876 4214
rect 21784 4176 21786 4185
rect 21824 4150 21876 4156
rect 21730 4111 21786 4120
rect 21836 4010 21864 4150
rect 22112 4078 22140 5102
rect 22204 4622 22232 5510
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22296 4826 22324 5170
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22388 4214 22416 4966
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21376 3590 21496 3618
rect 21916 3596 21968 3602
rect 21376 2825 21404 3590
rect 21916 3538 21968 3544
rect 21928 3505 21956 3538
rect 21914 3496 21970 3505
rect 21914 3431 21970 3440
rect 21454 3360 21510 3369
rect 21454 3295 21510 3304
rect 21468 2922 21496 3295
rect 22020 3058 22048 3878
rect 22098 3632 22154 3641
rect 22204 3602 22232 4150
rect 22480 4146 22508 4422
rect 22848 4282 22876 4558
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22940 4146 22968 19246
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23492 17882 23520 18158
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23676 17678 23704 20334
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23768 18834 23796 19246
rect 23756 18828 23808 18834
rect 23756 18770 23808 18776
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23032 17270 23060 17478
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23308 10674 23336 17614
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23400 16182 23428 16526
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23584 15910 23612 17070
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 14958 23612 15846
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23860 12434 23888 21966
rect 23492 12406 23888 12434
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 22098 3567 22154 3576
rect 22192 3596 22244 3602
rect 22112 3398 22140 3567
rect 22192 3538 22244 3544
rect 23032 3534 23060 4966
rect 23020 3528 23072 3534
rect 22650 3496 22706 3505
rect 23020 3470 23072 3476
rect 22650 3431 22652 3440
rect 22704 3431 22706 3440
rect 22652 3402 22704 3408
rect 23308 3398 23336 10610
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23400 3505 23428 4082
rect 23386 3496 23442 3505
rect 23386 3431 23442 3440
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 22204 3126 22232 3334
rect 22192 3120 22244 3126
rect 22284 3120 22336 3126
rect 22192 3062 22244 3068
rect 22282 3088 22284 3097
rect 22336 3088 22338 3097
rect 22008 3052 22060 3058
rect 22282 3023 22338 3032
rect 22008 2994 22060 3000
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21362 2816 21418 2825
rect 21362 2751 21418 2760
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21180 1896 21232 1902
rect 21180 1838 21232 1844
rect 21928 800 21956 2314
rect 22572 800 22600 2926
rect 22836 2916 22888 2922
rect 23020 2916 23072 2922
rect 22888 2876 23020 2904
rect 22836 2858 22888 2864
rect 23020 2858 23072 2864
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23216 800 23244 2790
rect 23400 2650 23428 3431
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23492 2310 23520 12406
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23584 2446 23612 4422
rect 23848 4208 23900 4214
rect 23848 4150 23900 4156
rect 23860 3398 23888 4150
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23768 3194 23796 3334
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23952 2038 23980 33594
rect 24030 24984 24086 24993
rect 24030 24919 24032 24928
rect 24084 24919 24086 24928
rect 24032 24890 24084 24896
rect 24228 23186 24256 41386
rect 25136 37936 25188 37942
rect 25136 37878 25188 37884
rect 25044 37800 25096 37806
rect 25044 37742 25096 37748
rect 25056 37466 25084 37742
rect 25044 37460 25096 37466
rect 25044 37402 25096 37408
rect 24860 36712 24912 36718
rect 24860 36654 24912 36660
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24412 33114 24440 35974
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24504 34202 24532 34478
rect 24492 34196 24544 34202
rect 24492 34138 24544 34144
rect 24780 34134 24808 34614
rect 24768 34128 24820 34134
rect 24768 34070 24820 34076
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24780 33590 24808 33866
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24872 33114 24900 36654
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24964 35290 24992 36518
rect 25148 36378 25176 37878
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 25136 36372 25188 36378
rect 25136 36314 25188 36320
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 24964 35170 24992 35226
rect 24964 35142 25176 35170
rect 24952 35012 25004 35018
rect 24952 34954 25004 34960
rect 24964 34066 24992 34954
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25056 33658 25084 33934
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25148 33538 25176 35142
rect 25240 35086 25268 36722
rect 25228 35080 25280 35086
rect 25228 35022 25280 35028
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 25056 33510 25176 33538
rect 25240 33522 25268 34002
rect 25228 33516 25280 33522
rect 24400 33108 24452 33114
rect 24400 33050 24452 33056
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 32570 24900 33050
rect 25056 32910 25084 33510
rect 25228 33458 25280 33464
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 25148 33046 25176 33254
rect 25136 33040 25188 33046
rect 25136 32982 25188 32988
rect 25044 32904 25096 32910
rect 25228 32904 25280 32910
rect 25096 32864 25228 32892
rect 25044 32846 25096 32852
rect 25228 32846 25280 32852
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 24780 31822 24808 32370
rect 25056 32298 25084 32846
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 25332 31822 25360 42162
rect 25412 34944 25464 34950
rect 25412 34886 25464 34892
rect 25424 33998 25452 34886
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 24780 31346 24808 31758
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24412 30870 24440 31078
rect 24400 30864 24452 30870
rect 24780 30818 24808 31282
rect 24400 30806 24452 30812
rect 24412 30258 24440 30806
rect 24688 30790 24808 30818
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24596 29034 24624 30330
rect 24688 30258 24716 30790
rect 24768 30660 24820 30666
rect 24768 30602 24820 30608
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24688 29646 24716 30194
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24596 28150 24624 28494
rect 24584 28144 24636 28150
rect 24584 28086 24636 28092
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24412 26790 24440 27338
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24504 26450 24532 27950
rect 24596 27538 24624 28086
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24584 27532 24636 27538
rect 24584 27474 24636 27480
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24688 25294 24716 27882
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 24400 25152 24452 25158
rect 24400 25094 24452 25100
rect 24412 24886 24440 25094
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 24308 24812 24360 24818
rect 24676 24812 24728 24818
rect 24308 24754 24360 24760
rect 24596 24772 24676 24800
rect 24320 24721 24348 24754
rect 24306 24712 24362 24721
rect 24306 24647 24362 24656
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 24596 22030 24624 24772
rect 24676 24754 24728 24760
rect 24780 24682 24808 30602
rect 24860 29776 24912 29782
rect 24860 29718 24912 29724
rect 24872 29170 24900 29718
rect 25148 29578 25176 31282
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25240 30054 25268 30194
rect 25228 30048 25280 30054
rect 25226 30016 25228 30025
rect 25280 30016 25282 30025
rect 25226 29951 25282 29960
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 24872 28558 24900 29106
rect 24950 29064 25006 29073
rect 24950 28999 25006 29008
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24964 27962 24992 28999
rect 24872 27934 24992 27962
rect 25056 27962 25084 29242
rect 25148 29034 25176 29514
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25136 29028 25188 29034
rect 25136 28970 25188 28976
rect 25136 28416 25188 28422
rect 25136 28358 25188 28364
rect 25148 28150 25176 28358
rect 25136 28144 25188 28150
rect 25136 28086 25188 28092
rect 25240 28082 25268 29446
rect 25332 28762 25360 31758
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25424 29850 25452 29990
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25320 28756 25372 28762
rect 25320 28698 25372 28704
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25056 27934 25176 27962
rect 24872 25906 24900 27934
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 25056 27402 25084 27814
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 25056 26858 25084 27338
rect 25044 26852 25096 26858
rect 25044 26794 25096 26800
rect 25056 26382 25084 26794
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25148 25906 25176 27934
rect 25424 27606 25452 28494
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25332 26926 25360 27406
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25044 25832 25096 25838
rect 25044 25774 25096 25780
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24872 24886 24900 25162
rect 24860 24880 24912 24886
rect 24858 24848 24860 24857
rect 24912 24848 24914 24857
rect 24858 24783 24914 24792
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24688 24138 24716 24550
rect 25056 24410 25084 25774
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 25498 25268 25638
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25332 25294 25360 26862
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25424 25906 25452 26182
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25148 24886 25176 25230
rect 25226 24984 25282 24993
rect 25226 24919 25282 24928
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 25148 24410 25176 24822
rect 25240 24818 25268 24919
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25226 24712 25282 24721
rect 25226 24647 25282 24656
rect 25240 24614 25268 24647
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25332 24274 25360 25230
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25056 23526 25084 23666
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 25056 23118 25084 23462
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25056 22642 25084 23054
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25056 22030 25084 22578
rect 25424 22094 25452 23122
rect 25516 22574 25544 43250
rect 25884 41414 25912 44134
rect 25964 43104 26016 43110
rect 25964 43046 26016 43052
rect 25976 42770 26004 43046
rect 25964 42764 26016 42770
rect 25964 42706 26016 42712
rect 25700 41386 25912 41414
rect 25596 33312 25648 33318
rect 25596 33254 25648 33260
rect 25608 29170 25636 33254
rect 25700 31770 25728 41386
rect 26240 37732 26292 37738
rect 26240 37674 26292 37680
rect 26148 37664 26200 37670
rect 26148 37606 26200 37612
rect 26160 36786 26188 37606
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26252 35630 26280 37674
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26252 35170 26280 35566
rect 26160 35154 26280 35170
rect 26148 35148 26280 35154
rect 26200 35142 26280 35148
rect 26148 35090 26200 35096
rect 25964 35012 26016 35018
rect 25964 34954 26016 34960
rect 25976 34474 26004 34954
rect 26148 34944 26200 34950
rect 26148 34886 26200 34892
rect 26056 34740 26108 34746
rect 26056 34682 26108 34688
rect 25964 34468 26016 34474
rect 25964 34410 26016 34416
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25792 33114 25820 33458
rect 25872 33312 25924 33318
rect 25872 33254 25924 33260
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25780 32768 25832 32774
rect 25780 32710 25832 32716
rect 25792 32434 25820 32710
rect 25884 32502 25912 33254
rect 25872 32496 25924 32502
rect 26068 32450 26096 34682
rect 26160 33522 26188 34886
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26160 32910 26188 33458
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26160 32502 26188 32846
rect 25872 32438 25924 32444
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25884 32230 25912 32438
rect 25976 32422 26096 32450
rect 26148 32496 26200 32502
rect 26148 32438 26200 32444
rect 25872 32224 25924 32230
rect 25872 32166 25924 32172
rect 25976 32178 26004 32422
rect 25976 32150 26188 32178
rect 25700 31742 26096 31770
rect 25976 31726 26096 31742
rect 25688 31136 25740 31142
rect 25688 31078 25740 31084
rect 25700 30190 25728 31078
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25688 30184 25740 30190
rect 25688 30126 25740 30132
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25792 28218 25820 30194
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25608 26382 25636 27814
rect 25976 26874 26004 31726
rect 26160 29306 26188 32150
rect 26252 31686 26280 35142
rect 26332 32836 26384 32842
rect 26332 32778 26384 32784
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26252 29714 26280 31622
rect 26344 31498 26372 32778
rect 26436 31754 26464 45526
rect 27252 37324 27304 37330
rect 27252 37266 27304 37272
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 27080 36718 27108 37062
rect 27264 36922 27292 37266
rect 27252 36916 27304 36922
rect 27252 36858 27304 36864
rect 27068 36712 27120 36718
rect 27068 36654 27120 36660
rect 26976 35692 27028 35698
rect 26976 35634 27028 35640
rect 26988 35290 27016 35634
rect 27160 35488 27212 35494
rect 27160 35430 27212 35436
rect 26976 35284 27028 35290
rect 26976 35226 27028 35232
rect 26988 34610 27016 35226
rect 27172 35018 27200 35430
rect 27160 35012 27212 35018
rect 27160 34954 27212 34960
rect 26976 34604 27028 34610
rect 26976 34546 27028 34552
rect 26976 33856 27028 33862
rect 26976 33798 27028 33804
rect 26988 33522 27016 33798
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26436 31726 26648 31754
rect 26344 31470 26556 31498
rect 26332 31408 26384 31414
rect 26332 31350 26384 31356
rect 26344 30938 26372 31350
rect 26528 31210 26556 31470
rect 26516 31204 26568 31210
rect 26516 31146 26568 31152
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 26344 29238 26372 30874
rect 26332 29232 26384 29238
rect 26332 29174 26384 29180
rect 26054 29064 26110 29073
rect 26054 28999 26110 29008
rect 26068 28490 26096 28999
rect 26056 28484 26108 28490
rect 26056 28426 26108 28432
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26344 28082 26372 28358
rect 26528 28150 26556 31146
rect 26516 28144 26568 28150
rect 26516 28086 26568 28092
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26160 27674 26188 27814
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 25976 26846 26096 26874
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25608 25974 25636 26318
rect 25964 26240 26016 26246
rect 25964 26182 26016 26188
rect 25596 25968 25648 25974
rect 25596 25910 25648 25916
rect 25976 25702 26004 26182
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25608 25362 25636 25638
rect 25596 25356 25648 25362
rect 25596 25298 25648 25304
rect 25976 24954 26004 25638
rect 25964 24948 26016 24954
rect 25964 24890 26016 24896
rect 25976 24750 26004 24890
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 25424 22066 25544 22094
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 25056 21622 25084 21830
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 24044 21146 24072 21422
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 24780 20942 24808 21286
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24780 20466 24808 20878
rect 25056 20534 25084 21558
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25044 20528 25096 20534
rect 25044 20470 25096 20476
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24780 19854 24808 20402
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24872 18902 24900 19246
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 15026 24072 15846
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 15162 24440 15438
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24412 14822 24440 15098
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24504 4214 24532 18702
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24596 3058 24624 3470
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 23940 2032 23992 2038
rect 23940 1974 23992 1980
rect 24504 800 24532 2314
rect 24688 1970 24716 18702
rect 24964 14618 24992 20334
rect 25148 18306 25176 20810
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25332 19378 25360 19722
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25240 18834 25268 19314
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25240 18698 25268 18770
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25148 18278 25268 18306
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3126 24808 3878
rect 24872 3641 24900 11018
rect 25148 4214 25176 18158
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 24858 3632 24914 3641
rect 24858 3567 24914 3576
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 24872 2961 24900 3062
rect 24858 2952 24914 2961
rect 24858 2887 24914 2896
rect 25056 2650 25084 4082
rect 25240 3466 25268 18278
rect 25424 18154 25452 19722
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25424 4146 25452 18090
rect 25516 17218 25544 22066
rect 25608 21554 25636 23666
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25608 18086 25636 21490
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25792 18290 25820 20470
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25792 17542 25820 18226
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25884 17746 25912 18022
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25516 17190 25636 17218
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25516 15570 25544 15846
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25608 3602 25636 17190
rect 25976 11762 26004 22510
rect 26068 16522 26096 26846
rect 26238 24848 26294 24857
rect 26238 24783 26240 24792
rect 26292 24783 26294 24792
rect 26240 24754 26292 24760
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 26344 23866 26372 24074
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 26620 22506 26648 31726
rect 26988 30938 27016 32370
rect 27160 31816 27212 31822
rect 27160 31758 27212 31764
rect 26976 30932 27028 30938
rect 26976 30874 27028 30880
rect 26700 30728 26752 30734
rect 26700 30670 26752 30676
rect 26712 29782 26740 30670
rect 26792 30660 26844 30666
rect 26792 30602 26844 30608
rect 26700 29776 26752 29782
rect 26700 29718 26752 29724
rect 26712 28626 26740 29718
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 26712 24070 26740 24754
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26608 22500 26660 22506
rect 26608 22442 26660 22448
rect 26606 21040 26662 21049
rect 26606 20975 26608 20984
rect 26660 20975 26662 20984
rect 26608 20946 26660 20952
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 26344 20602 26372 20810
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26160 19718 26188 20402
rect 26620 20058 26648 20402
rect 26608 20052 26660 20058
rect 26608 19994 26660 20000
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 26160 18766 26188 19654
rect 26436 19378 26464 19790
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26160 17338 26188 17682
rect 26252 17610 26280 18566
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26252 17202 26280 17546
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25976 11082 26004 11698
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25318 3496 25374 3505
rect 25228 3460 25280 3466
rect 25318 3431 25320 3440
rect 25228 3402 25280 3408
rect 25372 3431 25374 3440
rect 25320 3402 25372 3408
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 25148 800 25176 2926
rect 25792 2854 25820 3130
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25700 2446 25728 2790
rect 26344 2650 26372 18158
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26804 2514 26832 30602
rect 26976 30116 27028 30122
rect 26976 30058 27028 30064
rect 26988 29714 27016 30058
rect 26976 29708 27028 29714
rect 26976 29650 27028 29656
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 26976 29572 27028 29578
rect 26976 29514 27028 29520
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26896 27946 26924 28902
rect 26988 28762 27016 29514
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 27080 28558 27108 29582
rect 27172 29306 27200 31758
rect 27264 30598 27292 36858
rect 27528 35624 27580 35630
rect 27528 35566 27580 35572
rect 29000 35624 29052 35630
rect 29000 35566 29052 35572
rect 27540 34678 27568 35566
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 27620 35148 27672 35154
rect 27620 35090 27672 35096
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27632 32570 27660 35090
rect 28644 34610 28672 35430
rect 29012 34746 29040 35566
rect 28816 34740 28868 34746
rect 28816 34682 28868 34688
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 28828 34610 28856 34682
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28632 34604 28684 34610
rect 28632 34546 28684 34552
rect 28816 34604 28868 34610
rect 28868 34564 28948 34592
rect 28816 34546 28868 34552
rect 28460 34134 28488 34546
rect 28448 34128 28500 34134
rect 28448 34070 28500 34076
rect 28540 34128 28592 34134
rect 28540 34070 28592 34076
rect 28920 34082 28948 34564
rect 29000 34468 29052 34474
rect 29000 34410 29052 34416
rect 29012 34202 29040 34410
rect 29000 34196 29052 34202
rect 29000 34138 29052 34144
rect 28998 34096 29054 34105
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 28448 33992 28500 33998
rect 28448 33934 28500 33940
rect 27724 33454 27752 33934
rect 27896 33924 27948 33930
rect 27896 33866 27948 33872
rect 27908 33522 27936 33866
rect 28460 33522 28488 33934
rect 28552 33561 28580 34070
rect 28920 34054 28998 34082
rect 28998 34031 29054 34040
rect 29184 34060 29236 34066
rect 29184 34002 29236 34008
rect 29196 33833 29224 34002
rect 29274 33960 29330 33969
rect 29274 33895 29276 33904
rect 29328 33895 29330 33904
rect 29276 33866 29328 33872
rect 29182 33824 29238 33833
rect 29182 33759 29238 33768
rect 28816 33584 28868 33590
rect 28538 33552 28594 33561
rect 27896 33516 27948 33522
rect 27896 33458 27948 33464
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 28448 33516 28500 33522
rect 28868 33532 29316 33538
rect 28816 33526 29316 33532
rect 28828 33522 29316 33526
rect 28828 33516 29328 33522
rect 28828 33510 29276 33516
rect 28538 33487 28594 33496
rect 28448 33458 28500 33464
rect 29276 33458 29328 33464
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27724 32774 27752 33390
rect 27908 33318 27936 33458
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 28092 32910 28120 33458
rect 28460 33386 28488 33458
rect 28448 33380 28500 33386
rect 28448 33322 28500 33328
rect 29092 33040 29144 33046
rect 29092 32982 29144 32988
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 28448 32904 28500 32910
rect 28448 32846 28500 32852
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 27988 32836 28040 32842
rect 27988 32778 28040 32784
rect 27712 32768 27764 32774
rect 27712 32710 27764 32716
rect 27620 32564 27672 32570
rect 27620 32506 27672 32512
rect 27620 32428 27672 32434
rect 27620 32370 27672 32376
rect 27528 31952 27580 31958
rect 27528 31894 27580 31900
rect 27540 31686 27568 31894
rect 27632 31890 27660 32370
rect 27620 31884 27672 31890
rect 27620 31826 27672 31832
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 27540 31346 27568 31622
rect 27528 31340 27580 31346
rect 27528 31282 27580 31288
rect 27344 31136 27396 31142
rect 27344 31078 27396 31084
rect 27252 30592 27304 30598
rect 27252 30534 27304 30540
rect 27264 30258 27292 30534
rect 27252 30252 27304 30258
rect 27252 30194 27304 30200
rect 27356 30025 27384 31078
rect 27436 30184 27488 30190
rect 27436 30126 27488 30132
rect 27342 30016 27398 30025
rect 27342 29951 27398 29960
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27172 28558 27200 29242
rect 27068 28552 27120 28558
rect 26988 28512 27068 28540
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26988 26994 27016 28512
rect 27068 28494 27120 28500
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 27080 27062 27108 27338
rect 27068 27056 27120 27062
rect 27068 26998 27120 27004
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 26988 25906 27016 26930
rect 27356 26382 27384 29951
rect 27448 29782 27476 30126
rect 27436 29776 27488 29782
rect 27436 29718 27488 29724
rect 27620 29572 27672 29578
rect 27620 29514 27672 29520
rect 27632 29034 27660 29514
rect 27620 29028 27672 29034
rect 27620 28970 27672 28976
rect 27724 28082 27752 31690
rect 28000 31657 28028 32778
rect 28264 32496 28316 32502
rect 28264 32438 28316 32444
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 27986 31648 28042 31657
rect 27986 31583 28042 31592
rect 27804 31272 27856 31278
rect 27804 31214 27856 31220
rect 27816 30938 27844 31214
rect 27804 30932 27856 30938
rect 27804 30874 27856 30880
rect 28000 28558 28028 31583
rect 28184 31482 28212 31758
rect 28276 31754 28304 32438
rect 28460 31822 28488 32846
rect 28724 32836 28776 32842
rect 28724 32778 28776 32784
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28264 31748 28316 31754
rect 28264 31690 28316 31696
rect 28172 31476 28224 31482
rect 28172 31418 28224 31424
rect 28172 30864 28224 30870
rect 28172 30806 28224 30812
rect 28184 30394 28212 30806
rect 28276 30666 28304 31690
rect 28448 31408 28500 31414
rect 28448 31350 28500 31356
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28264 30660 28316 30666
rect 28264 30602 28316 30608
rect 28172 30388 28224 30394
rect 28172 30330 28224 30336
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27712 27532 27764 27538
rect 27712 27474 27764 27480
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27448 26382 27476 26522
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 25226 26924 25638
rect 26884 25220 26936 25226
rect 26884 25162 26936 25168
rect 26988 24954 27016 25842
rect 27080 25430 27108 26318
rect 27252 26308 27304 26314
rect 27252 26250 27304 26256
rect 27068 25424 27120 25430
rect 27068 25366 27120 25372
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26988 24290 27016 24890
rect 26896 24262 27016 24290
rect 27264 24274 27292 26250
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27356 24886 27384 25638
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27632 24818 27660 25162
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27252 24268 27304 24274
rect 26896 23730 26924 24262
rect 27252 24210 27304 24216
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26988 23866 27016 24142
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26884 23724 26936 23730
rect 26884 23666 26936 23672
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27172 22710 27200 22918
rect 27160 22704 27212 22710
rect 27160 22646 27212 22652
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26988 21962 27016 22510
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 26988 21418 27016 21898
rect 26976 21412 27028 21418
rect 26976 21354 27028 21360
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27158 15600 27214 15609
rect 27158 15535 27160 15544
rect 27212 15535 27214 15544
rect 27160 15506 27212 15512
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 26974 4176 27030 4185
rect 26974 4111 27030 4120
rect 26988 4010 27016 4111
rect 26976 4004 27028 4010
rect 26976 3946 27028 3952
rect 27172 3602 27200 8910
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 27264 2774 27292 17070
rect 27356 16590 27384 24006
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27448 18290 27476 19790
rect 27632 19514 27660 20334
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27632 18358 27660 18702
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 27356 13938 27384 16526
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27632 16182 27660 16390
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 27356 3602 27384 4966
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27632 3602 27660 4014
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27632 3369 27660 3538
rect 27618 3360 27674 3369
rect 27618 3295 27674 3304
rect 27724 2774 27752 27474
rect 27908 26926 27936 28358
rect 28184 27962 28212 30330
rect 28276 30054 28304 30602
rect 28368 30394 28396 30670
rect 28356 30388 28408 30394
rect 28356 30330 28408 30336
rect 28264 30048 28316 30054
rect 28264 29990 28316 29996
rect 28460 29850 28488 31350
rect 28552 30734 28580 32166
rect 28644 32026 28672 32370
rect 28632 32020 28684 32026
rect 28632 31962 28684 31968
rect 28736 31754 28764 32778
rect 29012 31822 29040 32846
rect 29104 32434 29132 32982
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 28644 31726 28764 31754
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28448 29844 28500 29850
rect 28448 29786 28500 29792
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 28276 28937 28304 28970
rect 28262 28928 28318 28937
rect 28262 28863 28318 28872
rect 28092 27934 28212 27962
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 28092 26450 28120 27934
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 27470 28212 27814
rect 28276 27606 28304 28863
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28264 27600 28316 27606
rect 28264 27542 28316 27548
rect 28172 27464 28224 27470
rect 28368 27452 28396 28018
rect 28172 27406 28224 27412
rect 28276 27424 28396 27452
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28184 27062 28212 27270
rect 28172 27056 28224 27062
rect 28172 26998 28224 27004
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28276 26314 28304 27424
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 28276 24614 28304 26250
rect 28644 24750 28672 31726
rect 29012 31142 29040 31758
rect 29288 31754 29316 33458
rect 29196 31726 29316 31754
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28816 30184 28868 30190
rect 28816 30126 28868 30132
rect 28828 29170 28856 30126
rect 28816 29164 28868 29170
rect 28816 29106 28868 29112
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28736 28014 28764 28494
rect 28724 28008 28776 28014
rect 28724 27950 28776 27956
rect 28828 25906 28856 29106
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28632 24744 28684 24750
rect 28632 24686 28684 24692
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28828 24342 28856 25842
rect 28816 24336 28868 24342
rect 28816 24278 28868 24284
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 27908 23798 27936 24006
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 28000 23322 28028 24074
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 27804 20528 27856 20534
rect 27802 20496 27804 20505
rect 27856 20496 27858 20505
rect 27802 20431 27858 20440
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 27802 19952 27858 19961
rect 27858 19910 27936 19938
rect 27802 19887 27804 19896
rect 27856 19887 27858 19896
rect 27804 19858 27856 19864
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27816 18902 27844 19722
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27816 18698 27844 18838
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27908 18426 27936 19910
rect 28276 19854 28304 20198
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28368 19718 28396 20742
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 28000 18970 28028 19246
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 28092 18290 28120 19450
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 28276 17882 28304 18158
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28368 8974 28396 19654
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28460 18834 28488 19314
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28552 16454 28580 23054
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28736 18766 28764 19314
rect 28816 19304 28868 19310
rect 28816 19246 28868 19252
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28828 18698 28856 19246
rect 28816 18692 28868 18698
rect 28816 18634 28868 18640
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28920 3194 28948 30194
rect 29196 29510 29224 31726
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29288 30666 29316 31078
rect 29276 30660 29328 30666
rect 29276 30602 29328 30608
rect 29184 29504 29236 29510
rect 29184 29446 29236 29452
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 29104 28082 29132 28494
rect 29092 28076 29144 28082
rect 29092 28018 29144 28024
rect 29000 23792 29052 23798
rect 29000 23734 29052 23740
rect 29012 23322 29040 23734
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 29012 20398 29040 21898
rect 29380 21010 29408 47126
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41206 49314 41318 50000
rect 40788 49286 41318 49314
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 31116 47048 31168 47054
rect 31116 46990 31168 46996
rect 29644 35692 29696 35698
rect 29644 35634 29696 35640
rect 29656 35290 29684 35634
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 29644 35284 29696 35290
rect 29644 35226 29696 35232
rect 29736 34536 29788 34542
rect 30024 34524 30052 35430
rect 29788 34496 30052 34524
rect 29736 34478 29788 34484
rect 29736 34400 29788 34406
rect 29736 34342 29788 34348
rect 29748 34202 29776 34342
rect 29736 34196 29788 34202
rect 29736 34138 29788 34144
rect 29644 34128 29696 34134
rect 29644 34070 29696 34076
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 29472 33658 29500 33934
rect 29460 33652 29512 33658
rect 29460 33594 29512 33600
rect 29458 33416 29514 33425
rect 29458 33351 29460 33360
rect 29512 33351 29514 33360
rect 29460 33322 29512 33328
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 29564 33114 29592 33254
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 29656 29850 29684 34070
rect 29736 33992 29788 33998
rect 29734 33960 29736 33969
rect 29788 33960 29790 33969
rect 29734 33895 29790 33904
rect 30024 33572 30052 34496
rect 30104 34536 30156 34542
rect 30104 34478 30156 34484
rect 30116 34202 30144 34478
rect 30196 34400 30248 34406
rect 30196 34342 30248 34348
rect 30104 34196 30156 34202
rect 30104 34138 30156 34144
rect 30102 34096 30158 34105
rect 30102 34031 30158 34040
rect 30116 33998 30144 34031
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30104 33584 30156 33590
rect 30024 33544 30104 33572
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29748 32910 29776 33458
rect 30024 33318 30052 33544
rect 30104 33526 30156 33532
rect 30208 33522 30236 34342
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30196 33516 30248 33522
rect 30196 33458 30248 33464
rect 30472 33448 30524 33454
rect 30378 33416 30434 33425
rect 30472 33390 30524 33396
rect 30378 33351 30380 33360
rect 30432 33351 30434 33360
rect 30380 33322 30432 33328
rect 30484 33318 30512 33390
rect 30012 33312 30064 33318
rect 30012 33254 30064 33260
rect 30288 33312 30340 33318
rect 30288 33254 30340 33260
rect 30472 33312 30524 33318
rect 30472 33254 30524 33260
rect 30300 33114 30328 33254
rect 30288 33108 30340 33114
rect 30288 33050 30340 33056
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 30576 32502 30604 33798
rect 30668 33522 30696 34138
rect 31024 34060 31076 34066
rect 31024 34002 31076 34008
rect 30932 33992 30984 33998
rect 30932 33934 30984 33940
rect 30748 33924 30800 33930
rect 30748 33866 30800 33872
rect 30760 33833 30788 33866
rect 30746 33824 30802 33833
rect 30746 33759 30802 33768
rect 30944 33590 30972 33934
rect 30932 33584 30984 33590
rect 30932 33526 30984 33532
rect 30656 33516 30708 33522
rect 30656 33458 30708 33464
rect 30668 33114 30696 33458
rect 30932 33312 30984 33318
rect 31036 33266 31064 34002
rect 30984 33260 31064 33266
rect 30932 33254 31064 33260
rect 30944 33238 31064 33254
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30656 32972 30708 32978
rect 30656 32914 30708 32920
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 30472 32360 30524 32366
rect 30472 32302 30524 32308
rect 30484 31890 30512 32302
rect 30472 31884 30524 31890
rect 30472 31826 30524 31832
rect 30484 30802 30512 31826
rect 30668 31822 30696 32914
rect 30932 32904 30984 32910
rect 30932 32846 30984 32852
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30852 32026 30880 32370
rect 30840 32020 30892 32026
rect 30840 31962 30892 31968
rect 30944 31958 30972 32846
rect 31036 32774 31064 33238
rect 31024 32768 31076 32774
rect 31024 32710 31076 32716
rect 31036 32434 31064 32710
rect 31024 32428 31076 32434
rect 31024 32370 31076 32376
rect 30932 31952 30984 31958
rect 30932 31894 30984 31900
rect 30656 31816 30708 31822
rect 30656 31758 30708 31764
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30576 30938 30604 31282
rect 30564 30932 30616 30938
rect 30564 30874 30616 30880
rect 30944 30802 30972 31894
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30932 30796 30984 30802
rect 30932 30738 30984 30744
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30024 30394 30052 30670
rect 30012 30388 30064 30394
rect 30012 30330 30064 30336
rect 29644 29844 29696 29850
rect 29644 29786 29696 29792
rect 29828 29572 29880 29578
rect 29828 29514 29880 29520
rect 29552 28960 29604 28966
rect 29552 28902 29604 28908
rect 29564 28082 29592 28902
rect 29644 28756 29696 28762
rect 29644 28698 29696 28704
rect 29656 28558 29684 28698
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29656 27470 29684 28494
rect 29644 27464 29696 27470
rect 29696 27424 29776 27452
rect 29644 27406 29696 27412
rect 29644 27056 29696 27062
rect 29644 26998 29696 27004
rect 29656 26586 29684 26998
rect 29748 26926 29776 27424
rect 29736 26920 29788 26926
rect 29736 26862 29788 26868
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 29460 26444 29512 26450
rect 29460 26386 29512 26392
rect 29472 25294 29500 26386
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 29472 24410 29500 25230
rect 29564 24886 29592 26318
rect 29840 25906 29868 29514
rect 30288 29504 30340 29510
rect 30288 29446 30340 29452
rect 30012 28960 30064 28966
rect 30012 28902 30064 28908
rect 30024 28558 30052 28902
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 30104 28552 30156 28558
rect 30104 28494 30156 28500
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29932 27402 29960 28358
rect 30024 27402 30052 28494
rect 30116 27996 30144 28494
rect 30196 28212 30248 28218
rect 30196 28154 30248 28160
rect 30208 28121 30236 28154
rect 30300 28150 30328 29446
rect 30288 28144 30340 28150
rect 30194 28112 30250 28121
rect 30288 28086 30340 28092
rect 30194 28047 30250 28056
rect 30196 28008 30248 28014
rect 30116 27968 30196 27996
rect 30196 27950 30248 27956
rect 29920 27396 29972 27402
rect 29920 27338 29972 27344
rect 30012 27396 30064 27402
rect 30012 27338 30064 27344
rect 30208 27334 30236 27950
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 30300 26790 30328 28086
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 30392 27674 30420 28018
rect 30380 27668 30432 27674
rect 30380 27610 30432 27616
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 30484 26586 30512 30738
rect 30840 30184 30892 30190
rect 30840 30126 30892 30132
rect 30564 29776 30616 29782
rect 30564 29718 30616 29724
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30576 26382 30604 29718
rect 30852 29714 30880 30126
rect 30840 29708 30892 29714
rect 30840 29650 30892 29656
rect 30852 29578 30880 29650
rect 30840 29572 30892 29578
rect 30840 29514 30892 29520
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30668 29238 30696 29446
rect 30656 29232 30708 29238
rect 30656 29174 30708 29180
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30760 28966 30788 29106
rect 30748 28960 30800 28966
rect 30748 28902 30800 28908
rect 30852 27996 30880 29514
rect 30932 28144 30984 28150
rect 30930 28112 30932 28121
rect 30984 28112 30986 28121
rect 31036 28098 31064 31758
rect 31128 31346 31156 46990
rect 32232 46442 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 45626 32352 46446
rect 33784 46368 33836 46374
rect 33784 46310 33836 46316
rect 32312 45620 32364 45626
rect 32312 45562 32364 45568
rect 32128 45484 32180 45490
rect 32128 45426 32180 45432
rect 32140 43314 32168 45426
rect 32128 43308 32180 43314
rect 32128 43250 32180 43256
rect 32140 37874 32168 43250
rect 33796 42770 33824 46310
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 38028 45554 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38384 46640 38436 46646
rect 38384 46582 38436 46588
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38396 45966 38424 46582
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 39960 46374 39988 49200
rect 40788 47410 40816 49286
rect 41206 49200 41318 49286
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 41892 47546 41920 49200
rect 41892 47518 42012 47546
rect 40052 47382 40816 47410
rect 39948 46368 40000 46374
rect 39948 46310 40000 46316
rect 38200 45960 38252 45966
rect 38200 45902 38252 45908
rect 38384 45960 38436 45966
rect 38384 45902 38436 45908
rect 37292 45526 38056 45554
rect 37188 45348 37240 45354
rect 37188 45290 37240 45296
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 37200 44334 37228 45290
rect 37188 44328 37240 44334
rect 37188 44270 37240 44276
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 33784 42764 33836 42770
rect 33784 42706 33836 42712
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 32128 37868 32180 37874
rect 32128 37810 32180 37816
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 37292 35894 37320 45526
rect 37292 35866 37412 35894
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 31220 34610 31248 34886
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 31772 33998 31800 35022
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31668 33856 31720 33862
rect 31668 33798 31720 33804
rect 31944 33856 31996 33862
rect 31944 33798 31996 33804
rect 31576 32836 31628 32842
rect 31576 32778 31628 32784
rect 31588 32570 31616 32778
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31312 31754 31340 32370
rect 31312 31726 31524 31754
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 31312 30802 31340 31078
rect 31300 30796 31352 30802
rect 31300 30738 31352 30744
rect 31300 30592 31352 30598
rect 31300 30534 31352 30540
rect 31312 30258 31340 30534
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 31116 29640 31168 29646
rect 31116 29582 31168 29588
rect 31312 29594 31340 30194
rect 31392 29640 31444 29646
rect 31312 29588 31392 29594
rect 31312 29582 31444 29588
rect 31128 28762 31156 29582
rect 31312 29566 31432 29582
rect 31208 29504 31260 29510
rect 31208 29446 31260 29452
rect 31220 29170 31248 29446
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31116 28756 31168 28762
rect 31116 28698 31168 28704
rect 31208 28484 31260 28490
rect 31312 28472 31340 29566
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31260 28444 31340 28472
rect 31208 28426 31260 28432
rect 31036 28070 31156 28098
rect 30930 28047 30986 28056
rect 30932 28008 30984 28014
rect 30852 27968 30932 27996
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30576 25974 30604 26318
rect 30564 25968 30616 25974
rect 30564 25910 30616 25916
rect 30852 25906 30880 27968
rect 30932 27950 30984 27956
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 30944 26994 30972 27814
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 31128 26586 31156 28070
rect 31220 27878 31248 28426
rect 31404 28082 31432 28562
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 31208 27872 31260 27878
rect 31208 27814 31260 27820
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31312 27402 31340 27814
rect 31300 27396 31352 27402
rect 31300 27338 31352 27344
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 29828 25900 29880 25906
rect 29828 25842 29880 25848
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29552 24880 29604 24886
rect 29552 24822 29604 24828
rect 29460 24404 29512 24410
rect 29460 24346 29512 24352
rect 29656 23662 29684 25230
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29748 23730 29776 24754
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 29460 23656 29512 23662
rect 29460 23598 29512 23604
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29840 23610 29868 25842
rect 30852 25498 30880 25842
rect 30840 25492 30892 25498
rect 30840 25434 30892 25440
rect 30012 25424 30064 25430
rect 30012 25366 30064 25372
rect 29920 25152 29972 25158
rect 29920 25094 29972 25100
rect 29932 24274 29960 25094
rect 30024 24818 30052 25366
rect 30288 25220 30340 25226
rect 30288 25162 30340 25168
rect 30116 24818 30236 24834
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 30104 24812 30236 24818
rect 30156 24806 30236 24812
rect 30104 24754 30156 24760
rect 30024 24698 30052 24754
rect 30024 24670 30144 24698
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 29932 23798 29960 24210
rect 29920 23792 29972 23798
rect 29920 23734 29972 23740
rect 30024 23746 30052 24550
rect 30116 24206 30144 24670
rect 30208 24410 30236 24806
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30024 23718 30236 23746
rect 29472 23322 29500 23598
rect 29840 23582 30144 23610
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 29460 23316 29512 23322
rect 29460 23258 29512 23264
rect 29552 23044 29604 23050
rect 29552 22986 29604 22992
rect 29368 21004 29420 21010
rect 29368 20946 29420 20952
rect 29564 20466 29592 22986
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 29012 17134 29040 20334
rect 29920 18216 29972 18222
rect 29920 18158 29972 18164
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29012 16658 29040 17070
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 12434 29040 16594
rect 29012 12406 29132 12434
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 29012 3602 29040 9454
rect 29104 4078 29132 12406
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 29104 2990 29132 4014
rect 29196 3398 29224 4082
rect 29460 4072 29512 4078
rect 29458 4040 29460 4049
rect 29512 4040 29514 4049
rect 29458 3975 29514 3984
rect 29932 3738 29960 18158
rect 30024 12714 30052 23462
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 30116 8362 30144 23582
rect 30208 23526 30236 23718
rect 30196 23520 30248 23526
rect 30196 23462 30248 23468
rect 30300 23118 30328 25162
rect 31128 24750 31156 26522
rect 31496 25770 31524 31726
rect 31576 29504 31628 29510
rect 31576 29446 31628 29452
rect 31588 29306 31616 29446
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 31484 25764 31536 25770
rect 31484 25706 31536 25712
rect 31392 25696 31444 25702
rect 31392 25638 31444 25644
rect 31404 25498 31432 25638
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31496 25362 31524 25434
rect 31484 25356 31536 25362
rect 31484 25298 31536 25304
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 30668 24138 30696 24550
rect 31036 24410 31064 24550
rect 31128 24426 31156 24686
rect 31024 24404 31076 24410
rect 31128 24398 31248 24426
rect 31024 24346 31076 24352
rect 30932 24336 30984 24342
rect 30932 24278 30984 24284
rect 30656 24132 30708 24138
rect 30656 24074 30708 24080
rect 30944 23730 30972 24278
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 31128 23866 31156 24210
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 23186 30420 23462
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30668 23118 30696 23666
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 31220 23050 31248 24398
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 31404 23322 31432 23666
rect 31484 23520 31536 23526
rect 31484 23462 31536 23468
rect 31392 23316 31444 23322
rect 31392 23258 31444 23264
rect 31496 23254 31524 23462
rect 31484 23248 31536 23254
rect 31484 23190 31536 23196
rect 31208 23044 31260 23050
rect 31208 22986 31260 22992
rect 31392 20868 31444 20874
rect 31392 20810 31444 20816
rect 31404 20398 31432 20810
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30484 19922 30512 20198
rect 31404 19990 31432 20334
rect 31392 19984 31444 19990
rect 31392 19926 31444 19932
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30104 8356 30156 8362
rect 30104 8298 30156 8304
rect 31680 4078 31708 33798
rect 31956 32842 31984 33798
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 31944 32836 31996 32842
rect 31944 32778 31996 32784
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32324 30326 32352 30602
rect 32312 30320 32364 30326
rect 32312 30262 32364 30268
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 31852 29844 31904 29850
rect 31852 29786 31904 29792
rect 31864 28966 31892 29786
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32036 29028 32088 29034
rect 32036 28970 32088 28976
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 32048 28558 32076 28970
rect 32324 28626 32352 29242
rect 32588 29096 32640 29102
rect 32588 29038 32640 29044
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 32312 28620 32364 28626
rect 32312 28562 32364 28568
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32128 27532 32180 27538
rect 32128 27474 32180 27480
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 32036 26354 32088 26360
rect 31772 26042 31800 26318
rect 32036 26296 32088 26302
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 32048 25702 32076 26296
rect 32140 25838 32168 27474
rect 32324 26994 32352 28358
rect 32508 27946 32536 28494
rect 32496 27940 32548 27946
rect 32496 27882 32548 27888
rect 32600 27538 32628 29038
rect 32876 28762 32904 29038
rect 32864 28756 32916 28762
rect 32864 28698 32916 28704
rect 33336 28558 33364 30194
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 33416 29232 33468 29238
rect 33416 29174 33468 29180
rect 33428 28762 33456 29174
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33324 28552 33376 28558
rect 33324 28494 33376 28500
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32680 27940 32732 27946
rect 32680 27882 32732 27888
rect 32588 27532 32640 27538
rect 32588 27474 32640 27480
rect 32496 27396 32548 27402
rect 32496 27338 32548 27344
rect 32404 27328 32456 27334
rect 32404 27270 32456 27276
rect 32416 26994 32444 27270
rect 32508 27062 32536 27338
rect 32496 27056 32548 27062
rect 32496 26998 32548 27004
rect 32692 26994 32720 27882
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32324 26518 32352 26930
rect 32588 26920 32640 26926
rect 32588 26862 32640 26868
rect 32312 26512 32364 26518
rect 32312 26454 32364 26460
rect 32496 26240 32548 26246
rect 32496 26182 32548 26188
rect 32508 25974 32536 26182
rect 32496 25968 32548 25974
rect 32496 25910 32548 25916
rect 32128 25832 32180 25838
rect 32128 25774 32180 25780
rect 32036 25696 32088 25702
rect 32036 25638 32088 25644
rect 31852 25424 31904 25430
rect 31852 25366 31904 25372
rect 31864 25294 31892 25366
rect 32048 25362 32076 25638
rect 32036 25356 32088 25362
rect 32036 25298 32088 25304
rect 31852 25288 31904 25294
rect 31852 25230 31904 25236
rect 31864 24410 31892 25230
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 32140 24274 32168 25774
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32416 24138 32444 24550
rect 32404 24132 32456 24138
rect 32404 24074 32456 24080
rect 31944 19780 31996 19786
rect 31944 19722 31996 19728
rect 32128 19780 32180 19786
rect 32128 19722 32180 19728
rect 31956 19514 31984 19722
rect 31944 19508 31996 19514
rect 31944 19450 31996 19456
rect 31956 18970 31984 19450
rect 31944 18964 31996 18970
rect 31944 18906 31996 18912
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 27172 2746 27292 2774
rect 27632 2746 27752 2774
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 27172 2446 27200 2746
rect 27632 2582 27660 2746
rect 27620 2576 27672 2582
rect 27620 2518 27672 2524
rect 30024 2514 30052 4014
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 26436 800 26464 2314
rect 27080 800 27108 2314
rect 28368 800 28396 2314
rect 29656 800 29684 2382
rect 30944 800 30972 3538
rect 31312 3058 31340 4014
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 32140 2922 32168 19722
rect 32128 2916 32180 2922
rect 32128 2858 32180 2864
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 32232 800 32260 2790
rect 32600 2774 32628 26862
rect 32692 26382 32720 26930
rect 32680 26376 32732 26382
rect 32680 26318 32732 26324
rect 32784 25498 32812 28018
rect 33140 27872 33192 27878
rect 33140 27814 33192 27820
rect 33152 27402 33180 27814
rect 33140 27396 33192 27402
rect 33140 27338 33192 27344
rect 33336 26234 33364 28494
rect 36360 28076 36412 28082
rect 36360 28018 36412 28024
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 33152 26206 33364 26234
rect 32772 25492 32824 25498
rect 32772 25434 32824 25440
rect 33152 25294 33180 26206
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 33244 25498 33272 25910
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 33152 24818 33180 25230
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 36372 22982 36400 28018
rect 37280 28008 37332 28014
rect 37280 27950 37332 27956
rect 37292 27674 37320 27950
rect 37280 27668 37332 27674
rect 37280 27610 37332 27616
rect 36360 22976 36412 22982
rect 36360 22918 36412 22924
rect 37384 22710 37412 35866
rect 37372 22704 37424 22710
rect 37372 22646 37424 22652
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 38212 16182 38240 45902
rect 40052 24410 40080 47382
rect 41880 47048 41932 47054
rect 41880 46990 41932 46996
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40420 26450 40448 46922
rect 41892 46578 41920 46990
rect 41880 46572 41932 46578
rect 41880 46514 41932 46520
rect 41328 46368 41380 46374
rect 41328 46310 41380 46316
rect 41340 46034 41368 46310
rect 41984 46034 42012 47518
rect 42536 46442 42564 49200
rect 43180 47122 43208 49200
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 42616 47048 42668 47054
rect 42616 46990 42668 46996
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41328 46028 41380 46034
rect 41328 45970 41380 45976
rect 41972 46028 42024 46034
rect 41972 45970 42024 45976
rect 41512 45892 41564 45898
rect 41512 45834 41564 45840
rect 41524 45626 41552 45834
rect 41512 45620 41564 45626
rect 41512 45562 41564 45568
rect 42628 45082 42656 46990
rect 42892 46980 42944 46986
rect 42892 46922 42944 46928
rect 42904 45558 42932 46922
rect 43536 46368 43588 46374
rect 43536 46310 43588 46316
rect 42892 45552 42944 45558
rect 42892 45494 42944 45500
rect 42800 45484 42852 45490
rect 42800 45426 42852 45432
rect 42616 45076 42668 45082
rect 42616 45018 42668 45024
rect 42812 45014 42840 45426
rect 42800 45008 42852 45014
rect 42800 44950 42852 44956
rect 40408 26444 40460 26450
rect 40408 26386 40460 26392
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 42800 23112 42852 23118
rect 42800 23054 42852 23060
rect 40684 21956 40736 21962
rect 40684 21898 40736 21904
rect 40696 21622 40724 21898
rect 40684 21616 40736 21622
rect 40684 21558 40736 21564
rect 40684 20596 40736 20602
rect 40684 20538 40736 20544
rect 39304 20392 39356 20398
rect 39304 20334 39356 20340
rect 38200 16176 38252 16182
rect 38200 16118 38252 16124
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 32956 4276 33008 4282
rect 32956 4218 33008 4224
rect 32680 4208 32732 4214
rect 32680 4150 32732 4156
rect 32692 2990 32720 4150
rect 32772 3188 32824 3194
rect 32824 3148 32904 3176
rect 32772 3130 32824 3136
rect 32680 2984 32732 2990
rect 32680 2926 32732 2932
rect 32876 2922 32904 3148
rect 32968 3126 32996 4218
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 33152 3942 33180 4082
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 39120 3936 39172 3942
rect 39120 3878 39172 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 39028 3732 39080 3738
rect 39028 3674 39080 3680
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 33048 3052 33100 3058
rect 33244 3040 33272 3538
rect 35900 3528 35952 3534
rect 39040 3505 39068 3674
rect 39132 3534 39160 3878
rect 39224 3738 39252 4082
rect 39212 3732 39264 3738
rect 39212 3674 39264 3680
rect 39120 3528 39172 3534
rect 35900 3470 35952 3476
rect 39026 3496 39082 3505
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 33416 3120 33468 3126
rect 33416 3062 33468 3068
rect 33100 3012 33272 3040
rect 33048 2994 33100 3000
rect 33324 2984 33376 2990
rect 33428 2972 33456 3062
rect 33376 2944 33456 2972
rect 33508 2984 33560 2990
rect 33324 2926 33376 2932
rect 33508 2926 33560 2932
rect 32864 2916 32916 2922
rect 32864 2858 32916 2864
rect 32508 2746 32628 2774
rect 32508 2582 32536 2746
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35820 2446 35848 3402
rect 35912 2990 35940 3470
rect 36176 3460 36228 3466
rect 39120 3470 39172 3476
rect 39026 3431 39082 3440
rect 36176 3402 36228 3408
rect 36188 3194 36216 3402
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35808 2440 35860 2446
rect 35808 2382 35860 2388
rect 35452 800 35480 2382
rect 36096 800 36124 2994
rect 39316 2582 39344 20334
rect 40592 19712 40644 19718
rect 40592 19654 40644 19660
rect 40604 19514 40632 19654
rect 40592 19508 40644 19514
rect 40592 19450 40644 19456
rect 40696 19378 40724 20538
rect 42812 20466 42840 23054
rect 43444 22636 43496 22642
rect 43444 22578 43496 22584
rect 42800 20460 42852 20466
rect 42800 20402 42852 20408
rect 40776 19780 40828 19786
rect 40776 19722 40828 19728
rect 42432 19780 42484 19786
rect 42432 19722 42484 19728
rect 40788 19514 40816 19722
rect 40776 19508 40828 19514
rect 40776 19450 40828 19456
rect 40684 19372 40736 19378
rect 40684 19314 40736 19320
rect 40684 16516 40736 16522
rect 40684 16458 40736 16464
rect 40696 16114 40724 16458
rect 40684 16108 40736 16114
rect 40684 16050 40736 16056
rect 42444 12434 42472 19722
rect 43260 19440 43312 19446
rect 43260 19382 43312 19388
rect 43272 18766 43300 19382
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 42352 12406 42472 12434
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 39868 4282 39896 4558
rect 39948 4480 40000 4486
rect 39948 4422 40000 4428
rect 39856 4276 39908 4282
rect 39856 4218 39908 4224
rect 39580 4140 39632 4146
rect 39580 4082 39632 4088
rect 39592 3194 39620 4082
rect 39960 4026 39988 4422
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 39868 3998 39988 4026
rect 39868 3602 39896 3998
rect 40052 3602 40080 4150
rect 40960 4140 41012 4146
rect 40960 4082 41012 4088
rect 39856 3596 39908 3602
rect 39856 3538 39908 3544
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 40224 3596 40276 3602
rect 40224 3538 40276 3544
rect 40408 3596 40460 3602
rect 40408 3538 40460 3544
rect 40132 3460 40184 3466
rect 40132 3402 40184 3408
rect 39580 3188 39632 3194
rect 39580 3130 39632 3136
rect 39684 3058 39896 3074
rect 40144 3058 40172 3402
rect 39672 3052 39908 3058
rect 39724 3046 39856 3052
rect 39672 2994 39724 3000
rect 39856 2994 39908 3000
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 40236 2990 40264 3538
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 39304 2576 39356 2582
rect 39304 2518 39356 2524
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 38028 800 38056 2314
rect 39316 800 39344 2314
rect 39960 800 39988 2926
rect 40420 2854 40448 3538
rect 40498 3496 40554 3505
rect 40498 3431 40554 3440
rect 40512 2854 40540 3431
rect 40592 3052 40644 3058
rect 40592 2994 40644 3000
rect 40408 2848 40460 2854
rect 40408 2790 40460 2796
rect 40500 2848 40552 2854
rect 40500 2790 40552 2796
rect 40604 800 40632 2994
rect 40972 2378 41000 4082
rect 41052 4072 41104 4078
rect 41052 4014 41104 4020
rect 41328 4072 41380 4078
rect 41420 4072 41472 4078
rect 41380 4020 41420 4026
rect 41328 4014 41472 4020
rect 41064 3126 41092 4014
rect 41340 3998 41460 4014
rect 42352 3738 42380 12406
rect 42800 4480 42852 4486
rect 42800 4422 42852 4428
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 42616 3936 42668 3942
rect 42616 3878 42668 3884
rect 42340 3732 42392 3738
rect 42340 3674 42392 3680
rect 42248 3664 42300 3670
rect 42248 3606 42300 3612
rect 41420 3460 41472 3466
rect 41420 3402 41472 3408
rect 41432 3194 41460 3402
rect 41420 3188 41472 3194
rect 41420 3130 41472 3136
rect 41052 3120 41104 3126
rect 41052 3062 41104 3068
rect 41328 3120 41380 3126
rect 41328 3062 41380 3068
rect 41340 2446 41368 3062
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 40960 2372 41012 2378
rect 40960 2314 41012 2320
rect 41248 800 41276 2382
rect 42260 1714 42288 3606
rect 42444 3058 42472 3878
rect 42628 3602 42656 3878
rect 42812 3602 42840 4422
rect 43076 4276 43128 4282
rect 43076 4218 43128 4224
rect 43088 4078 43116 4218
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43456 3738 43484 22578
rect 43548 17270 43576 46310
rect 43824 45966 43852 49200
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 44088 45824 44140 45830
rect 44088 45766 44140 45772
rect 43996 45280 44048 45286
rect 43996 45222 44048 45228
rect 43720 40928 43772 40934
rect 43720 40870 43772 40876
rect 43732 22642 43760 40870
rect 44008 28626 44036 45222
rect 44100 28762 44128 45766
rect 44180 45554 44232 45558
rect 44468 45554 44496 49200
rect 45112 45626 45140 49200
rect 45192 47048 45244 47054
rect 45192 46990 45244 46996
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 44180 45552 44496 45554
rect 44232 45526 44496 45552
rect 44180 45494 44232 45500
rect 44456 45416 44508 45422
rect 44456 45358 44508 45364
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 44468 45082 44496 45358
rect 45112 45082 45140 45358
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 44916 44872 44968 44878
rect 44916 44814 44968 44820
rect 44180 33312 44232 33318
rect 44180 33254 44232 33260
rect 44192 32366 44220 33254
rect 44180 32360 44232 32366
rect 44180 32302 44232 32308
rect 44088 28756 44140 28762
rect 44088 28698 44140 28704
rect 43996 28620 44048 28626
rect 43996 28562 44048 28568
rect 43720 22636 43772 22642
rect 43720 22578 43772 22584
rect 44548 22568 44600 22574
rect 44548 22510 44600 22516
rect 44180 22024 44232 22030
rect 44180 21966 44232 21972
rect 43720 21888 43772 21894
rect 43720 21830 43772 21836
rect 43732 21554 43760 21830
rect 44192 21690 44220 21966
rect 44456 21888 44508 21894
rect 44456 21830 44508 21836
rect 44180 21684 44232 21690
rect 44180 21626 44232 21632
rect 43720 21548 43772 21554
rect 43720 21490 43772 21496
rect 43732 21146 43760 21490
rect 44192 21146 44220 21626
rect 44468 21554 44496 21830
rect 44560 21554 44588 22510
rect 44928 22094 44956 44814
rect 45204 44402 45232 46990
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45388 45558 45416 46922
rect 45756 45966 45784 49200
rect 46400 46918 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46388 46912 46440 46918
rect 46388 46854 46440 46860
rect 45928 46640 45980 46646
rect 45928 46582 45980 46588
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 45560 45824 45612 45830
rect 45848 45778 45876 45902
rect 45560 45766 45612 45772
rect 45376 45552 45428 45558
rect 45376 45494 45428 45500
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 45572 37330 45600 45766
rect 45756 45750 45876 45778
rect 45652 45620 45704 45626
rect 45652 45562 45704 45568
rect 45664 45422 45692 45562
rect 45652 45416 45704 45422
rect 45652 45358 45704 45364
rect 45652 44872 45704 44878
rect 45652 44814 45704 44820
rect 45664 44470 45692 44814
rect 45652 44464 45704 44470
rect 45652 44406 45704 44412
rect 45560 37324 45612 37330
rect 45560 37266 45612 37272
rect 45376 29708 45428 29714
rect 45376 29650 45428 29656
rect 45284 23588 45336 23594
rect 45284 23530 45336 23536
rect 45296 22098 45324 23530
rect 45388 22710 45416 29650
rect 45468 23588 45520 23594
rect 45468 23530 45520 23536
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 44652 22066 44956 22094
rect 45284 22092 45336 22098
rect 44456 21548 44508 21554
rect 44456 21490 44508 21496
rect 44548 21548 44600 21554
rect 44548 21490 44600 21496
rect 43720 21140 43772 21146
rect 43720 21082 43772 21088
rect 44180 21140 44232 21146
rect 44180 21082 44232 21088
rect 43904 20936 43956 20942
rect 44364 20936 44416 20942
rect 43904 20878 43956 20884
rect 44100 20884 44364 20890
rect 44100 20878 44416 20884
rect 43812 20256 43864 20262
rect 43812 20198 43864 20204
rect 43824 19854 43852 20198
rect 43812 19848 43864 19854
rect 43812 19790 43864 19796
rect 43916 19378 43944 20878
rect 44100 20862 44404 20878
rect 44100 19514 44128 20862
rect 44456 20800 44508 20806
rect 44456 20742 44508 20748
rect 44180 20392 44232 20398
rect 44180 20334 44232 20340
rect 44364 20392 44416 20398
rect 44364 20334 44416 20340
rect 44192 19990 44220 20334
rect 44180 19984 44232 19990
rect 44180 19926 44232 19932
rect 44088 19508 44140 19514
rect 44088 19450 44140 19456
rect 44100 19378 44128 19450
rect 44192 19378 44220 19926
rect 44376 19922 44404 20334
rect 44468 20330 44496 20742
rect 44456 20324 44508 20330
rect 44456 20266 44508 20272
rect 44468 19922 44496 20266
rect 44364 19916 44416 19922
rect 44364 19858 44416 19864
rect 44456 19916 44508 19922
rect 44456 19858 44508 19864
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 44088 19372 44140 19378
rect 44088 19314 44140 19320
rect 44180 19372 44232 19378
rect 44180 19314 44232 19320
rect 43536 17264 43588 17270
rect 43536 17206 43588 17212
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 43168 3596 43220 3602
rect 43168 3538 43220 3544
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42260 1686 42564 1714
rect 42536 800 42564 1686
rect 43180 800 43208 3538
rect 43456 3466 43484 3674
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 43548 3398 43576 17206
rect 43916 12434 43944 19314
rect 44272 19304 44324 19310
rect 44272 19246 44324 19252
rect 44180 19236 44232 19242
rect 44180 19178 44232 19184
rect 44192 18766 44220 19178
rect 44284 18970 44312 19246
rect 44272 18964 44324 18970
rect 44272 18906 44324 18912
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44192 18290 44220 18702
rect 44180 18284 44232 18290
rect 44180 18226 44232 18232
rect 44456 18216 44508 18222
rect 44456 18158 44508 18164
rect 44468 17882 44496 18158
rect 44456 17876 44508 17882
rect 44456 17818 44508 17824
rect 44652 17814 44680 22066
rect 45284 22034 45336 22040
rect 44916 22024 44968 22030
rect 44916 21966 44968 21972
rect 45376 22024 45428 22030
rect 45376 21966 45428 21972
rect 44928 21554 44956 21966
rect 45388 21865 45416 21966
rect 45374 21856 45430 21865
rect 45374 21791 45430 21800
rect 44916 21548 44968 21554
rect 44916 21490 44968 21496
rect 45376 21548 45428 21554
rect 45376 21490 45428 21496
rect 44732 20868 44784 20874
rect 44732 20810 44784 20816
rect 44640 17808 44692 17814
rect 44640 17750 44692 17756
rect 44088 17672 44140 17678
rect 44088 17614 44140 17620
rect 44272 17672 44324 17678
rect 44272 17614 44324 17620
rect 44100 17270 44128 17614
rect 44088 17264 44140 17270
rect 44088 17206 44140 17212
rect 44284 17202 44312 17614
rect 44272 17196 44324 17202
rect 44272 17138 44324 17144
rect 43824 12406 43944 12434
rect 43536 3392 43588 3398
rect 43536 3334 43588 3340
rect 43824 3194 43852 12406
rect 43904 4072 43956 4078
rect 43904 4014 43956 4020
rect 44088 4072 44140 4078
rect 44088 4014 44140 4020
rect 43812 3188 43864 3194
rect 43812 3130 43864 3136
rect 43916 2446 43944 4014
rect 44100 3738 44128 4014
rect 44088 3732 44140 3738
rect 44088 3674 44140 3680
rect 44744 3670 44772 20810
rect 45388 19922 45416 21490
rect 45480 20534 45508 23530
rect 45560 23112 45612 23118
rect 45560 23054 45612 23060
rect 45572 22574 45600 23054
rect 45560 22568 45612 22574
rect 45560 22510 45612 22516
rect 45468 20528 45520 20534
rect 45468 20470 45520 20476
rect 45376 19916 45428 19922
rect 45376 19858 45428 19864
rect 44824 19848 44876 19854
rect 44824 19790 44876 19796
rect 44836 18154 44864 19790
rect 45008 19372 45060 19378
rect 45008 19314 45060 19320
rect 44916 18760 44968 18766
rect 44916 18702 44968 18708
rect 44928 18290 44956 18702
rect 45020 18358 45048 19314
rect 45572 19310 45600 22510
rect 45664 21978 45692 44406
rect 45756 44402 45784 45750
rect 45940 45554 45968 46582
rect 46860 46510 46888 47631
rect 46296 46504 46348 46510
rect 46296 46446 46348 46452
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 45848 45526 45968 45554
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 45848 41138 45876 45526
rect 46308 44538 46336 46446
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 47860 47184 47912 47190
rect 47860 47126 47912 47132
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47124 46912 47176 46918
rect 47124 46854 47176 46860
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46492 45082 46520 45834
rect 47136 45558 47164 46854
rect 47768 46436 47820 46442
rect 47768 46378 47820 46384
rect 47124 45552 47176 45558
rect 47124 45494 47176 45500
rect 46664 45484 46716 45490
rect 46664 45426 46716 45432
rect 46676 45354 46704 45426
rect 46664 45348 46716 45354
rect 46664 45290 46716 45296
rect 46480 45076 46532 45082
rect 46480 45018 46532 45024
rect 46296 44532 46348 44538
rect 46296 44474 46348 44480
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 45836 41132 45888 41138
rect 45836 41074 45888 41080
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46112 38956 46164 38962
rect 46112 38898 46164 38904
rect 45836 33856 45888 33862
rect 45836 33798 45888 33804
rect 45742 28656 45798 28665
rect 45742 28591 45798 28600
rect 45756 22098 45784 28591
rect 45744 22092 45796 22098
rect 45744 22034 45796 22040
rect 45664 21950 45784 21978
rect 45756 20534 45784 21950
rect 45744 20528 45796 20534
rect 45744 20470 45796 20476
rect 45848 19514 45876 33798
rect 46124 24750 46152 38898
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46308 37466 46336 38286
rect 46296 37460 46348 37466
rect 46296 37402 46348 37408
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 32434 46336 32846
rect 46296 32428 46348 32434
rect 46296 32370 46348 32376
rect 46676 32366 46704 45290
rect 47216 45280 47268 45286
rect 47216 45222 47268 45228
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 46940 44804 46992 44810
rect 46940 44746 46992 44752
rect 46952 44538 46980 44746
rect 46940 44532 46992 44538
rect 46940 44474 46992 44480
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 46754 39536 46810 39545
rect 46754 39471 46810 39480
rect 46664 32360 46716 32366
rect 46664 32302 46716 32308
rect 46386 31376 46442 31385
rect 46386 31311 46442 31320
rect 46296 25696 46348 25702
rect 46296 25638 46348 25644
rect 46308 25362 46336 25638
rect 46296 25356 46348 25362
rect 46296 25298 46348 25304
rect 45928 24744 45980 24750
rect 45928 24686 45980 24692
rect 46112 24744 46164 24750
rect 46112 24686 46164 24692
rect 45940 20602 45968 24686
rect 46296 24200 46348 24206
rect 46296 24142 46348 24148
rect 46308 23730 46336 24142
rect 46296 23724 46348 23730
rect 46296 23666 46348 23672
rect 46204 23656 46256 23662
rect 46204 23598 46256 23604
rect 46216 23225 46244 23598
rect 46202 23216 46258 23225
rect 46202 23151 46258 23160
rect 46020 22024 46072 22030
rect 46020 21966 46072 21972
rect 46032 21418 46060 21966
rect 46020 21412 46072 21418
rect 46020 21354 46072 21360
rect 45928 20596 45980 20602
rect 45928 20538 45980 20544
rect 45836 19508 45888 19514
rect 45836 19450 45888 19456
rect 45940 19394 45968 20538
rect 45756 19366 45968 19394
rect 45560 19304 45612 19310
rect 45560 19246 45612 19252
rect 45192 18760 45244 18766
rect 45192 18702 45244 18708
rect 45100 18692 45152 18698
rect 45100 18634 45152 18640
rect 45008 18352 45060 18358
rect 45008 18294 45060 18300
rect 44916 18284 44968 18290
rect 44916 18226 44968 18232
rect 44824 18148 44876 18154
rect 44824 18090 44876 18096
rect 44928 17882 44956 18226
rect 45112 18086 45140 18634
rect 45100 18080 45152 18086
rect 45100 18022 45152 18028
rect 44916 17876 44968 17882
rect 44916 17818 44968 17824
rect 45112 17678 45140 18022
rect 45100 17672 45152 17678
rect 45100 17614 45152 17620
rect 45204 17610 45232 18702
rect 45192 17604 45244 17610
rect 45192 17546 45244 17552
rect 45204 7342 45232 17546
rect 45558 15736 45614 15745
rect 45558 15671 45614 15680
rect 45572 15570 45600 15671
rect 45560 15564 45612 15570
rect 45560 15506 45612 15512
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 45192 7336 45244 7342
rect 45192 7278 45244 7284
rect 45204 5098 45232 7278
rect 45192 5092 45244 5098
rect 45192 5034 45244 5040
rect 45192 4616 45244 4622
rect 45192 4558 45244 4564
rect 44732 3664 44784 3670
rect 44732 3606 44784 3612
rect 45204 3058 45232 4558
rect 45756 4146 45784 19366
rect 45928 18284 45980 18290
rect 45928 18226 45980 18232
rect 45940 17338 45968 18226
rect 45928 17332 45980 17338
rect 45928 17274 45980 17280
rect 46032 7954 46060 21354
rect 46296 20936 46348 20942
rect 46296 20878 46348 20884
rect 46308 19310 46336 20878
rect 46296 19304 46348 19310
rect 46296 19246 46348 19252
rect 46296 19168 46348 19174
rect 46296 19110 46348 19116
rect 46308 18834 46336 19110
rect 46296 18828 46348 18834
rect 46296 18770 46348 18776
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 17202 46336 17614
rect 46296 17196 46348 17202
rect 46296 17138 46348 17144
rect 46400 16250 46428 31311
rect 46570 30016 46626 30025
rect 46570 29951 46626 29960
rect 46584 27130 46612 29951
rect 46572 27124 46624 27130
rect 46572 27066 46624 27072
rect 46570 26616 46626 26625
rect 46570 26551 46626 26560
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46584 22658 46612 26551
rect 46768 26234 46796 39471
rect 46940 39364 46992 39370
rect 46940 39306 46992 39312
rect 46952 39098 46980 39306
rect 46940 39092 46992 39098
rect 46940 39034 46992 39040
rect 46848 28008 46900 28014
rect 46846 27976 46848 27985
rect 46900 27976 46902 27985
rect 46846 27911 46902 27920
rect 46492 22630 46612 22658
rect 46676 26206 46796 26234
rect 46492 19666 46520 22630
rect 46572 22568 46624 22574
rect 46572 22510 46624 22516
rect 46584 20398 46612 22510
rect 46676 22386 46704 26206
rect 46846 25936 46902 25945
rect 46846 25871 46902 25880
rect 46756 24812 46808 24818
rect 46756 24754 46808 24760
rect 46768 23905 46796 24754
rect 46754 23896 46810 23905
rect 46754 23831 46810 23840
rect 46860 23186 46888 25871
rect 46756 23180 46808 23186
rect 46756 23122 46808 23128
rect 46848 23180 46900 23186
rect 46848 23122 46900 23128
rect 46768 22545 46796 23122
rect 46754 22536 46810 22545
rect 46754 22471 46810 22480
rect 46676 22358 46888 22386
rect 46860 22250 46888 22358
rect 46860 22222 46980 22250
rect 46848 22094 46900 22098
rect 46952 22094 46980 22222
rect 46848 22092 46980 22094
rect 46900 22066 46980 22092
rect 46848 22034 46900 22040
rect 47228 21010 47256 45222
rect 47400 45008 47452 45014
rect 47400 44950 47452 44956
rect 47412 42226 47440 44950
rect 47676 44192 47728 44198
rect 47676 44134 47728 44140
rect 47688 43858 47716 44134
rect 47676 43852 47728 43858
rect 47676 43794 47728 43800
rect 47780 43314 47808 46378
rect 47768 43308 47820 43314
rect 47768 43250 47820 43256
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47400 42220 47452 42226
rect 47400 42162 47452 42168
rect 47308 35080 47360 35086
rect 47308 35022 47360 35028
rect 47320 34105 47348 35022
rect 47306 34096 47362 34105
rect 47306 34031 47362 34040
rect 47306 32056 47362 32065
rect 47306 31991 47362 32000
rect 47320 31890 47348 31991
rect 47308 31884 47360 31890
rect 47308 31826 47360 31832
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47320 29345 47348 29582
rect 47306 29336 47362 29345
rect 47306 29271 47362 29280
rect 47216 21004 47268 21010
rect 47216 20946 47268 20952
rect 46940 20460 46992 20466
rect 46940 20402 46992 20408
rect 46572 20392 46624 20398
rect 46572 20334 46624 20340
rect 46492 19638 46704 19666
rect 46480 19508 46532 19514
rect 46480 19450 46532 19456
rect 46388 16244 46440 16250
rect 46388 16186 46440 16192
rect 46492 12434 46520 19450
rect 46572 17128 46624 17134
rect 46572 17070 46624 17076
rect 46400 12406 46520 12434
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46202 9616 46258 9625
rect 46202 9551 46204 9560
rect 46256 9551 46258 9560
rect 46204 9522 46256 9528
rect 46400 9110 46428 12406
rect 46480 11076 46532 11082
rect 46480 11018 46532 11024
rect 46492 10810 46520 11018
rect 46480 10804 46532 10810
rect 46480 10746 46532 10752
rect 46480 9512 46532 9518
rect 46480 9454 46532 9460
rect 46388 9104 46440 9110
rect 46388 9046 46440 9052
rect 46492 9042 46520 9454
rect 46480 9036 46532 9042
rect 46480 8978 46532 8984
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 46020 7948 46072 7954
rect 46020 7890 46072 7896
rect 46308 5370 46336 8910
rect 46584 5710 46612 17070
rect 46676 17066 46704 19638
rect 46846 18456 46902 18465
rect 46846 18391 46902 18400
rect 46860 18290 46888 18391
rect 46848 18284 46900 18290
rect 46848 18226 46900 18232
rect 46664 17060 46716 17066
rect 46664 17002 46716 17008
rect 46756 16516 46808 16522
rect 46756 16458 46808 16464
rect 46768 16250 46796 16458
rect 46756 16244 46808 16250
rect 46756 16186 46808 16192
rect 46952 15706 46980 20402
rect 47412 18290 47440 42162
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 40730 47716 41618
rect 47676 40724 47728 40730
rect 47676 40666 47728 40672
rect 47768 38956 47820 38962
rect 47768 38898 47820 38904
rect 47780 38865 47808 38898
rect 47766 38856 47822 38865
rect 47766 38791 47822 38800
rect 47768 38752 47820 38758
rect 47768 38694 47820 38700
rect 47676 38276 47728 38282
rect 47676 38218 47728 38224
rect 47688 38010 47716 38218
rect 47676 38004 47728 38010
rect 47676 37946 47728 37952
rect 47492 35080 47544 35086
rect 47492 35022 47544 35028
rect 47504 33930 47532 35022
rect 47492 33924 47544 33930
rect 47492 33866 47544 33872
rect 47676 32836 47728 32842
rect 47676 32778 47728 32784
rect 47688 32570 47716 32778
rect 47676 32564 47728 32570
rect 47676 32506 47728 32512
rect 47492 32496 47544 32502
rect 47492 32438 47544 32444
rect 47504 31890 47532 32438
rect 47492 31884 47544 31890
rect 47492 31826 47544 31832
rect 47676 25220 47728 25226
rect 47676 25162 47728 25168
rect 47688 24818 47716 25162
rect 47492 24812 47544 24818
rect 47492 24754 47544 24760
rect 47676 24812 47728 24818
rect 47676 24754 47728 24760
rect 47400 18284 47452 18290
rect 47400 18226 47452 18232
rect 47400 17808 47452 17814
rect 47400 17750 47452 17756
rect 47412 17202 47440 17750
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 46940 15700 46992 15706
rect 46940 15642 46992 15648
rect 46846 6216 46902 6225
rect 46846 6151 46902 6160
rect 46860 5778 46888 6151
rect 46848 5772 46900 5778
rect 46848 5714 46900 5720
rect 46572 5704 46624 5710
rect 46572 5646 46624 5652
rect 45836 5364 45888 5370
rect 45836 5306 45888 5312
rect 46296 5364 46348 5370
rect 46296 5306 46348 5312
rect 45848 4690 45876 5306
rect 46848 5228 46900 5234
rect 46848 5170 46900 5176
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45848 4282 45876 4626
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45836 4276 45888 4282
rect 45836 4218 45888 4224
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45100 2848 45152 2854
rect 45100 2790 45152 2796
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 43824 800 43852 2382
rect 45112 800 45140 2790
rect 46032 2446 46060 4490
rect 46664 4208 46716 4214
rect 46664 4150 46716 4156
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46492 3602 46520 3878
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46676 3505 46704 4150
rect 46662 3496 46718 3505
rect 46662 3431 46718 3440
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 46020 2440 46072 2446
rect 46020 2382 46072 2388
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 46400 800 46428 2314
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46768 105 46796 2994
rect 46860 921 46888 5170
rect 46952 4758 46980 15642
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47320 6866 47348 7511
rect 47308 6860 47360 6866
rect 47308 6802 47360 6808
rect 46940 4752 46992 4758
rect 46940 4694 46992 4700
rect 47032 4684 47084 4690
rect 47032 4626 47084 4632
rect 47044 3670 47072 4626
rect 47032 3664 47084 3670
rect 47032 3606 47084 3612
rect 47412 3466 47440 17138
rect 47504 16726 47532 24754
rect 47780 23866 47808 38694
rect 47872 33674 47900 47126
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47952 46572 48004 46578
rect 47952 46514 48004 46520
rect 47964 46345 47992 46514
rect 48044 46368 48096 46374
rect 47950 46336 48006 46345
rect 48044 46310 48096 46316
rect 47950 46271 48006 46280
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47964 40905 47992 41074
rect 47950 40896 48006 40905
rect 47950 40831 48006 40840
rect 47952 34400 48004 34406
rect 47952 34342 48004 34348
rect 47964 34066 47992 34342
rect 47952 34060 48004 34066
rect 47952 34002 48004 34008
rect 47872 33646 47992 33674
rect 47860 33516 47912 33522
rect 47860 33458 47912 33464
rect 47872 33425 47900 33458
rect 47858 33416 47914 33425
rect 47858 33351 47914 33360
rect 47964 30122 47992 33646
rect 47952 30116 48004 30122
rect 47952 30058 48004 30064
rect 47768 23860 47820 23866
rect 47768 23802 47820 23808
rect 47676 23044 47728 23050
rect 47676 22986 47728 22992
rect 47688 22778 47716 22986
rect 47676 22772 47728 22778
rect 47676 22714 47728 22720
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47596 21554 47624 22578
rect 47676 21956 47728 21962
rect 47676 21898 47728 21904
rect 47688 21690 47716 21898
rect 47676 21684 47728 21690
rect 47676 21626 47728 21632
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47596 19446 47624 21490
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 20602 47716 20810
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 47952 20392 48004 20398
rect 47952 20334 48004 20340
rect 47964 19802 47992 20334
rect 48056 19922 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48148 34610 48176 34711
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48134 25256 48190 25265
rect 48134 25191 48136 25200
rect 48188 25191 48190 25200
rect 48136 25162 48188 25168
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48044 19916 48096 19922
rect 48044 19858 48096 19864
rect 47964 19786 48084 19802
rect 47964 19780 48096 19786
rect 47964 19774 48044 19780
rect 48044 19722 48096 19728
rect 47584 19440 47636 19446
rect 47584 19382 47636 19388
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47676 17604 47728 17610
rect 47676 17546 47728 17552
rect 47688 17338 47716 17546
rect 47676 17332 47728 17338
rect 47676 17274 47728 17280
rect 47492 16720 47544 16726
rect 47492 16662 47544 16668
rect 47504 9586 47532 16662
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47780 16114 47808 16594
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47768 12640 47820 12646
rect 47768 12582 47820 12588
rect 47780 12306 47808 12582
rect 47768 12300 47820 12306
rect 47768 12242 47820 12248
rect 47676 12164 47728 12170
rect 47676 12106 47728 12112
rect 47688 11898 47716 12106
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47768 11212 47820 11218
rect 47768 11154 47820 11160
rect 47780 10674 47808 11154
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47492 9580 47544 9586
rect 47492 9522 47544 9528
rect 47766 8936 47822 8945
rect 47766 8871 47822 8880
rect 47780 8566 47808 8871
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 48056 7954 48084 19722
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48136 17604 48188 17610
rect 48136 17546 48188 17552
rect 48148 17105 48176 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48136 16516 48188 16522
rect 48136 16458 48188 16464
rect 48148 16425 48176 16458
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48134 12336 48190 12345
rect 48134 12271 48136 12280
rect 48188 12271 48190 12280
rect 48136 12242 48188 12248
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48044 7948 48096 7954
rect 48044 7890 48096 7896
rect 47492 7812 47544 7818
rect 47492 7754 47544 7760
rect 47504 6866 47532 7754
rect 47492 6860 47544 6866
rect 47492 6802 47544 6808
rect 47952 6112 48004 6118
rect 47952 6054 48004 6060
rect 47964 5302 47992 6054
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 47768 4208 47820 4214
rect 47768 4150 47820 4156
rect 47400 3460 47452 3466
rect 47400 3402 47452 3408
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 46846 912 46902 921
rect 46846 847 46902 856
rect 47044 800 47072 2450
rect 47688 800 47716 2926
rect 47780 1465 47808 4150
rect 48056 3194 48084 7890
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48134 6831 48190 6840
rect 48136 6316 48188 6322
rect 48136 6258 48188 6264
rect 48148 4185 48176 6258
rect 48134 4176 48190 4185
rect 48134 4111 48190 4120
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 48320 2372 48372 2378
rect 48320 2314 48372 2320
rect 47766 1456 47822 1465
rect 47766 1391 47822 1400
rect 48332 800 48360 2314
rect 48976 800 49004 3402
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1858 47640 1914 47696
rect 3422 46960 3478 47016
rect 1858 42880 1914 42936
rect 1858 41520 1914 41576
rect 1858 40160 1914 40216
rect 1582 35400 1638 35456
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 32680 1638 32736
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1398 12280 1454 12336
rect 1858 23160 1914 23216
rect 1950 20440 2006 20496
rect 2226 19080 2282 19136
rect 3054 46280 3110 46336
rect 2778 36760 2834 36816
rect 2778 32000 2834 32056
rect 1858 17720 1914 17776
rect 2778 16360 2834 16416
rect 3238 19896 3294 19952
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3514 44920 3570 44976
rect 3698 43560 3754 43616
rect 3606 39480 3662 39536
rect 3790 31320 3846 31376
rect 3974 28600 4030 28656
rect 3974 19760 4030 19816
rect 3974 18400 4030 18456
rect 3974 17040 4030 17096
rect 2778 15000 2834 15056
rect 3790 13676 3792 13696
rect 3792 13676 3844 13696
rect 3844 13676 3846 13696
rect 3790 13640 3846 13676
rect 2778 10240 2834 10296
rect 3146 7520 3202 7576
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3974 3984 4030 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3606 3440 3662 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3330 1400 3386 1456
rect 16670 32428 16726 32464
rect 16670 32408 16672 32428
rect 16672 32408 16724 32428
rect 16724 32408 16726 32428
rect 17406 32444 17408 32464
rect 17408 32444 17460 32464
rect 17460 32444 17462 32464
rect 17406 32408 17462 32444
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19338 33496 19394 33552
rect 17682 13948 17684 13968
rect 17684 13948 17736 13968
rect 17736 13948 17738 13968
rect 17682 13912 17738 13948
rect 18786 13948 18788 13968
rect 18788 13948 18840 13968
rect 18840 13948 18842 13968
rect 18786 13912 18842 13948
rect 17682 2760 17738 2816
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20074 21004 20130 21040
rect 20074 20984 20076 21004
rect 20076 20984 20128 21004
rect 20128 20984 20130 21004
rect 20350 28872 20406 28928
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19246 3032 19302 3088
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19890 2932 19892 2952
rect 19892 2932 19944 2952
rect 19944 2932 19946 2952
rect 19890 2896 19946 2932
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21546 29044 21548 29064
rect 21548 29044 21600 29064
rect 21600 29044 21602 29064
rect 21546 29008 21602 29044
rect 22190 33516 22246 33552
rect 22190 33496 22192 33516
rect 22192 33496 22244 33516
rect 22244 33496 22246 33516
rect 23018 31592 23074 31648
rect 21730 4156 21732 4176
rect 21732 4156 21784 4176
rect 21784 4156 21786 4176
rect 21730 4120 21786 4156
rect 21914 3440 21970 3496
rect 21454 3304 21510 3360
rect 22098 3576 22154 3632
rect 22650 3460 22706 3496
rect 22650 3440 22652 3460
rect 22652 3440 22704 3460
rect 22704 3440 22706 3460
rect 23386 3440 23442 3496
rect 22282 3068 22284 3088
rect 22284 3068 22336 3088
rect 22336 3068 22338 3088
rect 22282 3032 22338 3068
rect 21362 2760 21418 2816
rect 24030 24948 24086 24984
rect 24030 24928 24032 24948
rect 24032 24928 24084 24948
rect 24084 24928 24086 24948
rect 24306 24656 24362 24712
rect 25226 29996 25228 30016
rect 25228 29996 25280 30016
rect 25280 29996 25282 30016
rect 25226 29960 25282 29996
rect 24950 29008 25006 29064
rect 24858 24828 24860 24848
rect 24860 24828 24912 24848
rect 24912 24828 24914 24848
rect 24858 24792 24914 24828
rect 25226 24928 25282 24984
rect 25226 24656 25282 24712
rect 26054 29008 26110 29064
rect 24858 3576 24914 3632
rect 24858 2896 24914 2952
rect 26238 24812 26294 24848
rect 26238 24792 26240 24812
rect 26240 24792 26292 24812
rect 26292 24792 26294 24812
rect 26606 21004 26662 21040
rect 26606 20984 26608 21004
rect 26608 20984 26660 21004
rect 26660 20984 26662 21004
rect 25318 3460 25374 3496
rect 25318 3440 25320 3460
rect 25320 3440 25372 3460
rect 25372 3440 25374 3460
rect 28998 34040 29054 34096
rect 29274 33924 29330 33960
rect 29274 33904 29276 33924
rect 29276 33904 29328 33924
rect 29328 33904 29330 33924
rect 29182 33768 29238 33824
rect 28538 33496 28594 33552
rect 27342 29960 27398 30016
rect 27986 31592 28042 31648
rect 27158 15564 27214 15600
rect 27158 15544 27160 15564
rect 27160 15544 27212 15564
rect 27212 15544 27214 15564
rect 26974 4120 27030 4176
rect 27618 3304 27674 3360
rect 28262 28872 28318 28928
rect 27802 20476 27804 20496
rect 27804 20476 27856 20496
rect 27856 20476 27858 20496
rect 27802 20440 27858 20476
rect 27802 19916 27858 19952
rect 27802 19896 27804 19916
rect 27804 19896 27856 19916
rect 27856 19896 27858 19916
rect 29458 33380 29514 33416
rect 29458 33360 29460 33380
rect 29460 33360 29512 33380
rect 29512 33360 29514 33380
rect 29734 33940 29736 33960
rect 29736 33940 29788 33960
rect 29788 33940 29790 33960
rect 29734 33904 29790 33940
rect 30102 34040 30158 34096
rect 30378 33380 30434 33416
rect 30378 33360 30380 33380
rect 30380 33360 30432 33380
rect 30432 33360 30434 33380
rect 30746 33768 30802 33824
rect 30194 28056 30250 28112
rect 30930 28092 30932 28112
rect 30932 28092 30984 28112
rect 30984 28092 30986 28112
rect 30930 28056 30986 28092
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 29458 4020 29460 4040
rect 29460 4020 29512 4040
rect 29512 4020 29514 4040
rect 29458 3984 29514 4020
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39026 3440 39082 3496
rect 40498 3440 40554 3496
rect 46846 47640 46902 47696
rect 45374 21800 45430 21856
rect 45742 28600 45798 28656
rect 46754 39480 46810 39536
rect 46386 31320 46442 31376
rect 46202 23160 46258 23216
rect 45558 15680 45614 15736
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 46570 29960 46626 30016
rect 46570 26560 46626 26616
rect 46846 27956 46848 27976
rect 46848 27956 46900 27976
rect 46900 27956 46902 27976
rect 46846 27920 46902 27956
rect 46846 25880 46902 25936
rect 46754 23840 46810 23896
rect 46754 22480 46810 22536
rect 47306 34040 47362 34096
rect 47306 32000 47362 32056
rect 47306 29280 47362 29336
rect 46202 9580 46258 9616
rect 46202 9560 46204 9580
rect 46204 9560 46256 9580
rect 46256 9560 46258 9580
rect 46846 18400 46902 18456
rect 47766 38800 47822 38856
rect 46846 6160 46902 6216
rect 46662 3440 46718 3496
rect 2962 720 3018 776
rect 47306 7520 47362 7576
rect 47950 46280 48006 46336
rect 47950 40840 48006 40896
rect 47858 33360 47914 33416
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48134 32680 48190 32736
rect 48134 25220 48190 25256
rect 48134 25200 48136 25220
rect 48136 25200 48188 25220
rect 48188 25200 48190 25220
rect 48134 24520 48190 24576
rect 48134 21120 48190 21176
rect 47766 8880 47822 8936
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 12300 48190 12336
rect 48134 12280 48136 12300
rect 48136 12280 48188 12300
rect 48188 12280 48190 12300
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 46846 856 46902 912
rect 48134 6840 48190 6896
rect 48134 4120 48190 4176
rect 47766 1400 47822 1456
rect 46754 40 46810 96
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1853 47698 1919 47701
rect 0 47696 1919 47698
rect 0 47640 1858 47696
rect 1914 47640 1919 47696
rect 0 47638 1919 47640
rect 0 47548 800 47638
rect 1853 47635 1919 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3417 47018 3483 47021
rect 0 47016 3483 47018
rect 0 46960 3422 47016
rect 3478 46960 3483 47016
rect 0 46958 3483 46960
rect 0 46868 800 46958
rect 3417 46955 3483 46958
rect 46054 46956 46060 47020
rect 46124 47018 46130 47020
rect 49200 47018 50000 47108
rect 46124 46958 50000 47018
rect 46124 46956 46130 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 3049 46338 3115 46341
rect 0 46336 3115 46338
rect 0 46280 3054 46336
rect 3110 46280 3115 46336
rect 0 46278 3115 46280
rect 0 46188 800 46278
rect 3049 46275 3115 46278
rect 47945 46338 48011 46341
rect 49200 46338 50000 46428
rect 47945 46336 50000 46338
rect 47945 46280 47950 46336
rect 48006 46280 50000 46336
rect 47945 46278 50000 46280
rect 47945 46275 48011 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3509 44978 3575 44981
rect 0 44976 3575 44978
rect 0 44920 3514 44976
rect 3570 44920 3575 44976
rect 0 44918 3575 44920
rect 0 44828 800 44918
rect 3509 44915 3575 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3693 43618 3759 43621
rect 0 43616 3759 43618
rect 0 43560 3698 43616
rect 3754 43560 3759 43616
rect 0 43558 3759 43560
rect 0 43468 800 43558
rect 3693 43555 3759 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1853 42938 1919 42941
rect 0 42936 1919 42938
rect 0 42880 1858 42936
rect 1914 42880 1919 42936
rect 0 42878 1919 42880
rect 0 42788 800 42878
rect 1853 42875 1919 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 47945 40898 48011 40901
rect 49200 40898 50000 40988
rect 47945 40896 50000 40898
rect 47945 40840 47950 40896
rect 48006 40840 50000 40896
rect 47945 40838 50000 40840
rect 47945 40835 48011 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40068 800 40158
rect 1853 40155 1919 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3601 39538 3667 39541
rect 0 39536 3667 39538
rect 0 39480 3606 39536
rect 3662 39480 3667 39536
rect 0 39478 3667 39480
rect 0 39388 800 39478
rect 3601 39475 3667 39478
rect 46749 39538 46815 39541
rect 49200 39538 50000 39628
rect 46749 39536 50000 39538
rect 46749 39480 46754 39536
rect 46810 39480 50000 39536
rect 46749 39478 50000 39480
rect 46749 39475 46815 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47761 38858 47827 38861
rect 49200 38858 50000 38948
rect 47761 38856 50000 38858
rect 47761 38800 47766 38856
rect 47822 38800 50000 38856
rect 47761 38798 50000 38800
rect 47761 38795 47827 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 28993 34098 29059 34101
rect 30097 34098 30163 34101
rect 28993 34096 30163 34098
rect 28993 34040 28998 34096
rect 29054 34040 30102 34096
rect 30158 34040 30163 34096
rect 28993 34038 30163 34040
rect 28993 34035 29059 34038
rect 30097 34035 30163 34038
rect 47301 34098 47367 34101
rect 49200 34098 50000 34188
rect 47301 34096 50000 34098
rect 47301 34040 47306 34096
rect 47362 34040 50000 34096
rect 47301 34038 50000 34040
rect 47301 34035 47367 34038
rect 29269 33962 29335 33965
rect 29729 33962 29795 33965
rect 29269 33960 29795 33962
rect 29269 33904 29274 33960
rect 29330 33904 29734 33960
rect 29790 33904 29795 33960
rect 49200 33948 50000 34038
rect 29269 33902 29795 33904
rect 29269 33899 29335 33902
rect 29729 33899 29795 33902
rect 29177 33826 29243 33829
rect 30741 33826 30807 33829
rect 29177 33824 30807 33826
rect 29177 33768 29182 33824
rect 29238 33768 30746 33824
rect 30802 33768 30807 33824
rect 29177 33766 30807 33768
rect 29177 33763 29243 33766
rect 30741 33763 30807 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 19333 33554 19399 33557
rect 22185 33554 22251 33557
rect 28533 33554 28599 33557
rect 19333 33552 28599 33554
rect 0 33418 800 33508
rect 19333 33496 19338 33552
rect 19394 33496 22190 33552
rect 22246 33496 28538 33552
rect 28594 33496 28599 33552
rect 19333 33494 28599 33496
rect 19333 33491 19399 33494
rect 22185 33491 22251 33494
rect 28533 33491 28599 33494
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 29453 33418 29519 33421
rect 30373 33418 30439 33421
rect 29453 33416 30439 33418
rect 29453 33360 29458 33416
rect 29514 33360 30378 33416
rect 30434 33360 30439 33416
rect 29453 33358 30439 33360
rect 29453 33355 29519 33358
rect 30373 33355 30439 33358
rect 47853 33418 47919 33421
rect 49200 33418 50000 33508
rect 47853 33416 50000 33418
rect 47853 33360 47858 33416
rect 47914 33360 50000 33416
rect 47853 33358 50000 33360
rect 47853 33355 47919 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32828
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32588 800 32678
rect 1577 32675 1643 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 16665 32466 16731 32469
rect 17401 32466 17467 32469
rect 16665 32464 17467 32466
rect 16665 32408 16670 32464
rect 16726 32408 17406 32464
rect 17462 32408 17467 32464
rect 16665 32406 17467 32408
rect 16665 32403 16731 32406
rect 17401 32403 17467 32406
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31908 800 31998
rect 2773 31995 2839 31998
rect 47301 32058 47367 32061
rect 49200 32058 50000 32148
rect 47301 32056 50000 32058
rect 47301 32000 47306 32056
rect 47362 32000 50000 32056
rect 47301 31998 50000 32000
rect 47301 31995 47367 31998
rect 49200 31908 50000 31998
rect 23013 31650 23079 31653
rect 27981 31650 28047 31653
rect 23013 31648 28047 31650
rect 23013 31592 23018 31648
rect 23074 31592 27986 31648
rect 28042 31592 28047 31648
rect 23013 31590 28047 31592
rect 23013 31587 23079 31590
rect 27981 31587 28047 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3785 31378 3851 31381
rect 0 31376 3851 31378
rect 0 31320 3790 31376
rect 3846 31320 3851 31376
rect 0 31318 3851 31320
rect 0 31228 800 31318
rect 3785 31315 3851 31318
rect 46381 31378 46447 31381
rect 49200 31378 50000 31468
rect 46381 31376 50000 31378
rect 46381 31320 46386 31376
rect 46442 31320 50000 31376
rect 46381 31318 50000 31320
rect 46381 31315 46447 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 25221 30018 25287 30021
rect 27337 30018 27403 30021
rect 25221 30016 27403 30018
rect 25221 29960 25226 30016
rect 25282 29960 27342 30016
rect 27398 29960 27403 30016
rect 25221 29958 27403 29960
rect 25221 29955 25287 29958
rect 27337 29955 27403 29958
rect 46565 30018 46631 30021
rect 49200 30018 50000 30108
rect 46565 30016 50000 30018
rect 46565 29960 46570 30016
rect 46626 29960 50000 30016
rect 46565 29958 50000 29960
rect 46565 29955 46631 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47301 29338 47367 29341
rect 49200 29338 50000 29428
rect 47301 29336 50000 29338
rect 47301 29280 47306 29336
rect 47362 29280 50000 29336
rect 47301 29278 50000 29280
rect 47301 29275 47367 29278
rect 49200 29188 50000 29278
rect 21541 29066 21607 29069
rect 24945 29066 25011 29069
rect 26049 29066 26115 29069
rect 21541 29064 26115 29066
rect 21541 29008 21546 29064
rect 21602 29008 24950 29064
rect 25006 29008 26054 29064
rect 26110 29008 26115 29064
rect 21541 29006 26115 29008
rect 21541 29003 21607 29006
rect 24945 29003 25011 29006
rect 26049 29003 26115 29006
rect 20345 28930 20411 28933
rect 28257 28930 28323 28933
rect 20345 28928 28323 28930
rect 20345 28872 20350 28928
rect 20406 28872 28262 28928
rect 28318 28872 28323 28928
rect 20345 28870 28323 28872
rect 20345 28867 20411 28870
rect 28257 28867 28323 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3969 28658 4035 28661
rect 0 28656 4035 28658
rect 0 28600 3974 28656
rect 4030 28600 4035 28656
rect 0 28598 4035 28600
rect 0 28508 800 28598
rect 3969 28595 4035 28598
rect 45737 28658 45803 28661
rect 49200 28658 50000 28748
rect 45737 28656 50000 28658
rect 45737 28600 45742 28656
rect 45798 28600 50000 28656
rect 45737 28598 50000 28600
rect 45737 28595 45803 28598
rect 49200 28508 50000 28598
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 30189 28114 30255 28117
rect 30925 28114 30991 28117
rect 30189 28112 30991 28114
rect 0 27828 800 28068
rect 30189 28056 30194 28112
rect 30250 28056 30930 28112
rect 30986 28056 30991 28112
rect 30189 28054 30991 28056
rect 30189 28051 30255 28054
rect 30925 28051 30991 28054
rect 46841 27978 46907 27981
rect 49200 27978 50000 28068
rect 46841 27976 50000 27978
rect 46841 27920 46846 27976
rect 46902 27920 50000 27976
rect 46841 27918 50000 27920
rect 46841 27915 46907 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 46565 26618 46631 26621
rect 49200 26618 50000 26708
rect 46565 26616 50000 26618
rect 46565 26560 46570 26616
rect 46626 26560 50000 26616
rect 46565 26558 50000 26560
rect 46565 26555 46631 26558
rect 49200 26468 50000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 46841 25938 46907 25941
rect 49200 25938 50000 26028
rect 46841 25936 50000 25938
rect 46841 25880 46846 25936
rect 46902 25880 50000 25936
rect 46841 25878 50000 25880
rect 46841 25875 46907 25878
rect 49200 25788 50000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 48129 25258 48195 25261
rect 49200 25258 50000 25348
rect 48129 25256 50000 25258
rect 48129 25200 48134 25256
rect 48190 25200 50000 25256
rect 48129 25198 50000 25200
rect 48129 25195 48195 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 24025 24986 24091 24989
rect 25221 24986 25287 24989
rect 24025 24984 25287 24986
rect 24025 24928 24030 24984
rect 24086 24928 25226 24984
rect 25282 24928 25287 24984
rect 24025 24926 25287 24928
rect 24025 24923 24091 24926
rect 25221 24923 25287 24926
rect 24853 24850 24919 24853
rect 26233 24850 26299 24853
rect 24853 24848 26299 24850
rect 24853 24792 24858 24848
rect 24914 24792 26238 24848
rect 26294 24792 26299 24848
rect 24853 24790 26299 24792
rect 24853 24787 24919 24790
rect 26233 24787 26299 24790
rect 24301 24714 24367 24717
rect 25221 24714 25287 24717
rect 24301 24712 25287 24714
rect 0 24428 800 24668
rect 24301 24656 24306 24712
rect 24362 24656 25226 24712
rect 25282 24656 25287 24712
rect 24301 24654 25287 24656
rect 24301 24651 24367 24654
rect 25221 24651 25287 24654
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46749 23898 46815 23901
rect 49200 23898 50000 23988
rect 46749 23896 50000 23898
rect 46749 23840 46754 23896
rect 46810 23840 50000 23896
rect 46749 23838 50000 23840
rect 46749 23835 46815 23838
rect 49200 23748 50000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 46197 23218 46263 23221
rect 49200 23218 50000 23308
rect 46197 23216 50000 23218
rect 46197 23160 46202 23216
rect 46258 23160 50000 23216
rect 46197 23158 50000 23160
rect 46197 23155 46263 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46749 22538 46815 22541
rect 49200 22538 50000 22628
rect 46749 22536 50000 22538
rect 46749 22480 46754 22536
rect 46810 22480 50000 22536
rect 46749 22478 50000 22480
rect 46749 22475 46815 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 45369 21858 45435 21861
rect 49200 21858 50000 21948
rect 45369 21856 50000 21858
rect 45369 21800 45374 21856
rect 45430 21800 50000 21856
rect 45369 21798 50000 21800
rect 45369 21795 45435 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 20069 21042 20135 21045
rect 26601 21042 26667 21045
rect 20069 21040 26667 21042
rect 20069 20984 20074 21040
rect 20130 20984 26606 21040
rect 26662 20984 26667 21040
rect 49200 21028 50000 21118
rect 20069 20982 26667 20984
rect 20069 20979 20135 20982
rect 26601 20979 26667 20982
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 1945 20498 2011 20501
rect 27797 20498 27863 20501
rect 1945 20496 27863 20498
rect 1945 20440 1950 20496
rect 2006 20440 27802 20496
rect 27858 20440 27863 20496
rect 1945 20438 27863 20440
rect 1945 20435 2011 20438
rect 27797 20435 27863 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 3233 19954 3299 19957
rect 27797 19954 27863 19957
rect 3233 19952 27863 19954
rect 0 19818 800 19908
rect 3233 19896 3238 19952
rect 3294 19896 27802 19952
rect 27858 19896 27863 19952
rect 3233 19894 27863 19896
rect 3233 19891 3299 19894
rect 27797 19891 27863 19894
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18308 800 18398
rect 3969 18395 4035 18398
rect 46841 18458 46907 18461
rect 49200 18458 50000 18548
rect 46841 18456 50000 18458
rect 46841 18400 46846 18456
rect 46902 18400 50000 18456
rect 46841 18398 50000 18400
rect 46841 18395 46907 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 1853 17778 1919 17781
rect 0 17776 1919 17778
rect 0 17720 1858 17776
rect 1914 17720 1919 17776
rect 0 17718 1919 17720
rect 0 17628 800 17718
rect 1853 17715 1919 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3969 17098 4035 17101
rect 0 17096 4035 17098
rect 0 17040 3974 17096
rect 4030 17040 4035 17096
rect 0 17038 4035 17040
rect 0 16948 800 17038
rect 3969 17035 4035 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16268 800 16358
rect 2773 16355 2839 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16508
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 45553 15738 45619 15741
rect 49200 15738 50000 15828
rect 45553 15736 50000 15738
rect 45553 15680 45558 15736
rect 45614 15680 50000 15736
rect 45553 15678 50000 15680
rect 45553 15675 45619 15678
rect 27153 15602 27219 15605
rect 46054 15602 46060 15604
rect 27153 15600 46060 15602
rect 27153 15544 27158 15600
rect 27214 15544 46060 15600
rect 27153 15542 46060 15544
rect 27153 15539 27219 15542
rect 46054 15540 46060 15542
rect 46124 15540 46130 15604
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 17677 13970 17743 13973
rect 18781 13970 18847 13973
rect 17677 13968 18847 13970
rect 17677 13912 17682 13968
rect 17738 13912 18786 13968
rect 18842 13912 18847 13968
rect 17677 13910 18847 13912
rect 17677 13907 17743 13910
rect 18781 13907 18847 13910
rect 0 13698 800 13788
rect 3785 13698 3851 13701
rect 0 13696 3851 13698
rect 0 13640 3790 13696
rect 3846 13640 3851 13696
rect 0 13638 3851 13640
rect 0 13548 800 13638
rect 3785 13635 3851 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10148 800 10238
rect 2773 10235 2839 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 46197 9618 46263 9621
rect 49200 9618 50000 9708
rect 46197 9616 50000 9618
rect 46197 9560 46202 9616
rect 46258 9560 50000 9616
rect 46197 9558 50000 9560
rect 46197 9555 46263 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3141 7578 3207 7581
rect 0 7576 3207 7578
rect 0 7520 3146 7576
rect 3202 7520 3207 7576
rect 0 7518 3207 7520
rect 0 7428 800 7518
rect 3141 7515 3207 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 46841 6218 46907 6221
rect 49200 6218 50000 6308
rect 46841 6216 50000 6218
rect 46841 6160 46846 6216
rect 46902 6160 50000 6216
rect 46841 6158 50000 6160
rect 46841 6155 46907 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 21725 4178 21791 4181
rect 26969 4178 27035 4181
rect 21725 4176 27035 4178
rect 21725 4120 21730 4176
rect 21786 4120 26974 4176
rect 27030 4120 27035 4176
rect 21725 4118 27035 4120
rect 21725 4115 21791 4118
rect 26969 4115 27035 4118
rect 48129 4178 48195 4181
rect 49200 4178 50000 4268
rect 48129 4176 50000 4178
rect 48129 4120 48134 4176
rect 48190 4120 50000 4176
rect 48129 4118 50000 4120
rect 48129 4115 48195 4118
rect 3969 4042 4035 4045
rect 29453 4042 29519 4045
rect 3969 4040 29519 4042
rect 3969 3984 3974 4040
rect 4030 3984 29458 4040
rect 29514 3984 29519 4040
rect 49200 4028 50000 4118
rect 3969 3982 29519 3984
rect 3969 3979 4035 3982
rect 29453 3979 29519 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 22093 3634 22159 3637
rect 24853 3634 24919 3637
rect 22093 3632 24919 3634
rect 0 3498 800 3588
rect 22093 3576 22098 3632
rect 22154 3576 24858 3632
rect 24914 3576 24919 3632
rect 22093 3574 24919 3576
rect 22093 3571 22159 3574
rect 24853 3571 24919 3574
rect 3601 3498 3667 3501
rect 0 3496 3667 3498
rect 0 3440 3606 3496
rect 3662 3440 3667 3496
rect 0 3438 3667 3440
rect 0 3348 800 3438
rect 3601 3435 3667 3438
rect 21909 3498 21975 3501
rect 22645 3498 22711 3501
rect 21909 3496 22711 3498
rect 21909 3440 21914 3496
rect 21970 3440 22650 3496
rect 22706 3440 22711 3496
rect 21909 3438 22711 3440
rect 21909 3435 21975 3438
rect 22645 3435 22711 3438
rect 23381 3498 23447 3501
rect 25313 3498 25379 3501
rect 23381 3496 25379 3498
rect 23381 3440 23386 3496
rect 23442 3440 25318 3496
rect 25374 3440 25379 3496
rect 23381 3438 25379 3440
rect 23381 3435 23447 3438
rect 25313 3435 25379 3438
rect 39021 3498 39087 3501
rect 40493 3498 40559 3501
rect 39021 3496 40559 3498
rect 39021 3440 39026 3496
rect 39082 3440 40498 3496
rect 40554 3440 40559 3496
rect 39021 3438 40559 3440
rect 39021 3435 39087 3438
rect 40493 3435 40559 3438
rect 46657 3498 46723 3501
rect 49200 3498 50000 3588
rect 46657 3496 50000 3498
rect 46657 3440 46662 3496
rect 46718 3440 50000 3496
rect 46657 3438 50000 3440
rect 46657 3435 46723 3438
rect 21449 3362 21515 3365
rect 27613 3362 27679 3365
rect 21449 3360 27679 3362
rect 21449 3304 21454 3360
rect 21510 3304 27618 3360
rect 27674 3304 27679 3360
rect 49200 3348 50000 3438
rect 21449 3302 27679 3304
rect 21449 3299 21515 3302
rect 27613 3299 27679 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 19241 3090 19307 3093
rect 22277 3090 22343 3093
rect 19241 3088 22343 3090
rect 19241 3032 19246 3088
rect 19302 3032 22282 3088
rect 22338 3032 22343 3088
rect 19241 3030 22343 3032
rect 19241 3027 19307 3030
rect 22277 3027 22343 3030
rect 19885 2954 19951 2957
rect 24853 2954 24919 2957
rect 19885 2952 24919 2954
rect 0 2668 800 2908
rect 19885 2896 19890 2952
rect 19946 2896 24858 2952
rect 24914 2896 24919 2952
rect 19885 2894 24919 2896
rect 19885 2891 19951 2894
rect 24853 2891 24919 2894
rect 17677 2818 17743 2821
rect 21357 2818 21423 2821
rect 17677 2816 21423 2818
rect 17677 2760 17682 2816
rect 17738 2760 21362 2816
rect 21418 2760 21423 2816
rect 17677 2758 21423 2760
rect 17677 2755 17743 2758
rect 21357 2755 21423 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1308 800 1398
rect 3325 1395 3391 1398
rect 47761 1458 47827 1461
rect 49200 1458 50000 1548
rect 47761 1456 50000 1458
rect 47761 1400 47766 1456
rect 47822 1400 50000 1456
rect 47761 1398 50000 1400
rect 47761 1395 47827 1398
rect 49200 1308 50000 1398
rect 46841 914 46907 917
rect 46841 912 47042 914
rect 0 778 800 868
rect 46841 856 46846 912
rect 46902 856 47042 912
rect 46841 854 47042 856
rect 46841 851 46907 854
rect 2957 778 3023 781
rect 0 776 3023 778
rect 0 720 2962 776
rect 3018 720 3023 776
rect 0 718 3023 720
rect 46982 778 47042 854
rect 49200 778 50000 868
rect 46982 718 50000 778
rect 0 628 800 718
rect 2957 715 3023 718
rect 49200 628 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 188
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 46060 46956 46124 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 46060 15540 46124 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 46059 47020 46125 47021
rect 46059 46956 46060 47020
rect 46124 46956 46125 47020
rect 46059 46955 46125 46956
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 46062 15605 46122 46955
rect 46059 15604 46125 15605
rect 46059 15540 46060 15604
rect 46124 15540 46125 15604
rect 46059 15539 46125 15540
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 29164 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 27784 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 30544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 26220 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_242
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1644511149
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1644511149
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_64
timestamp 1644511149
transform 1 0 6992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_68
timestamp 1644511149
transform 1 0 7360 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_95
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_177
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1644511149
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_203
timestamp 1644511149
transform 1 0 19780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1644511149
transform 1 0 20792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1644511149
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_345
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_368
timestamp 1644511149
transform 1 0 34960 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_380
timestamp 1644511149
transform 1 0 36064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1644511149
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_88
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1644511149
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1644511149
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_125
timestamp 1644511149
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1644511149
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1644511149
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_262
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_282
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_350
timestamp 1644511149
transform 1 0 33304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1644511149
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_399
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_411
timestamp 1644511149
transform 1 0 38916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_442
timestamp 1644511149
transform 1 0 41768 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_450
timestamp 1644511149
transform 1 0 42504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_116
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp 1644511149
transform 1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1644511149
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_209
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1644511149
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1644511149
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_262
timestamp 1644511149
transform 1 0 25208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1644511149
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_345
timestamp 1644511149
transform 1 0 32844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_351
timestamp 1644511149
transform 1 0 33396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_363
timestamp 1644511149
transform 1 0 34500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_375
timestamp 1644511149
transform 1 0 35604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_413
timestamp 1644511149
transform 1 0 39100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_418
timestamp 1644511149
transform 1 0 39560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_425
timestamp 1644511149
transform 1 0 40204 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_433
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_442
timestamp 1644511149
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_490
timestamp 1644511149
transform 1 0 46184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1644511149
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_104
timestamp 1644511149
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_116
timestamp 1644511149
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1644511149
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_200
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_211
timestamp 1644511149
transform 1 0 20516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1644511149
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1644511149
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_424
timestamp 1644511149
transform 1 0 40112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_436
timestamp 1644511149
transform 1 0 41216 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_448
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_455
timestamp 1644511149
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_467
timestamp 1644511149
transform 1 0 44068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_482
timestamp 1644511149
transform 1 0 45448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_507
timestamp 1644511149
transform 1 0 47748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_515
timestamp 1644511149
transform 1 0 48484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1644511149
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_203
timestamp 1644511149
transform 1 0 19780 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1644511149
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_247
timestamp 1644511149
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_259
timestamp 1644511149
transform 1 0 24932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1644511149
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_494
timestamp 1644511149
transform 1 0 46552 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1644511149
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1644511149
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_217
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1644511149
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1644511149
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1644511149
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1644511149
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_486
timestamp 1644511149
transform 1 0 45816 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1644511149
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_146
timestamp 1644511149
transform 1 0 14536 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_158
timestamp 1644511149
transform 1 0 15640 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1644511149
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_194
timestamp 1644511149
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1644511149
transform 1 0 19596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1644511149
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1644511149
transform 1 0 15640 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1644511149
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_200
timestamp 1644511149
transform 1 0 19504 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_236
timestamp 1644511149
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1644511149
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_489
timestamp 1644511149
transform 1 0 46092 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1644511149
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1644511149
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_492
timestamp 1644511149
transform 1 0 46368 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1644511149
transform 1 0 47012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1644511149
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_212
timestamp 1644511149
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_224
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1644511149
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_156
timestamp 1644511149
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_182
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_206
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1644511149
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1644511149
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1644511149
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_175
timestamp 1644511149
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_206
timestamp 1644511149
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_210
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_234
timestamp 1644511149
transform 1 0 22632 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1644511149
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1644511149
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1644511149
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1644511149
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1644511149
transform 1 0 17020 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_188
timestamp 1644511149
transform 1 0 18400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_228
timestamp 1644511149
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_240
timestamp 1644511149
transform 1 0 23184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_252
timestamp 1644511149
transform 1 0 24288 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_264
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1644511149
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1644511149
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 1644511149
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_208
timestamp 1644511149
transform 1 0 20240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1644511149
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1644511149
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_157
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1644511149
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_186
timestamp 1644511149
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_233
timestamp 1644511149
transform 1 0 22540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1644511149
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1644511149
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_173
timestamp 1644511149
transform 1 0 17020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_218
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1644511149
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1644511149
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_153
timestamp 1644511149
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1644511149
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_197
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_209
timestamp 1644511149
transform 1 0 20332 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_267
timestamp 1644511149
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1644511149
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1644511149
transform 1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1644511149
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_163
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1644511149
transform 1 0 17204 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1644511149
transform 1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_210
timestamp 1644511149
transform 1 0 20424 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1644511149
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_240
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_284
timestamp 1644511149
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_296
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_133
timestamp 1644511149
transform 1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1644511149
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_252
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_493
timestamp 1644511149
transform 1 0 46460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1644511149
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1644511149
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_73
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1644511149
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1644511149
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1644511149
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1644511149
transform 1 0 12880 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1644511149
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1644511149
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1644511149
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1644511149
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1644511149
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_101
timestamp 1644511149
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_173
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1644511149
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1644511149
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_302
timestamp 1644511149
transform 1 0 28888 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_314
timestamp 1644511149
transform 1 0 29992 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_326
timestamp 1644511149
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_472
timestamp 1644511149
transform 1 0 44528 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_484
timestamp 1644511149
transform 1 0 45632 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_496
timestamp 1644511149
transform 1 0 46736 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_14
timestamp 1644511149
transform 1 0 2392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1644511149
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_92
timestamp 1644511149
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_117
timestamp 1644511149
transform 1 0 11868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1644511149
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1644511149
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_201
timestamp 1644511149
transform 1 0 19596 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1644511149
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_241
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1644511149
transform 1 0 27600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_465
timestamp 1644511149
transform 1 0 43884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_482
timestamp 1644511149
transform 1 0 45448 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_490
timestamp 1644511149
transform 1 0 46184 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1644511149
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1644511149
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1644511149
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_102
timestamp 1644511149
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1644511149
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_119
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_145
timestamp 1644511149
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_194
timestamp 1644511149
transform 1 0 18952 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_202
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1644511149
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1644511149
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_289
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1644511149
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1644511149
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_465
timestamp 1644511149
transform 1 0 43884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_483
timestamp 1644511149
transform 1 0 45540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_492
timestamp 1644511149
transform 1 0 46368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_496
timestamp 1644511149
transform 1 0 46736 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_105
timestamp 1644511149
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1644511149
transform 1 0 12972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1644511149
transform 1 0 14536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1644511149
transform 1 0 15272 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_161
timestamp 1644511149
transform 1 0 15916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_231
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_266
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_285
timestamp 1644511149
transform 1 0 27324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_336
timestamp 1644511149
transform 1 0 32016 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_348
timestamp 1644511149
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_463
timestamp 1644511149
transform 1 0 43700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_467
timestamp 1644511149
transform 1 0 44068 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1644511149
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_482
timestamp 1644511149
transform 1 0 45448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_490
timestamp 1644511149
transform 1 0 46184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1644511149
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1644511149
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_230
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_257
timestamp 1644511149
transform 1 0 24748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1644511149
transform 1 0 28152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1644511149
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_433
timestamp 1644511149
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1644511149
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_468
timestamp 1644511149
transform 1 0 44160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1644511149
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1644511149
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1644511149
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_180
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_217
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1644511149
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_256
timestamp 1644511149
transform 1 0 24656 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_278
timestamp 1644511149
transform 1 0 26680 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_284
timestamp 1644511149
transform 1 0 27232 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_290
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_338
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_350
timestamp 1644511149
transform 1 0 33304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1644511149
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_450
timestamp 1644511149
transform 1 0 42504 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_458
timestamp 1644511149
transform 1 0 43240 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_484
timestamp 1644511149
transform 1 0 45632 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_490
timestamp 1644511149
transform 1 0 46184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1644511149
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_96
timestamp 1644511149
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_210
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1644511149
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_230
timestamp 1644511149
transform 1 0 22264 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_434
timestamp 1644511149
transform 1 0 41032 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1644511149
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_475
timestamp 1644511149
transform 1 0 44804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1644511149
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_95
timestamp 1644511149
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_119
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1644511149
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_173
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1644511149
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_208
timestamp 1644511149
transform 1 0 20240 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1644511149
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_267
timestamp 1644511149
transform 1 0 25668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_271
timestamp 1644511149
transform 1 0 26036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_293
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1644511149
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_330
timestamp 1644511149
transform 1 0 31464 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_342
timestamp 1644511149
transform 1 0 32568 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_461
timestamp 1644511149
transform 1 0 43516 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_465
timestamp 1644511149
transform 1 0 43884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_472
timestamp 1644511149
transform 1 0 44528 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_485
timestamp 1644511149
transform 1 0 45724 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_73
timestamp 1644511149
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_95
timestamp 1644511149
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_116
timestamp 1644511149
transform 1 0 11776 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_123
timestamp 1644511149
transform 1 0 12420 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1644511149
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1644511149
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_228
timestamp 1644511149
transform 1 0 22080 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_236
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_456
timestamp 1644511149
transform 1 0 43056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_482
timestamp 1644511149
transform 1 0 45448 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_499
timestamp 1644511149
transform 1 0 47012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_508
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1644511149
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_182
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1644511149
transform 1 0 21804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_237
timestamp 1644511149
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1644511149
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_290
timestamp 1644511149
transform 1 0 27784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_463
timestamp 1644511149
transform 1 0 43700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1644511149
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_487
timestamp 1644511149
transform 1 0 45908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_89
timestamp 1644511149
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_96
timestamp 1644511149
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_121
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_130
timestamp 1644511149
transform 1 0 13064 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_138
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_142
timestamp 1644511149
transform 1 0 14168 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_150
timestamp 1644511149
transform 1 0 14904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_154
timestamp 1644511149
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1644511149
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1644511149
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_228
timestamp 1644511149
transform 1 0 22080 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_302
timestamp 1644511149
transform 1 0 28888 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_314
timestamp 1644511149
transform 1 0 29992 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_326
timestamp 1644511149
transform 1 0 31096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1644511149
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_470
timestamp 1644511149
transform 1 0 44344 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_478
timestamp 1644511149
transform 1 0 45080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_123
timestamp 1644511149
transform 1 0 12420 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_145
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_157
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_161
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_169
timestamp 1644511149
transform 1 0 16652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_178
timestamp 1644511149
transform 1 0 17480 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_204
timestamp 1644511149
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_268
timestamp 1644511149
transform 1 0 25760 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_278
timestamp 1644511149
transform 1 0 26680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_285
timestamp 1644511149
transform 1 0 27324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_294
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_315
timestamp 1644511149
transform 1 0 30084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_322
timestamp 1644511149
transform 1 0 30728 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_334
timestamp 1644511149
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_346
timestamp 1644511149
transform 1 0 32936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1644511149
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1644511149
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_92
timestamp 1644511149
transform 1 0 9568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_120
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_128
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_152
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_156
timestamp 1644511149
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_175
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_184
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_190
timestamp 1644511149
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_196
timestamp 1644511149
transform 1 0 19136 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_209
timestamp 1644511149
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1644511149
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1644511149
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1644511149
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_314
timestamp 1644511149
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_325
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_489
timestamp 1644511149
transform 1 0 46092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_73
timestamp 1644511149
transform 1 0 7820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1644511149
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1644511149
transform 1 0 10764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_116
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_178
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1644511149
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_273
timestamp 1644511149
transform 1 0 26220 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_322
timestamp 1644511149
transform 1 0 30728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_346
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1644511149
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1644511149
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_128
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_136
timestamp 1644511149
transform 1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1644511149
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1644511149
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_214
timestamp 1644511149
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1644511149
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_238
timestamp 1644511149
transform 1 0 23000 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1644511149
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_267
timestamp 1644511149
transform 1 0 25668 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_299
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_307
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_316
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_320
timestamp 1644511149
transform 1 0 30544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_341
timestamp 1644511149
transform 1 0 32476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_353
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_365
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_92
timestamp 1644511149
transform 1 0 9568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1644511149
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1644511149
transform 1 0 11592 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1644511149
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_158
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_179
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1644511149
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_212
timestamp 1644511149
transform 1 0 20608 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_220
timestamp 1644511149
transform 1 0 21344 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_229
timestamp 1644511149
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1644511149
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_283
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1644511149
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_314
timestamp 1644511149
transform 1 0 29992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_335
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_347
timestamp 1644511149
transform 1 0 33028 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1644511149
transform 1 0 33396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_85
timestamp 1644511149
transform 1 0 8924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_130
timestamp 1644511149
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_151
timestamp 1644511149
transform 1 0 14996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_190
timestamp 1644511149
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_214
timestamp 1644511149
transform 1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_245
timestamp 1644511149
transform 1 0 23644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_265
timestamp 1644511149
transform 1 0 25484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_284
timestamp 1644511149
transform 1 0 27232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_296
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_330
timestamp 1644511149
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_358
timestamp 1644511149
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_370
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1644511149
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_106
timestamp 1644511149
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_117
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_125
timestamp 1644511149
transform 1 0 12604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1644511149
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_171
timestamp 1644511149
transform 1 0 16836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_183
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_206
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_214
timestamp 1644511149
transform 1 0 20792 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1644511149
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_232
timestamp 1644511149
transform 1 0 22448 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1644511149
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_260
timestamp 1644511149
transform 1 0 25024 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_267
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_279
timestamp 1644511149
transform 1 0 26772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_300
timestamp 1644511149
transform 1 0 28704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_312
timestamp 1644511149
transform 1 0 29808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_320
timestamp 1644511149
transform 1 0 30544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_328
timestamp 1644511149
transform 1 0 31280 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_332
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_342
timestamp 1644511149
transform 1 0 32568 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_354
timestamp 1644511149
transform 1 0 33672 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1644511149
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_80
timestamp 1644511149
transform 1 0 8464 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_88
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_100
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1644511149
transform 1 0 14536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1644511149
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_188
timestamp 1644511149
transform 1 0 18400 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_210
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_244
timestamp 1644511149
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_256
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_268
timestamp 1644511149
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_284
timestamp 1644511149
transform 1 0 27232 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_290
timestamp 1644511149
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_311
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_323
timestamp 1644511149
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_346
timestamp 1644511149
transform 1 0 32936 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_358
timestamp 1644511149
transform 1 0 34040 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_370
timestamp 1644511149
transform 1 0 35144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_382
timestamp 1644511149
transform 1 0 36248 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1644511149
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_118
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_130
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1644511149
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_218
timestamp 1644511149
transform 1 0 21160 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_227
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_235
timestamp 1644511149
transform 1 0 22724 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_241
timestamp 1644511149
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1644511149
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_257
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_263
timestamp 1644511149
transform 1 0 25300 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_284
timestamp 1644511149
transform 1 0 27232 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1644511149
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_313
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_319
timestamp 1644511149
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_331
timestamp 1644511149
transform 1 0 31556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_337
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_358
timestamp 1644511149
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_394
timestamp 1644511149
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_406
timestamp 1644511149
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1644511149
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_77
timestamp 1644511149
transform 1 0 8188 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_100
timestamp 1644511149
transform 1 0 10304 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_133
timestamp 1644511149
transform 1 0 13340 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_139
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_147
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_154
timestamp 1644511149
transform 1 0 15272 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1644511149
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_207
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1644511149
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1644511149
transform 1 0 23644 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_255
timestamp 1644511149
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_268
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1644511149
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_312
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_323
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_343
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_347
timestamp 1644511149
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_359
timestamp 1644511149
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_371
timestamp 1644511149
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1644511149
transform 1 0 36616 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_414
timestamp 1644511149
transform 1 0 39192 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_426
timestamp 1644511149
transform 1 0 40296 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_438
timestamp 1644511149
transform 1 0 41400 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1644511149
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1644511149
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_174
timestamp 1644511149
transform 1 0 17112 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_186
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1644511149
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_232
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1644511149
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_264
timestamp 1644511149
transform 1 0 25392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_288
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_293
timestamp 1644511149
transform 1 0 28060 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_297
timestamp 1644511149
transform 1 0 28428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_314
timestamp 1644511149
transform 1 0 29992 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_320
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_327
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_335
timestamp 1644511149
transform 1 0 31924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_349
timestamp 1644511149
transform 1 0 33212 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_353
timestamp 1644511149
transform 1 0 33580 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1644511149
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_157
timestamp 1644511149
transform 1 0 15548 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_212
timestamp 1644511149
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_234
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_243
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_260
timestamp 1644511149
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_309
timestamp 1644511149
transform 1 0 29532 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_315
timestamp 1644511149
transform 1 0 30084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_323
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1644511149
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_341
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_362
timestamp 1644511149
transform 1 0 34408 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_374
timestamp 1644511149
transform 1 0 35512 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1644511149
transform 1 0 36616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_149
timestamp 1644511149
transform 1 0 14812 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_171
timestamp 1644511149
transform 1 0 16836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_184
timestamp 1644511149
transform 1 0 18032 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_203
timestamp 1644511149
transform 1 0 19780 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1644511149
transform 1 0 20884 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1644511149
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1644511149
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_257
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_298
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1644511149
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_313
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_322
timestamp 1644511149
transform 1 0 30728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_332
timestamp 1644511149
transform 1 0 31648 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_340
timestamp 1644511149
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_352
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 1644511149
transform 1 0 17480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_198
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_204
timestamp 1644511149
transform 1 0 19872 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1644511149
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1644511149
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_263
timestamp 1644511149
transform 1 0 25300 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_288
timestamp 1644511149
transform 1 0 27600 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_292
timestamp 1644511149
transform 1 0 27968 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_299
timestamp 1644511149
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_318
timestamp 1644511149
transform 1 0 30360 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_326
timestamp 1644511149
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1644511149
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_341
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_353
timestamp 1644511149
transform 1 0 33580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_365
timestamp 1644511149
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_377
timestamp 1644511149
transform 1 0 35788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1644511149
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_161
timestamp 1644511149
transform 1 0 15916 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_166
timestamp 1644511149
transform 1 0 16376 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_174
timestamp 1644511149
transform 1 0 17112 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1644511149
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_202
timestamp 1644511149
transform 1 0 19688 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_214
timestamp 1644511149
transform 1 0 20792 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_222
timestamp 1644511149
transform 1 0 21528 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_238
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_288
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_313
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_188
timestamp 1644511149
transform 1 0 18400 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_200
timestamp 1644511149
transform 1 0 19504 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_208
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_241
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_255
timestamp 1644511149
transform 1 0 24564 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_272
timestamp 1644511149
transform 1 0 26128 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_319
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_327
timestamp 1644511149
transform 1 0 31188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_10
timestamp 1644511149
transform 1 0 2024 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_14
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_149
timestamp 1644511149
transform 1 0 14812 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_174
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_204
timestamp 1644511149
transform 1 0 19872 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1644511149
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_224
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_229
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_237
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1644511149
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_263
timestamp 1644511149
transform 1 0 25300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_275
timestamp 1644511149
transform 1 0 26404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_281
timestamp 1644511149
transform 1 0 26956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_326
timestamp 1644511149
transform 1 0 31096 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_338
timestamp 1644511149
transform 1 0 32200 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_350
timestamp 1644511149
transform 1 0 33304 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 1644511149
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_29
timestamp 1644511149
transform 1 0 3772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_41
timestamp 1644511149
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1644511149
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_153
timestamp 1644511149
transform 1 0 15180 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1644511149
transform 1 0 17296 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_180
timestamp 1644511149
transform 1 0 17664 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_189
timestamp 1644511149
transform 1 0 18492 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_198
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_206
timestamp 1644511149
transform 1 0 20056 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_253
timestamp 1644511149
transform 1 0 24380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_263
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp 1644511149
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_289
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1644511149
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_314
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_173
timestamp 1644511149
transform 1 0 17020 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 1644511149
transform 1 0 17940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_207
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_211
timestamp 1644511149
transform 1 0 20516 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_216
timestamp 1644511149
transform 1 0 20976 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_220
timestamp 1644511149
transform 1 0 21344 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_232
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_238
timestamp 1644511149
transform 1 0 23000 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_262
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_272
timestamp 1644511149
transform 1 0 26128 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_279
timestamp 1644511149
transform 1 0 26772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_295
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_322
timestamp 1644511149
transform 1 0 30728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_326
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_347
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1644511149
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_177
timestamp 1644511149
transform 1 0 17388 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_185
timestamp 1644511149
transform 1 0 18124 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_201
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_212
timestamp 1644511149
transform 1 0 20608 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_232
timestamp 1644511149
transform 1 0 22448 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_242
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_264
timestamp 1644511149
transform 1 0 25392 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1644511149
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_294
timestamp 1644511149
transform 1 0 28152 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_307
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_326
timestamp 1644511149
transform 1 0 31096 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1644511149
transform 1 0 16560 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1644511149
transform 1 0 17664 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_205
timestamp 1644511149
transform 1 0 19964 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1644511149
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_263
timestamp 1644511149
transform 1 0 25300 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_272
timestamp 1644511149
transform 1 0 26128 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_284
timestamp 1644511149
transform 1 0 27232 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_291
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_318
timestamp 1644511149
transform 1 0 30360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_328
timestamp 1644511149
transform 1 0 31280 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_332
timestamp 1644511149
transform 1 0 31648 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_336
timestamp 1644511149
transform 1 0 32016 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_348
timestamp 1644511149
transform 1 0 33120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_157
timestamp 1644511149
transform 1 0 15548 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_176
timestamp 1644511149
transform 1 0 17296 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_180
timestamp 1644511149
transform 1 0 17664 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_190
timestamp 1644511149
transform 1 0 18584 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_213
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1644511149
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_234
timestamp 1644511149
transform 1 0 22632 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_246
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_250
timestamp 1644511149
transform 1 0 24104 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_284
timestamp 1644511149
transform 1 0 27232 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_292
timestamp 1644511149
transform 1 0 27968 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_304
timestamp 1644511149
transform 1 0 29072 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_10
timestamp 1644511149
transform 1 0 2024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_14
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1644511149
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_168
timestamp 1644511149
transform 1 0 16560 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_218
timestamp 1644511149
transform 1 0 21160 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_271
timestamp 1644511149
transform 1 0 26036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_292
timestamp 1644511149
transform 1 0 27968 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_312
timestamp 1644511149
transform 1 0 29808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_324
timestamp 1644511149
transform 1 0 30912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_329
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_341
timestamp 1644511149
transform 1 0 32476 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_353
timestamp 1644511149
transform 1 0 33580 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_361
timestamp 1644511149
transform 1 0 34316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1644511149
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1644511149
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1644511149
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1644511149
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_235
timestamp 1644511149
transform 1 0 22724 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_243
timestamp 1644511149
transform 1 0 23460 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_250
timestamp 1644511149
transform 1 0 24104 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_262
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1644511149
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_286
timestamp 1644511149
transform 1 0 27416 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_294
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_315
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1644511149
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_201
timestamp 1644511149
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_211
timestamp 1644511149
transform 1 0 20516 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_223
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1644511149
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1644511149
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_256
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_292
timestamp 1644511149
transform 1 0 27968 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_200
timestamp 1644511149
transform 1 0 19504 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_213
timestamp 1644511149
transform 1 0 20700 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_254
timestamp 1644511149
transform 1 0 24472 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_268
timestamp 1644511149
transform 1 0 25760 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_217
timestamp 1644511149
transform 1 0 21068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_229
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_243
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_263
timestamp 1644511149
transform 1 0 25300 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_271
timestamp 1644511149
transform 1 0 26036 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_275
timestamp 1644511149
transform 1 0 26404 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_286
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_298
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1644511149
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_507
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_202
timestamp 1644511149
transform 1 0 19688 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_214
timestamp 1644511149
transform 1 0 20792 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1644511149
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1644511149
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1644511149
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_14
timestamp 1644511149
transform 1 0 2392 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_499
timestamp 1644511149
transform 1 0 47012 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_512
timestamp 1644511149
transform 1 0 48208 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_264
timestamp 1644511149
transform 1 0 25392 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_37
timestamp 1644511149
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1644511149
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_272
timestamp 1644511149
transform 1 0 26128 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_479
timestamp 1644511149
transform 1 0 45172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_451
timestamp 1644511149
transform 1 0 42596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_455
timestamp 1644511149
transform 1 0 42964 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_467
timestamp 1644511149
transform 1 0 44068 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_9
timestamp 1644511149
transform 1 0 1932 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_31
timestamp 1644511149
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_43
timestamp 1644511149
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_140
timestamp 1644511149
transform 1 0 13984 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_152
timestamp 1644511149
transform 1 0 15088 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_340
timestamp 1644511149
transform 1 0 32384 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_376
timestamp 1644511149
transform 1 0 35696 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_437
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_456
timestamp 1644511149
transform 1 0 43056 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_468
timestamp 1644511149
transform 1 0 44160 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1644511149
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_22
timestamp 1644511149
transform 1 0 3128 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_39
timestamp 1644511149
transform 1 0 4692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_51
timestamp 1644511149
transform 1 0 5796 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_63
timestamp 1644511149
transform 1 0 6900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_75
timestamp 1644511149
transform 1 0 8004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_112
timestamp 1644511149
transform 1 0 11408 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_124
timestamp 1644511149
transform 1 0 12512 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_205
timestamp 1644511149
transform 1 0 19964 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_458
timestamp 1644511149
transform 1 0 43240 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1644511149
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_24
timestamp 1644511149
transform 1 0 3312 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1644511149
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1644511149
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_316
timestamp 1644511149
transform 1 0 30176 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_328
timestamp 1644511149
transform 1 0 31280 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_9
timestamp 1644511149
transform 1 0 1932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_16
timestamp 1644511149
transform 1 0 2576 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1644511149
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1644511149
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_191
timestamp 1644511149
transform 1 0 18676 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_228
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_240
timestamp 1644511149
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1644511149
transform 1 0 24840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_262
timestamp 1644511149
transform 1 0 25208 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_266
timestamp 1644511149
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_406
timestamp 1644511149
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_418
timestamp 1644511149
transform 1 0 39560 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_444
timestamp 1644511149
transform 1 0 41952 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0572_
timestamp 1644511149
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0574_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0577_
timestamp 1644511149
transform 1 0 21988 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0579_
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0580_
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0582_
timestamp 1644511149
transform 1 0 25668 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0583_
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0589_
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0590_
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0591_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0593_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0594_
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0600_
timestamp 1644511149
transform 1 0 27232 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0601_
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0602_
timestamp 1644511149
transform 1 0 23184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0604_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0605_
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_2  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0607_
timestamp 1644511149
transform 1 0 27876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0608_
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0611_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0612_
timestamp 1644511149
transform 1 0 17664 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0615_
timestamp 1644511149
transform 1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0616_
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0617_
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0620_
timestamp 1644511149
transform 1 0 16468 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0621_
timestamp 1644511149
transform 1 0 32016 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0622_
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0623_
timestamp 1644511149
transform 1 0 20148 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18952 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0625_
timestamp 1644511149
transform 1 0 18952 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1644511149
transform 1 0 19872 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1644511149
transform 1 0 19688 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0630_
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0632_
timestamp 1644511149
transform 1 0 30912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0633_
timestamp 1644511149
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0635_
timestamp 1644511149
transform 1 0 28704 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0636_
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0638_
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0639_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0640_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0641_
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1644511149
transform 1 0 25760 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0646_
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0647_
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0648_
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0649_
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0650_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0651_
timestamp 1644511149
transform 1 0 22724 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0652_
timestamp 1644511149
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0653_
timestamp 1644511149
transform 1 0 26496 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0656_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0657_
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0662_
timestamp 1644511149
transform 1 0 28612 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0663_
timestamp 1644511149
transform 1 0 30636 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0664_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28704 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0665_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0666_
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0667_
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0668_
timestamp 1644511149
transform 1 0 28244 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0669_
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 1644511149
transform 1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0671_
timestamp 1644511149
transform 1 0 30912 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0672_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0673_
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0674_
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0675_
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0676_
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0677_
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0678_
timestamp 1644511149
transform 1 0 23000 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0679_
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0681_
timestamp 1644511149
transform -1 0 29808 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0682_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1644511149
transform 1 0 25392 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0684_
timestamp 1644511149
transform 1 0 26036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1644511149
transform 1 0 24656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0686_
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0687_
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0689_
timestamp 1644511149
transform 1 0 24564 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0690_
timestamp 1644511149
transform 1 0 25852 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0691_
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1644511149
transform 1 0 22080 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0693_
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0694_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0695_
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform 1 0 26128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0702_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0704_
timestamp 1644511149
transform 1 0 21712 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0705_
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0706_
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0707_
timestamp 1644511149
transform 1 0 21252 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0708_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0710_
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0711_
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0712_
timestamp 1644511149
transform 1 0 31188 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0713_
timestamp 1644511149
transform 1 0 29992 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0715_
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0716_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0718_
timestamp 1644511149
transform 1 0 28428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0720_
timestamp 1644511149
transform 1 0 31096 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0721_
timestamp 1644511149
transform 1 0 30912 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0722_
timestamp 1644511149
transform 1 0 32016 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0723_
timestamp 1644511149
transform 1 0 30452 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1644511149
transform 1 0 29992 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0725_
timestamp 1644511149
transform 1 0 30636 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0727_
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0728_
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0729_
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1644511149
transform 1 0 30084 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0731_
timestamp 1644511149
transform 1 0 29532 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0732_
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1644511149
transform 1 0 30452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0735_
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0736_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0738_
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0739_
timestamp 1644511149
transform 1 0 14260 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0740_
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0743_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0745_
timestamp 1644511149
transform 1 0 12972 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0746_
timestamp 1644511149
transform 1 0 12696 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp 1644511149
transform 1 0 16744 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0748_
timestamp 1644511149
transform 1 0 16744 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0750_
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0751_
timestamp 1644511149
transform 1 0 13432 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0752_
timestamp 1644511149
transform 1 0 13892 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0754_
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0755_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0756_
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1644511149
transform 1 0 19044 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0758_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0759_
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0761_
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0762_
timestamp 1644511149
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0764_
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0766_
timestamp 1644511149
transform 1 0 18676 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0767_
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0768_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0769_
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0771_
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1644511149
transform 1 0 18124 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0775_
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0777_
timestamp 1644511149
transform 1 0 18308 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0778_
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1644511149
transform 1 0 16560 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0780_
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0781_
timestamp 1644511149
transform 1 0 13248 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0782_
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0785_
timestamp 1644511149
transform 1 0 12696 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _0786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0788_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0790_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1644511149
transform 1 0 11224 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0793_
timestamp 1644511149
transform 1 0 10580 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0794_
timestamp 1644511149
transform 1 0 8280 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0796_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0797_
timestamp 1644511149
transform 1 0 9016 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1644511149
transform 1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1644511149
transform 1 0 13892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0803_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0804_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0806_
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0809_
timestamp 1644511149
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0810_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0811_
timestamp 1644511149
transform 1 0 12144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0813_
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0814_
timestamp 1644511149
transform 1 0 11684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0816_
timestamp 1644511149
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1644511149
transform 1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0819_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0820_
timestamp 1644511149
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1644511149
transform 1 0 13064 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0823_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0826_
timestamp 1644511149
transform 1 0 13156 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1644511149
transform 1 0 15824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 1644511149
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform 1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0832_
timestamp 1644511149
transform 1 0 12972 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1644511149
transform 1 0 14720 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0834_
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0835_
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1644511149
transform 1 0 16744 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0837_
timestamp 1644511149
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0839_
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1644511149
transform 1 0 15364 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0844_
timestamp 1644511149
transform 1 0 16836 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1644511149
transform 1 0 18124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0846_
timestamp 1644511149
transform 1 0 18584 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0847_
timestamp 1644511149
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0848_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1644511149
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0850_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0853_
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0854_
timestamp 1644511149
transform 1 0 19872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1644511149
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0857_
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0858_
timestamp 1644511149
transform 1 0 21896 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1644511149
transform 1 0 22632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1644511149
transform 1 0 21068 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0861_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0862_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0864_
timestamp 1644511149
transform 1 0 16468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1644511149
transform 1 0 7360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0876_
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0882_
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0889_
timestamp 1644511149
transform 1 0 24564 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform 1 0 42780 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 41400 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0901_
timestamp 1644511149
transform 1 0 24564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 45908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0907_
timestamp 1644511149
transform 1 0 23368 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 46736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0913_
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 22908 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0919_
timestamp 1644511149
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0920_
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 8096 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1644511149
transform 1 0 8188 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0926_
timestamp 1644511149
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1644511149
transform 1 0 27968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0932_
timestamp 1644511149
transform 1 0 26128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 40664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1644511149
transform 1 0 27048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0938_
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0944_
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0951_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 46644 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 2852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 33120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0957_
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 42688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0963_
timestamp 1644511149
transform 1 0 20700 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 46736 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0969_
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 19320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0975_
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 16744 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0982_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0983_
timestamp 1644511149
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 20148 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _0985_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0988_
timestamp 1644511149
transform 1 0 26036 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0989_
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0991_
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0992_
timestamp 1644511149
transform 1 0 23460 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _0994_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0996_
timestamp 1644511149
transform 1 0 27508 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0997_
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0998_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0999_
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1000_
timestamp 1644511149
transform 1 0 43240 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29992 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1003_
timestamp 1644511149
transform 1 0 44252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1004_
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1005_
timestamp 1644511149
transform 1 0 45908 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1644511149
transform 1 0 44160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44528 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1644511149
transform 1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1011_
timestamp 1644511149
transform 1 0 44252 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _1012_
timestamp 1644511149
transform 1 0 43976 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1013_
timestamp 1644511149
transform 1 0 43332 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1644511149
transform 1 0 43608 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1644511149
transform 1 0 45264 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1644511149
transform 1 0 42780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1018_
timestamp 1644511149
transform 1 0 45816 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _1019_
timestamp 1644511149
transform 1 0 43792 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1644511149
transform 1 0 43148 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1021_
timestamp 1644511149
transform 1 0 43424 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1022_
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 20792 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1024_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1026_
timestamp 1644511149
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1028_
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1029_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 17572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1031_
timestamp 1644511149
transform 1 0 15824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1032_
timestamp 1644511149
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1033_
timestamp 1644511149
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1034_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1035_
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1036_
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1037_
timestamp 1644511149
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1039_
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1040_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1042_
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1043_
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 12972 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1045_
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1046_
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1047_
timestamp 1644511149
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1048_
timestamp 1644511149
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1049_
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1050_
timestamp 1644511149
transform 1 0 14168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1051_
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1052_
timestamp 1644511149
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1053_
timestamp 1644511149
transform 1 0 16836 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1054_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1055_
timestamp 1644511149
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1056_
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1059_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1063_
timestamp 1644511149
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1644511149
transform 1 0 32200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform 1 0 33120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1644511149
transform 1 0 32200 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1644511149
transform 1 0 33304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1069_
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1644511149
transform 1 0 32752 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1644511149
transform 1 0 19780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1075_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1644511149
transform 1 0 26956 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1081_
timestamp 1644511149
transform 1 0 23736 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1644511149
transform 1 0 31096 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1644511149
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1087_
timestamp 1644511149
transform 1 0 22724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1644511149
transform 1 0 23552 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1644511149
transform 1 0 22448 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1093_
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1644511149
transform 1 0 15272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1102_
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1103_
timestamp 1644511149
transform 1 0 19136 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1644511149
transform 1 0 16376 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1105_
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1644511149
transform 1 0 13800 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1108_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1644511149
transform 1 0 14628 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1112_
timestamp 1644511149
transform 1 0 9936 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1644511149
transform 1 0 9476 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1115_
timestamp 1644511149
transform 1 0 10212 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1116_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1117_
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1644511149
transform 1 0 9476 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1120_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1121_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1644511149
transform 1 0 14628 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1644511149
transform 1 0 16744 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1644511149
transform 1 0 18952 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1128_
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1133_
timestamp 1644511149
transform 1 0 28152 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1644511149
transform 1 0 31096 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1644511149
transform 1 0 32200 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1644511149
transform 1 0 31004 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1644511149
transform 1 0 32568 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1644511149
transform 1 0 32200 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1140_
timestamp 1644511149
transform 1 0 18768 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1644511149
transform 1 0 19780 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1644511149
transform 1 0 25392 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1147_
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1644511149
transform 1 0 31188 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1644511149
transform 1 0 28244 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1644511149
transform 1 0 24196 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1644511149
transform 1 0 26128 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1644511149
transform 1 0 22632 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1155_
timestamp 1644511149
transform 1 0 24380 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1644511149
transform 1 0 20148 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1644511149
transform 1 0 16928 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1644511149
transform 1 0 14904 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1644511149
transform 1 0 14720 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _1164__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__83
timestamp 1644511149
transform 1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__84
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__85
timestamp 1644511149
transform 1 0 37076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__86
timestamp 1644511149
transform 1 0 20700 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__87
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__88
timestamp 1644511149
transform 1 0 24564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__90
timestamp 1644511149
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__91
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__92
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__93
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__94
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__95
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__96
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__98
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__99
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__100
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1184__101
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185__102
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1186__103
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1187__104
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1188__105
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1189__106
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1190__107
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1191__108
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1192__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1193__110
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1194__111
timestamp 1644511149
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1195__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1196__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1197__114
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1198__115
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1199__116
timestamp 1644511149
transform 1 0 42688 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1201__118
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1202__119
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1203__120
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1204__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1205__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1206__123
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1207__124
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1208__125
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1209__126
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1210__127
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1211__128
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1212__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1213__130
timestamp 1644511149
transform 1 0 46092 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1214__131
timestamp 1644511149
transform 1 0 1840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1215__132
timestamp 1644511149
transform 1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1216__133
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1217__134
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1218__135
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1220_
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1224_
timestamp 1644511149
transform 1 0 40572 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1225_
timestamp 1644511149
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1226_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1227_
timestamp 1644511149
transform 1 0 25760 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1228_
timestamp 1644511149
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1229_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1230_
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1231_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1232_
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1233_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1234_
timestamp 1644511149
transform 1 0 10672 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1235_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1236_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1237_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1238_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1239_
timestamp 1644511149
transform 1 0 2024 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1240_
timestamp 1644511149
transform 1 0 33028 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1241_
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1242_
timestamp 1644511149
transform 1 0 2024 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1243_
timestamp 1644511149
transform 1 0 42596 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1244_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1245_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1246_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1247_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1248_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1249_
timestamp 1644511149
transform 1 0 7912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1250_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1251_
timestamp 1644511149
transform 1 0 22816 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1252_
timestamp 1644511149
transform 1 0 25300 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1253_
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1254_
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1255_
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1256_
timestamp 1644511149
transform 1 0 19412 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1257_
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1258_
timestamp 1644511149
transform 1 0 14168 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1259_
timestamp 1644511149
transform 1 0 15364 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1260_
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1261_
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1262_
timestamp 1644511149
transform 1 0 7912 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1263_
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1264_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1265_
timestamp 1644511149
transform 1 0 8004 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1266_
timestamp 1644511149
transform 1 0 7912 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1267_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1268_
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1269_
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1270_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1271_
timestamp 1644511149
transform 1 0 7728 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1272_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1273_
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1274_
timestamp 1644511149
transform 1 0 8372 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1275_
timestamp 1644511149
transform 1 0 17940 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1276_
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1277_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1644511149
transform 1 0 23000 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1644511149
transform 1 0 23276 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1644511149
transform 1 0 41308 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24748 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22080 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 47656 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 2944 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 47288 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 47932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1644511149
transform 1 0 46184 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 46184 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 2024 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1644511149
transform 1 0 47288 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 47656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 43792 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 47288 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 41308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 38916 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 39100 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 28244 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 29440 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 15272 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 22816 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1840 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45356 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 45816 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 43056 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 27140 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 25852 0 1 21760
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
