magic
tech sky130A
magscale 1 2
timestamp 1654174654
<< viali >>
rect 12449 47141 12483 47175
rect 19441 47141 19475 47175
rect 29929 47141 29963 47175
rect 20085 47073 20119 47107
rect 30757 47073 30791 47107
rect 43177 47073 43211 47107
rect 47041 47073 47075 47107
rect 1961 47005 1995 47039
rect 2697 47005 2731 47039
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6837 47005 6871 47039
rect 7757 47005 7791 47039
rect 9137 47005 9171 47039
rect 11621 47005 11655 47039
rect 12265 47005 12299 47039
rect 13093 47005 13127 47039
rect 14565 47005 14599 47039
rect 19257 47005 19291 47039
rect 20361 47005 20395 47039
rect 24869 47005 24903 47039
rect 25513 47005 25547 47039
rect 28641 47005 28675 47039
rect 29745 47005 29779 47039
rect 31033 47005 31067 47039
rect 38301 47005 38335 47039
rect 42625 47005 42659 47039
rect 45201 47005 45235 47039
rect 47777 47005 47811 47039
rect 4077 46937 4111 46971
rect 4997 46937 5031 46971
rect 7941 46937 7975 46971
rect 11805 46937 11839 46971
rect 13461 46937 13495 46971
rect 14749 46937 14783 46971
rect 17141 46937 17175 46971
rect 17325 46937 17359 46971
rect 40325 46937 40359 46971
rect 40509 46937 40543 46971
rect 42809 46937 42843 46971
rect 45385 46937 45419 46971
rect 2145 46869 2179 46903
rect 2881 46869 2915 46903
rect 6929 46869 6963 46903
rect 9321 46869 9355 46903
rect 28457 46869 28491 46903
rect 47961 46869 47995 46903
rect 28365 46597 28399 46631
rect 1409 46529 1443 46563
rect 24593 46529 24627 46563
rect 28181 46529 28215 46563
rect 38117 46529 38151 46563
rect 47869 46529 47903 46563
rect 3985 46461 4019 46495
rect 4169 46461 4203 46495
rect 5181 46461 5215 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 12449 46461 12483 46495
rect 13829 46461 13863 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 19257 46461 19291 46495
rect 19441 46461 19475 46495
rect 20637 46461 20671 46495
rect 24777 46461 24811 46495
rect 25145 46461 25179 46495
rect 29377 46461 29411 46495
rect 31585 46461 31619 46495
rect 32137 46461 32171 46495
rect 32321 46461 32355 46495
rect 32597 46461 32631 46495
rect 38301 46461 38335 46495
rect 38669 46461 38703 46495
rect 41889 46461 41923 46495
rect 42441 46461 42475 46495
rect 42625 46461 42659 46495
rect 42901 46461 42935 46495
rect 45201 46461 45235 46495
rect 45385 46461 45419 46495
rect 46857 46461 46891 46495
rect 1593 46325 1627 46359
rect 22017 46325 22051 46359
rect 41245 46325 41279 46359
rect 48053 46325 48087 46359
rect 4445 46121 4479 46155
rect 5089 46121 5123 46155
rect 12173 46121 12207 46155
rect 13553 46121 13587 46155
rect 14197 46121 14231 46155
rect 18613 46121 18647 46155
rect 19441 46121 19475 46155
rect 24685 46121 24719 46155
rect 31861 46121 31895 46155
rect 38301 46121 38335 46155
rect 20729 45985 20763 46019
rect 21281 45985 21315 46019
rect 25237 45985 25271 46019
rect 25789 45985 25823 46019
rect 41245 45985 41279 46019
rect 41889 45985 41923 46019
rect 47041 45985 47075 46019
rect 2053 45917 2087 45951
rect 4997 45917 5031 45951
rect 12081 45917 12115 45951
rect 14105 45917 14139 45951
rect 18521 45917 18555 45951
rect 24593 45917 24627 45951
rect 31769 45917 31803 45951
rect 38209 45917 38243 45951
rect 44005 45917 44039 45951
rect 45569 45917 45603 45951
rect 46305 45917 46339 45951
rect 20913 45849 20947 45883
rect 25421 45849 25455 45883
rect 41429 45849 41463 45883
rect 44189 45849 44223 45883
rect 46489 45849 46523 45883
rect 45753 45781 45787 45815
rect 20913 45577 20947 45611
rect 25421 45577 25455 45611
rect 41429 45577 41463 45611
rect 42533 45577 42567 45611
rect 43177 45509 43211 45543
rect 43913 45509 43947 45543
rect 46949 45509 46983 45543
rect 1777 45441 1811 45475
rect 20821 45441 20855 45475
rect 25329 45441 25363 45475
rect 41337 45441 41371 45475
rect 42441 45441 42475 45475
rect 43085 45441 43119 45475
rect 46857 45441 46891 45475
rect 47593 45441 47627 45475
rect 1961 45373 1995 45407
rect 2789 45373 2823 45407
rect 44557 45373 44591 45407
rect 44741 45373 44775 45407
rect 45569 45373 45603 45407
rect 44005 45237 44039 45271
rect 47777 45237 47811 45271
rect 2237 45033 2271 45067
rect 42993 45033 43027 45067
rect 44465 45033 44499 45067
rect 45109 45033 45143 45067
rect 45753 45033 45787 45067
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 2145 44829 2179 44863
rect 45017 44829 45051 44863
rect 45661 44829 45695 44863
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 47685 44489 47719 44523
rect 44833 44353 44867 44387
rect 45753 44353 45787 44387
rect 46213 44353 46247 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 46949 44149 46983 44183
rect 46489 43809 46523 43843
rect 48145 43809 48179 43843
rect 45845 43741 45879 43775
rect 46305 43741 46339 43775
rect 1409 43265 1443 43299
rect 47041 43265 47075 43299
rect 47777 43265 47811 43299
rect 1685 43197 1719 43231
rect 46305 42653 46339 42687
rect 46489 42585 46523 42619
rect 48145 42585 48179 42619
rect 47685 42313 47719 42347
rect 47041 42177 47075 42211
rect 47593 42177 47627 42211
rect 2053 41973 2087 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 27353 41565 27387 41599
rect 48145 41565 48179 41599
rect 1593 41497 1627 41531
rect 46489 41497 46523 41531
rect 27445 41429 27479 41463
rect 2145 41225 2179 41259
rect 46765 41225 46799 41259
rect 27169 41157 27203 41191
rect 28825 41157 28859 41191
rect 2053 41089 2087 41123
rect 46673 41089 46707 41123
rect 47777 41089 47811 41123
rect 26985 41021 27019 41055
rect 46857 40613 46891 40647
rect 26065 40545 26099 40579
rect 1409 40477 1443 40511
rect 45109 40477 45143 40511
rect 45477 40477 45511 40511
rect 47041 40477 47075 40511
rect 47685 40477 47719 40511
rect 26249 40409 26283 40443
rect 27905 40409 27939 40443
rect 1593 40341 1627 40375
rect 46121 40341 46155 40375
rect 45845 40001 45879 40035
rect 46121 40001 46155 40035
rect 47593 40001 47627 40035
rect 46121 39865 46155 39899
rect 47685 39797 47719 39831
rect 46305 39457 46339 39491
rect 46489 39457 46523 39491
rect 48145 39457 48179 39491
rect 45201 39049 45235 39083
rect 45017 38913 45051 38947
rect 45845 38913 45879 38947
rect 47869 38913 47903 38947
rect 46397 38845 46431 38879
rect 48053 38777 48087 38811
rect 45569 38369 45603 38403
rect 45201 38301 45235 38335
rect 46305 38301 46339 38335
rect 46489 38233 46523 38267
rect 48145 38233 48179 38267
rect 47685 37961 47719 37995
rect 45845 37825 45879 37859
rect 47593 37825 47627 37859
rect 46213 37757 46247 37791
rect 47685 37417 47719 37451
rect 2053 37213 2087 37247
rect 45845 37213 45879 37247
rect 46397 37145 46431 37179
rect 46397 36805 46431 36839
rect 1777 36737 1811 36771
rect 45845 36737 45879 36771
rect 1961 36669 1995 36703
rect 2789 36669 2823 36703
rect 2237 36329 2271 36363
rect 2145 36125 2179 36159
rect 1593 35649 1627 35683
rect 1409 35445 1443 35479
rect 48145 35037 48179 35071
rect 47961 34901 47995 34935
rect 29561 34561 29595 34595
rect 30573 34561 30607 34595
rect 48145 34561 48179 34595
rect 29653 34493 29687 34527
rect 30389 34357 30423 34391
rect 47961 34357 47995 34391
rect 24961 34017 24995 34051
rect 30021 34017 30055 34051
rect 47133 34017 47167 34051
rect 47409 34017 47443 34051
rect 1593 33949 1627 33983
rect 20545 33949 20579 33983
rect 20821 33881 20855 33915
rect 24869 33881 24903 33915
rect 30297 33881 30331 33915
rect 47225 33881 47259 33915
rect 1409 33813 1443 33847
rect 22293 33813 22327 33847
rect 24409 33813 24443 33847
rect 24777 33813 24811 33847
rect 31769 33813 31803 33847
rect 30481 33609 30515 33643
rect 31217 33609 31251 33643
rect 31309 33609 31343 33643
rect 32689 33609 32723 33643
rect 22385 33541 22419 33575
rect 19349 33473 19383 33507
rect 21281 33473 21315 33507
rect 23489 33473 23523 33507
rect 30021 33473 30055 33507
rect 30205 33473 30239 33507
rect 32321 33473 32355 33507
rect 47777 33473 47811 33507
rect 1409 33405 1443 33439
rect 1685 33405 1719 33439
rect 22477 33405 22511 33439
rect 22661 33405 22695 33439
rect 23949 33405 23983 33439
rect 24225 33405 24259 33439
rect 27905 33405 27939 33439
rect 28181 33405 28215 33439
rect 31493 33405 31527 33439
rect 32229 33405 32263 33439
rect 19441 33269 19475 33303
rect 21097 33269 21131 33303
rect 22017 33269 22051 33303
rect 23305 33269 23339 33303
rect 25697 33269 25731 33303
rect 29653 33269 29687 33303
rect 30021 33269 30055 33303
rect 30849 33269 30883 33303
rect 47869 33269 47903 33303
rect 18613 33065 18647 33099
rect 21649 33065 21683 33099
rect 24409 33065 24443 33099
rect 25697 33065 25731 33099
rect 28641 33065 28675 33099
rect 30573 33065 30607 33099
rect 31861 33065 31895 33099
rect 35725 32997 35759 33031
rect 1409 32929 1443 32963
rect 1593 32929 1627 32963
rect 22109 32929 22143 32963
rect 22293 32929 22327 32963
rect 24961 32929 24995 32963
rect 28273 32929 28307 32963
rect 31033 32929 31067 32963
rect 31217 32929 31251 32963
rect 36369 32929 36403 32963
rect 12449 32861 12483 32895
rect 12633 32861 12667 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 22845 32861 22879 32895
rect 23581 32861 23615 32895
rect 24777 32861 24811 32895
rect 24869 32861 24903 32895
rect 25605 32861 25639 32895
rect 27905 32861 27939 32895
rect 28089 32861 28123 32895
rect 28181 32861 28215 32895
rect 28457 32861 28491 32895
rect 29745 32861 29779 32895
rect 29929 32861 29963 32895
rect 30021 32861 30055 32895
rect 30941 32861 30975 32895
rect 31769 32861 31803 32895
rect 32689 32861 32723 32895
rect 33609 32861 33643 32895
rect 36093 32861 36127 32895
rect 46305 32861 46339 32895
rect 3249 32793 3283 32827
rect 19441 32793 19475 32827
rect 21097 32793 21131 32827
rect 46489 32793 46523 32827
rect 48145 32793 48179 32827
rect 12541 32725 12575 32759
rect 22017 32725 22051 32759
rect 23029 32725 23063 32759
rect 23765 32725 23799 32759
rect 29561 32725 29595 32759
rect 32873 32725 32907 32759
rect 33425 32725 33459 32759
rect 36185 32725 36219 32759
rect 22385 32521 22419 32555
rect 24869 32521 24903 32555
rect 29009 32521 29043 32555
rect 35725 32521 35759 32555
rect 46857 32521 46891 32555
rect 47685 32521 47719 32555
rect 2329 32453 2363 32487
rect 19349 32453 19383 32487
rect 21005 32453 21039 32487
rect 32505 32453 32539 32487
rect 34805 32453 34839 32487
rect 11713 32385 11747 32419
rect 12817 32385 12851 32419
rect 14657 32385 14691 32419
rect 15669 32385 15703 32419
rect 16681 32385 16715 32419
rect 22017 32385 22051 32419
rect 24501 32385 24535 32419
rect 25329 32385 25363 32419
rect 28457 32385 28491 32419
rect 28825 32385 28859 32419
rect 29929 32385 29963 32419
rect 30113 32385 30147 32419
rect 32229 32385 32263 32419
rect 36093 32385 36127 32419
rect 37473 32385 37507 32419
rect 47041 32385 47075 32419
rect 47593 32385 47627 32419
rect 2145 32317 2179 32351
rect 3249 32317 3283 32351
rect 12909 32317 12943 32351
rect 19165 32317 19199 32351
rect 21925 32317 21959 32351
rect 24593 32317 24627 32351
rect 34897 32317 34931 32351
rect 34989 32317 35023 32351
rect 36185 32317 36219 32351
rect 36369 32317 36403 32351
rect 34437 32249 34471 32283
rect 1685 32181 1719 32215
rect 11713 32181 11747 32215
rect 13185 32181 13219 32215
rect 14749 32181 14783 32215
rect 15485 32181 15519 32215
rect 16773 32181 16807 32215
rect 25513 32181 25547 32215
rect 28825 32181 28859 32215
rect 30297 32181 30331 32215
rect 33977 32181 34011 32215
rect 37289 32181 37323 32215
rect 14289 31977 14323 32011
rect 14473 31977 14507 32011
rect 21649 31977 21683 32011
rect 32781 31977 32815 32011
rect 34069 31977 34103 32011
rect 37565 31977 37599 32011
rect 47685 31977 47719 32011
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 11713 31841 11747 31875
rect 11989 31841 12023 31875
rect 15209 31841 15243 31875
rect 15485 31841 15519 31875
rect 16957 31841 16991 31875
rect 18061 31841 18095 31875
rect 18613 31841 18647 31875
rect 19441 31841 19475 31875
rect 19717 31841 19751 31875
rect 27261 31841 27295 31875
rect 27537 31841 27571 31875
rect 33333 31841 33367 31875
rect 35817 31841 35851 31875
rect 36093 31841 36127 31875
rect 17601 31773 17635 31807
rect 17693 31773 17727 31807
rect 18521 31773 18555 31807
rect 19257 31773 19291 31807
rect 21557 31773 21591 31807
rect 25605 31773 25639 31807
rect 33977 31773 34011 31807
rect 1593 31705 1627 31739
rect 14105 31705 14139 31739
rect 14321 31705 14355 31739
rect 17969 31705 18003 31739
rect 33241 31705 33275 31739
rect 13461 31637 13495 31671
rect 17417 31637 17451 31671
rect 17785 31637 17819 31671
rect 25697 31637 25731 31671
rect 29009 31637 29043 31671
rect 33149 31637 33183 31671
rect 2237 31433 2271 31467
rect 11621 31433 11655 31467
rect 12357 31433 12391 31467
rect 14657 31433 14691 31467
rect 15761 31433 15795 31467
rect 16957 31433 16991 31467
rect 27353 31433 27387 31467
rect 28641 31433 28675 31467
rect 36645 31433 36679 31467
rect 37381 31433 37415 31467
rect 12173 31365 12207 31399
rect 13185 31365 13219 31399
rect 16681 31365 16715 31399
rect 29469 31365 29503 31399
rect 2145 31297 2179 31331
rect 9137 31297 9171 31331
rect 10057 31297 10091 31331
rect 10701 31297 10735 31331
rect 11529 31297 11563 31331
rect 12449 31297 12483 31331
rect 15577 31297 15611 31331
rect 16865 31297 16899 31331
rect 17049 31297 17083 31331
rect 22293 31297 22327 31331
rect 22477 31297 22511 31331
rect 24593 31297 24627 31331
rect 27261 31297 27295 31331
rect 27905 31297 27939 31331
rect 28089 31297 28123 31331
rect 28181 31297 28215 31331
rect 28457 31297 28491 31331
rect 29285 31297 29319 31331
rect 33609 31297 33643 31331
rect 36553 31297 36587 31331
rect 36737 31297 36771 31331
rect 37289 31297 37323 31331
rect 9229 31229 9263 31263
rect 12909 31229 12943 31263
rect 15393 31229 15427 31263
rect 17877 31229 17911 31263
rect 18153 31229 18187 31263
rect 19625 31229 19659 31263
rect 22569 31229 22603 31263
rect 24869 31229 24903 31263
rect 28273 31229 28307 31263
rect 29101 31229 29135 31263
rect 33517 31229 33551 31263
rect 33977 31229 34011 31263
rect 12173 31161 12207 31195
rect 9505 31093 9539 31127
rect 10149 31093 10183 31127
rect 10793 31093 10827 31127
rect 17233 31093 17267 31127
rect 22109 31093 22143 31127
rect 26341 31093 26375 31127
rect 12909 30889 12943 30923
rect 14197 30889 14231 30923
rect 18061 30889 18095 30923
rect 19349 30889 19383 30923
rect 23397 30889 23431 30923
rect 25697 30889 25731 30923
rect 26525 30889 26559 30923
rect 27813 30889 27847 30923
rect 28181 30889 28215 30923
rect 29653 30889 29687 30923
rect 31033 30889 31067 30923
rect 32965 30889 32999 30923
rect 33701 30889 33735 30923
rect 36185 30889 36219 30923
rect 18613 30821 18647 30855
rect 31217 30821 31251 30855
rect 9689 30753 9723 30787
rect 9965 30753 9999 30787
rect 17601 30753 17635 30787
rect 20453 30753 20487 30787
rect 20729 30753 20763 30787
rect 22931 30753 22965 30787
rect 12909 30685 12943 30719
rect 14105 30685 14139 30719
rect 15669 30685 15703 30719
rect 16129 30685 16163 30719
rect 16313 30685 16347 30719
rect 17693 30685 17727 30719
rect 18521 30685 18555 30719
rect 19257 30685 19291 30719
rect 22661 30685 22695 30719
rect 22845 30685 22879 30719
rect 23029 30685 23063 30719
rect 23213 30685 23247 30719
rect 24961 30685 24995 30719
rect 25145 30685 25179 30719
rect 25237 30685 25271 30719
rect 25329 30685 25363 30719
rect 25513 30685 25547 30719
rect 27813 30685 27847 30719
rect 27997 30685 28031 30719
rect 28641 30685 28675 30719
rect 29561 30685 29595 30719
rect 29745 30685 29779 30719
rect 30849 30685 30883 30719
rect 31033 30685 31067 30719
rect 32321 30685 32355 30719
rect 32505 30685 32539 30719
rect 32965 30685 32999 30719
rect 33149 30685 33183 30719
rect 33609 30685 33643 30719
rect 36093 30685 36127 30719
rect 36277 30685 36311 30719
rect 36921 30685 36955 30719
rect 11713 30617 11747 30651
rect 15485 30617 15519 30651
rect 26249 30617 26283 30651
rect 28825 30617 28859 30651
rect 32413 30617 32447 30651
rect 36737 30617 36771 30651
rect 16221 30549 16255 30583
rect 22201 30549 22235 30583
rect 29009 30549 29043 30583
rect 34069 30549 34103 30583
rect 37105 30549 37139 30583
rect 17509 30345 17543 30379
rect 22569 30345 22603 30379
rect 26065 30345 26099 30379
rect 17233 30277 17267 30311
rect 21189 30277 21223 30311
rect 23029 30277 23063 30311
rect 24777 30277 24811 30311
rect 30021 30277 30055 30311
rect 31309 30277 31343 30311
rect 9873 30209 9907 30243
rect 13001 30209 13035 30243
rect 17141 30209 17175 30243
rect 17325 30209 17359 30243
rect 21097 30209 21131 30243
rect 22017 30209 22051 30243
rect 22385 30209 22419 30243
rect 23213 30209 23247 30243
rect 23949 30209 23983 30243
rect 24133 30209 24167 30243
rect 24961 30209 24995 30243
rect 25697 30209 25731 30243
rect 25881 30209 25915 30243
rect 28641 30209 28675 30243
rect 30297 30209 30331 30243
rect 31125 30209 31159 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 37473 30209 37507 30243
rect 38485 30209 38519 30243
rect 13185 30141 13219 30175
rect 13461 30141 13495 30175
rect 25237 30141 25271 30175
rect 28457 30141 28491 30175
rect 30205 30141 30239 30175
rect 33517 30141 33551 30175
rect 33793 30141 33827 30175
rect 37381 30141 37415 30175
rect 38301 30141 38335 30175
rect 16957 30073 16991 30107
rect 25145 30073 25179 30107
rect 9965 30005 9999 30039
rect 22109 30005 22143 30039
rect 23397 30005 23431 30039
rect 24133 30005 24167 30039
rect 24317 30005 24351 30039
rect 25881 30005 25915 30039
rect 28825 30005 28859 30039
rect 30021 30005 30055 30039
rect 30481 30005 30515 30039
rect 31493 30005 31527 30039
rect 32229 30005 32263 30039
rect 35265 30005 35299 30039
rect 37749 30005 37783 30039
rect 38669 30005 38703 30039
rect 12541 29801 12575 29835
rect 13277 29801 13311 29835
rect 23397 29801 23431 29835
rect 24593 29801 24627 29835
rect 25421 29801 25455 29835
rect 27524 29801 27558 29835
rect 29009 29801 29043 29835
rect 31309 29801 31343 29835
rect 31677 29801 31711 29835
rect 33977 29801 34011 29835
rect 35357 29801 35391 29835
rect 36001 29801 36035 29835
rect 36921 29801 36955 29835
rect 17233 29665 17267 29699
rect 17693 29665 17727 29699
rect 23489 29665 23523 29699
rect 27261 29665 27295 29699
rect 31401 29665 31435 29699
rect 32413 29665 32447 29699
rect 36185 29665 36219 29699
rect 36829 29665 36863 29699
rect 37565 29665 37599 29699
rect 47593 29665 47627 29699
rect 8401 29597 8435 29631
rect 8953 29597 8987 29631
rect 11437 29597 11471 29631
rect 12449 29597 12483 29631
rect 13093 29597 13127 29631
rect 14289 29597 14323 29631
rect 15853 29597 15887 29631
rect 17325 29597 17359 29631
rect 18153 29597 18187 29631
rect 19257 29597 19291 29631
rect 22477 29597 22511 29631
rect 22661 29597 22695 29631
rect 23305 29597 23339 29631
rect 23581 29597 23615 29631
rect 24409 29597 24443 29631
rect 24501 29597 24535 29631
rect 25329 29597 25363 29631
rect 25513 29597 25547 29631
rect 26525 29597 26559 29631
rect 31309 29597 31343 29631
rect 32229 29597 32263 29631
rect 32873 29597 32907 29631
rect 33149 29597 33183 29631
rect 33885 29597 33919 29631
rect 34713 29597 34747 29631
rect 34806 29597 34840 29631
rect 35081 29597 35115 29631
rect 35178 29597 35212 29631
rect 35909 29597 35943 29631
rect 36921 29597 36955 29631
rect 47317 29597 47351 29631
rect 9229 29529 9263 29563
rect 14565 29529 14599 29563
rect 30021 29529 30055 29563
rect 33057 29529 33091 29563
rect 34989 29529 35023 29563
rect 36645 29529 36679 29563
rect 37841 29529 37875 29563
rect 8217 29461 8251 29495
rect 10701 29461 10735 29495
rect 11529 29461 11563 29495
rect 15945 29461 15979 29495
rect 18337 29461 18371 29495
rect 19349 29461 19383 29495
rect 22569 29461 22603 29495
rect 23765 29461 23799 29495
rect 24777 29461 24811 29495
rect 26617 29461 26651 29495
rect 30113 29461 30147 29495
rect 32965 29461 32999 29495
rect 36185 29461 36219 29495
rect 37105 29461 37139 29495
rect 39313 29461 39347 29495
rect 9229 29257 9263 29291
rect 11989 29257 12023 29291
rect 19717 29257 19751 29291
rect 20729 29257 20763 29291
rect 22937 29257 22971 29291
rect 25237 29257 25271 29291
rect 28733 29257 28767 29291
rect 8217 29189 8251 29223
rect 14841 29189 14875 29223
rect 18245 29189 18279 29223
rect 26249 29189 26283 29223
rect 29929 29189 29963 29223
rect 30573 29189 30607 29223
rect 34989 29189 35023 29223
rect 38485 29189 38519 29223
rect 7941 29121 7975 29155
rect 8769 29121 8803 29155
rect 10425 29121 10459 29155
rect 11805 29121 11839 29155
rect 15485 29121 15519 29155
rect 17233 29121 17267 29155
rect 17969 29121 18003 29155
rect 20545 29121 20579 29155
rect 22293 29121 22327 29155
rect 23121 29121 23155 29155
rect 24869 29121 24903 29155
rect 24961 29121 24995 29155
rect 27353 29121 27387 29155
rect 27537 29119 27571 29153
rect 27997 29121 28031 29155
rect 28181 29121 28215 29155
rect 28273 29121 28307 29155
rect 28549 29121 28583 29155
rect 29745 29121 29779 29155
rect 30849 29121 30883 29155
rect 32689 29121 32723 29155
rect 34897 29121 34931 29155
rect 36001 29121 36035 29155
rect 37289 29121 37323 29155
rect 37437 29121 37471 29155
rect 37565 29121 37599 29155
rect 37657 29121 37691 29155
rect 37795 29121 37829 29155
rect 38393 29121 38427 29155
rect 13001 29053 13035 29087
rect 13185 29053 13219 29087
rect 15577 29053 15611 29087
rect 17141 29053 17175 29087
rect 17325 29053 17359 29087
rect 17417 29053 17451 29087
rect 23581 29053 23615 29087
rect 23857 29053 23891 29087
rect 27445 29053 27479 29087
rect 28365 29053 28399 29087
rect 30757 29053 30791 29087
rect 34437 29053 34471 29087
rect 35725 29053 35759 29087
rect 9045 28985 9079 29019
rect 26433 28985 26467 29019
rect 30113 28985 30147 29019
rect 31033 28985 31067 29019
rect 37933 28985 37967 29019
rect 10425 28917 10459 28951
rect 15761 28917 15795 28951
rect 16957 28917 16991 28951
rect 22385 28917 22419 28951
rect 24869 28917 24903 28951
rect 30849 28917 30883 28951
rect 32946 28917 32980 28951
rect 12173 28713 12207 28747
rect 12725 28713 12759 28747
rect 16405 28713 16439 28747
rect 24501 28713 24535 28747
rect 26985 28713 27019 28747
rect 28457 28713 28491 28747
rect 30849 28713 30883 28747
rect 31033 28713 31067 28747
rect 32413 28713 32447 28747
rect 33793 28713 33827 28747
rect 38853 28713 38887 28747
rect 17417 28645 17451 28679
rect 9505 28577 9539 28611
rect 10425 28577 10459 28611
rect 14657 28577 14691 28611
rect 14933 28577 14967 28611
rect 17141 28577 17175 28611
rect 24685 28577 24719 28611
rect 30757 28577 30791 28611
rect 36461 28577 36495 28611
rect 38485 28577 38519 28611
rect 46489 28577 46523 28611
rect 47041 28577 47075 28611
rect 9597 28509 9631 28543
rect 12633 28509 12667 28543
rect 13369 28509 13403 28543
rect 18061 28509 18095 28543
rect 18245 28509 18279 28543
rect 20177 28509 20211 28543
rect 22753 28509 22787 28543
rect 22845 28509 22879 28543
rect 22937 28509 22971 28543
rect 23121 28509 23155 28543
rect 23673 28509 23707 28543
rect 23857 28509 23891 28543
rect 24409 28509 24443 28543
rect 25237 28509 25271 28543
rect 27629 28509 27663 28543
rect 28365 28509 28399 28543
rect 29653 28509 29687 28543
rect 29745 28509 29779 28543
rect 30573 28509 30607 28543
rect 30849 28509 30883 28543
rect 31677 28509 31711 28543
rect 31861 28509 31895 28543
rect 31953 28509 31987 28543
rect 32091 28509 32125 28543
rect 32229 28509 32263 28543
rect 33057 28509 33091 28543
rect 35173 28509 35207 28543
rect 35357 28509 35391 28543
rect 38669 28509 38703 28543
rect 46305 28509 46339 28543
rect 10701 28441 10735 28475
rect 18429 28441 18463 28475
rect 20361 28441 20395 28475
rect 22017 28441 22051 28475
rect 24685 28441 24719 28475
rect 25513 28441 25547 28475
rect 27813 28441 27847 28475
rect 29929 28441 29963 28475
rect 33701 28441 33735 28475
rect 36185 28441 36219 28475
rect 9965 28373 9999 28407
rect 13461 28373 13495 28407
rect 17601 28373 17635 28407
rect 22477 28373 22511 28407
rect 23857 28373 23891 28407
rect 32873 28373 32907 28407
rect 35357 28373 35391 28407
rect 35817 28373 35851 28407
rect 36277 28373 36311 28407
rect 15945 28169 15979 28203
rect 17157 28169 17191 28203
rect 17325 28169 17359 28203
rect 20269 28169 20303 28203
rect 25881 28169 25915 28203
rect 36093 28169 36127 28203
rect 16957 28101 16991 28135
rect 18061 28101 18095 28135
rect 22109 28101 22143 28135
rect 27445 28101 27479 28135
rect 32781 28101 32815 28135
rect 7941 28033 7975 28067
rect 11529 28033 11563 28067
rect 15761 28033 15795 28067
rect 20177 28033 20211 28067
rect 21833 28033 21867 28067
rect 24041 28033 24075 28067
rect 24225 28033 24259 28067
rect 24317 28033 24351 28067
rect 24501 28033 24535 28067
rect 24593 28033 24627 28067
rect 25237 28033 25271 28067
rect 25330 28033 25364 28067
rect 25513 28033 25547 28067
rect 25605 28033 25639 28067
rect 25743 28033 25777 28067
rect 27629 28033 27663 28067
rect 29745 28033 29779 28067
rect 30941 28033 30975 28067
rect 31125 28033 31159 28067
rect 31217 28033 31251 28067
rect 33609 28033 33643 28067
rect 36001 28033 36035 28067
rect 37473 28033 37507 28067
rect 37933 28033 37967 28067
rect 47593 28033 47627 28067
rect 8125 27965 8159 27999
rect 8401 27965 8435 27999
rect 12725 27965 12759 27999
rect 12909 27965 12943 27999
rect 13185 27965 13219 27999
rect 17785 27965 17819 27999
rect 19533 27965 19567 27999
rect 23581 27965 23615 27999
rect 30021 27965 30055 27999
rect 36185 27965 36219 27999
rect 29929 27897 29963 27931
rect 32965 27897 32999 27931
rect 35633 27897 35667 27931
rect 11713 27829 11747 27863
rect 17141 27829 17175 27863
rect 29837 27829 29871 27863
rect 31217 27829 31251 27863
rect 31401 27829 31435 27863
rect 33425 27829 33459 27863
rect 37289 27829 37323 27863
rect 38025 27829 38059 27863
rect 47041 27829 47075 27863
rect 47685 27829 47719 27863
rect 7665 27625 7699 27659
rect 13185 27625 13219 27659
rect 23581 27625 23615 27659
rect 32137 27625 32171 27659
rect 36356 27625 36390 27659
rect 9045 27557 9079 27591
rect 10149 27557 10183 27591
rect 17233 27557 17267 27591
rect 18061 27557 18095 27591
rect 19349 27557 19383 27591
rect 23857 27557 23891 27591
rect 24961 27557 24995 27591
rect 31401 27557 31435 27591
rect 32597 27557 32631 27591
rect 34897 27557 34931 27591
rect 9229 27489 9263 27523
rect 9321 27489 9355 27523
rect 23489 27489 23523 27523
rect 32229 27489 32263 27523
rect 36093 27489 36127 27523
rect 37841 27489 37875 27523
rect 46305 27489 46339 27523
rect 48145 27489 48179 27523
rect 7573 27421 7607 27455
rect 8401 27421 8435 27455
rect 9689 27421 9723 27455
rect 10333 27421 10367 27455
rect 11161 27421 11195 27455
rect 13093 27421 13127 27455
rect 17417 27421 17451 27455
rect 18061 27421 18095 27455
rect 19257 27421 19291 27455
rect 22753 27421 22787 27455
rect 22937 27421 22971 27455
rect 23673 27421 23707 27455
rect 24777 27421 24811 27455
rect 26249 27421 26283 27455
rect 32413 27421 32447 27455
rect 33609 27421 33643 27455
rect 34713 27421 34747 27455
rect 38301 27421 38335 27455
rect 10517 27353 10551 27387
rect 22845 27353 22879 27387
rect 23397 27353 23431 27387
rect 29929 27353 29963 27387
rect 32137 27353 32171 27387
rect 46489 27353 46523 27387
rect 8217 27285 8251 27319
rect 9413 27285 9447 27319
rect 9597 27285 9631 27319
rect 10425 27285 10459 27319
rect 10701 27285 10735 27319
rect 11345 27285 11379 27319
rect 26341 27285 26375 27319
rect 33793 27285 33827 27319
rect 38393 27285 38427 27319
rect 13277 27081 13311 27115
rect 27905 27081 27939 27115
rect 29561 27081 29595 27115
rect 8401 27013 8435 27047
rect 9229 27013 9263 27047
rect 17233 27013 17267 27047
rect 17969 27013 18003 27047
rect 30205 27013 30239 27047
rect 30389 27013 30423 27047
rect 32505 27013 32539 27047
rect 9413 26945 9447 26979
rect 9505 26945 9539 26979
rect 10333 26945 10367 26979
rect 11529 26945 11563 26979
rect 14933 26945 14967 26979
rect 17141 26945 17175 26979
rect 17785 26945 17819 26979
rect 20085 26945 20119 26979
rect 22569 26945 22603 26979
rect 23489 26945 23523 26979
rect 24133 26945 24167 26979
rect 24869 26945 24903 26979
rect 27169 26945 27203 26979
rect 27721 26945 27755 26979
rect 29653 26945 29687 26979
rect 34713 26945 34747 26979
rect 38393 26945 38427 26979
rect 38577 26945 38611 26979
rect 10057 26877 10091 26911
rect 11805 26877 11839 26911
rect 19625 26877 19659 26911
rect 22845 26877 22879 26911
rect 24961 26877 24995 26911
rect 29193 26877 29227 26911
rect 32229 26877 32263 26911
rect 33977 26877 34011 26911
rect 8033 26809 8067 26843
rect 8401 26741 8435 26775
rect 8585 26741 8619 26775
rect 9505 26741 9539 26775
rect 15025 26741 15059 26775
rect 20177 26741 20211 26775
rect 22385 26741 22419 26775
rect 22753 26741 22787 26775
rect 23581 26741 23615 26775
rect 24317 26741 24351 26775
rect 26985 26741 27019 26775
rect 29377 26741 29411 26775
rect 34805 26741 34839 26775
rect 38761 26741 38795 26775
rect 12265 26537 12299 26571
rect 17141 26537 17175 26571
rect 18429 26537 18463 26571
rect 23305 26537 23339 26571
rect 33793 26537 33827 26571
rect 11253 26469 11287 26503
rect 12817 26469 12851 26503
rect 35081 26469 35115 26503
rect 9321 26401 9355 26435
rect 10885 26401 10919 26435
rect 13001 26401 13035 26435
rect 15025 26401 15059 26435
rect 16497 26401 16531 26435
rect 19257 26401 19291 26435
rect 19441 26401 19475 26435
rect 21557 26401 21591 26435
rect 25697 26401 25731 26435
rect 29561 26401 29595 26435
rect 31309 26401 31343 26435
rect 32413 26401 32447 26435
rect 37565 26401 37599 26435
rect 41153 26401 41187 26435
rect 7205 26333 7239 26367
rect 7389 26333 7423 26367
rect 8033 26333 8067 26367
rect 8309 26333 8343 26367
rect 9781 26333 9815 26367
rect 9965 26333 9999 26367
rect 12173 26333 12207 26367
rect 13093 26333 13127 26367
rect 13461 26333 13495 26367
rect 14841 26333 14875 26367
rect 17417 26333 17451 26367
rect 17509 26333 17543 26367
rect 17601 26333 17635 26367
rect 17785 26333 17819 26367
rect 18245 26333 18279 26367
rect 24869 26333 24903 26367
rect 32689 26333 32723 26367
rect 33701 26333 33735 26367
rect 34897 26333 34931 26367
rect 40877 26333 40911 26367
rect 47685 26333 47719 26367
rect 7297 26265 7331 26299
rect 8971 26265 9005 26299
rect 9137 26265 9171 26299
rect 13369 26265 13403 26299
rect 21097 26265 21131 26299
rect 21833 26265 21867 26299
rect 25053 26265 25087 26299
rect 25973 26265 26007 26299
rect 29837 26265 29871 26299
rect 37841 26265 37875 26299
rect 7849 26197 7883 26231
rect 8217 26197 8251 26231
rect 10149 26197 10183 26231
rect 11345 26197 11379 26231
rect 13277 26197 13311 26231
rect 27445 26197 27479 26231
rect 39313 26197 39347 26231
rect 11529 25993 11563 26027
rect 13093 25993 13127 26027
rect 14013 25993 14047 26027
rect 14289 25993 14323 26027
rect 15761 25993 15795 26027
rect 21833 25993 21867 26027
rect 26985 25993 27019 26027
rect 28549 25993 28583 26027
rect 29745 25993 29779 26027
rect 30297 25993 30331 26027
rect 31585 25993 31619 26027
rect 37473 25993 37507 26027
rect 7573 25925 7607 25959
rect 13737 25925 13771 25959
rect 15393 25925 15427 25959
rect 16957 25925 16991 25959
rect 19625 25925 19659 25959
rect 22201 25925 22235 25959
rect 22293 25925 22327 25959
rect 25329 25925 25363 25959
rect 28181 25925 28215 25959
rect 29377 25925 29411 25959
rect 32505 25925 32539 25959
rect 33517 25925 33551 25959
rect 41061 25925 41095 25959
rect 6745 25857 6779 25891
rect 11713 25857 11747 25891
rect 12449 25857 12483 25891
rect 12909 25857 12943 25891
rect 13921 25857 13955 25891
rect 14105 25857 14139 25891
rect 14749 25857 14783 25891
rect 15669 25857 15703 25891
rect 15853 25857 15887 25891
rect 20637 25857 20671 25891
rect 21097 25857 21131 25891
rect 21281 25857 21315 25891
rect 22845 25857 22879 25891
rect 23397 25857 23431 25891
rect 24685 25857 24719 25891
rect 24869 25857 24903 25891
rect 24961 25857 24995 25891
rect 25054 25857 25088 25891
rect 25789 25857 25823 25891
rect 25973 25857 26007 25891
rect 27353 25857 27387 25891
rect 28365 25857 28399 25891
rect 29101 25857 29135 25891
rect 29249 25857 29283 25891
rect 29469 25857 29503 25891
rect 29607 25857 29641 25891
rect 30205 25857 30239 25891
rect 31217 25857 31251 25891
rect 37749 25857 37783 25891
rect 37841 25857 37875 25891
rect 37933 25857 37967 25891
rect 38117 25857 38151 25891
rect 38577 25857 38611 25891
rect 38761 25857 38795 25891
rect 40233 25857 40267 25891
rect 46489 25857 46523 25891
rect 6837 25789 6871 25823
rect 7297 25789 7331 25823
rect 16129 25789 16163 25823
rect 17785 25789 17819 25823
rect 17969 25789 18003 25823
rect 22477 25789 22511 25823
rect 23673 25789 23707 25823
rect 27445 25789 27479 25823
rect 27629 25789 27663 25823
rect 31309 25789 31343 25823
rect 32597 25789 32631 25823
rect 32781 25789 32815 25823
rect 34253 25789 34287 25823
rect 34529 25789 34563 25823
rect 16037 25721 16071 25755
rect 21097 25721 21131 25755
rect 38945 25721 38979 25755
rect 9045 25653 9079 25687
rect 12265 25653 12299 25687
rect 14841 25653 14875 25687
rect 17049 25653 17083 25687
rect 20453 25653 20487 25687
rect 26157 25653 26191 25687
rect 28089 25653 28123 25687
rect 32137 25653 32171 25687
rect 33609 25653 33643 25687
rect 36001 25653 36035 25687
rect 38577 25653 38611 25687
rect 46581 25653 46615 25687
rect 47777 25653 47811 25687
rect 9045 25449 9079 25483
rect 13553 25449 13587 25483
rect 21005 25449 21039 25483
rect 22201 25449 22235 25483
rect 25513 25449 25547 25483
rect 27169 25449 27203 25483
rect 35357 25449 35391 25483
rect 37013 25449 37047 25483
rect 19901 25381 19935 25415
rect 22937 25381 22971 25415
rect 24777 25381 24811 25415
rect 30205 25381 30239 25415
rect 31953 25381 31987 25415
rect 33241 25381 33275 25415
rect 12081 25313 12115 25347
rect 15853 25313 15887 25347
rect 17509 25313 17543 25347
rect 26709 25313 26743 25347
rect 32413 25313 32447 25347
rect 32505 25313 32539 25347
rect 33425 25313 33459 25347
rect 33977 25313 34011 25347
rect 38393 25313 38427 25347
rect 40785 25313 40819 25347
rect 46489 25313 46523 25347
rect 48145 25313 48179 25347
rect 1409 25245 1443 25279
rect 7573 25245 7607 25279
rect 8953 25245 8987 25279
rect 9781 25245 9815 25279
rect 11805 25245 11839 25279
rect 14289 25245 14323 25279
rect 14565 25245 14599 25279
rect 15669 25245 15703 25279
rect 18521 25245 18555 25279
rect 20913 25245 20947 25279
rect 22845 25245 22879 25279
rect 23029 25245 23063 25279
rect 23121 25245 23155 25279
rect 23305 25245 23339 25279
rect 24623 25245 24657 25279
rect 24869 25245 24903 25279
rect 26801 25245 26835 25279
rect 30021 25245 30055 25279
rect 32321 25245 32355 25279
rect 33149 25245 33183 25279
rect 33885 25245 33919 25279
rect 34069 25245 34103 25279
rect 34713 25245 34747 25279
rect 34806 25245 34840 25279
rect 35081 25245 35115 25279
rect 35219 25245 35253 25279
rect 36737 25245 36771 25279
rect 37013 25245 37047 25279
rect 38117 25245 38151 25279
rect 40233 25245 40267 25279
rect 46305 25245 46339 25279
rect 1685 25177 1719 25211
rect 18337 25177 18371 25211
rect 18705 25177 18739 25211
rect 19717 25177 19751 25211
rect 21833 25177 21867 25211
rect 22017 25177 22051 25211
rect 24409 25177 24443 25211
rect 25421 25177 25455 25211
rect 33425 25177 33459 25211
rect 34989 25177 35023 25211
rect 36921 25177 36955 25211
rect 7757 25109 7791 25143
rect 9597 25109 9631 25143
rect 14105 25109 14139 25143
rect 14473 25109 14507 25143
rect 22661 25109 22695 25143
rect 13093 24905 13127 24939
rect 17233 24905 17267 24939
rect 24409 24905 24443 24939
rect 26065 24905 26099 24939
rect 33517 24905 33551 24939
rect 7573 24769 7607 24803
rect 10333 24769 10367 24803
rect 11529 24769 11563 24803
rect 12909 24769 12943 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 13829 24769 13863 24803
rect 15761 24769 15795 24803
rect 16037 24769 16071 24803
rect 17141 24769 17175 24803
rect 17785 24769 17819 24803
rect 21005 24769 21039 24803
rect 22569 24769 22603 24803
rect 22661 24769 22695 24803
rect 23489 24769 23523 24803
rect 23673 24769 23707 24803
rect 23765 24769 23799 24803
rect 24317 24769 24351 24803
rect 25973 24769 26007 24803
rect 26157 24769 26191 24803
rect 26433 24769 26467 24803
rect 27077 24769 27111 24803
rect 28641 24769 28675 24803
rect 29377 24769 29411 24803
rect 29561 24769 29595 24803
rect 30389 24769 30423 24803
rect 30573 24769 30607 24803
rect 32137 24769 32171 24803
rect 32413 24769 32447 24803
rect 33149 24769 33183 24803
rect 33333 24769 33367 24803
rect 37289 24769 37323 24803
rect 46489 24769 46523 24803
rect 47593 24769 47627 24803
rect 7849 24701 7883 24735
rect 12725 24701 12759 24735
rect 22385 24701 22419 24735
rect 22477 24701 22511 24735
rect 25697 24701 25731 24735
rect 27261 24701 27295 24735
rect 29837 24701 29871 24735
rect 32229 24701 32263 24735
rect 37565 24701 37599 24735
rect 46213 24701 46247 24735
rect 13645 24633 13679 24667
rect 23305 24633 23339 24667
rect 9321 24565 9355 24599
rect 10425 24565 10459 24599
rect 11621 24565 11655 24599
rect 15577 24565 15611 24599
rect 15945 24565 15979 24599
rect 17969 24565 18003 24599
rect 21097 24565 21131 24599
rect 22201 24565 22235 24599
rect 26341 24565 26375 24599
rect 28825 24565 28859 24599
rect 30481 24565 30515 24599
rect 32321 24565 32355 24599
rect 32597 24565 32631 24599
rect 33149 24565 33183 24599
rect 37381 24565 37415 24599
rect 37473 24565 37507 24599
rect 47685 24565 47719 24599
rect 13001 24361 13035 24395
rect 21833 24361 21867 24395
rect 22109 24361 22143 24395
rect 26249 24361 26283 24395
rect 28825 24361 28859 24395
rect 31309 24361 31343 24395
rect 31769 24361 31803 24395
rect 36921 24361 36955 24395
rect 37841 24361 37875 24395
rect 9045 24293 9079 24327
rect 12357 24293 12391 24327
rect 17509 24293 17543 24327
rect 26157 24293 26191 24327
rect 26893 24293 26927 24327
rect 29009 24293 29043 24327
rect 29699 24293 29733 24327
rect 29837 24293 29871 24327
rect 30481 24293 30515 24327
rect 37105 24293 37139 24327
rect 20085 24225 20119 24259
rect 23121 24225 23155 24259
rect 31493 24225 31527 24259
rect 33057 24225 33091 24259
rect 36829 24225 36863 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 8953 24157 8987 24191
rect 9965 24157 9999 24191
rect 12265 24157 12299 24191
rect 12909 24157 12943 24191
rect 16681 24157 16715 24191
rect 17417 24157 17451 24191
rect 19625 24157 19659 24191
rect 22845 24157 22879 24191
rect 25973 24157 26007 24191
rect 26065 24157 26099 24191
rect 26433 24157 26467 24191
rect 26893 24157 26927 24191
rect 27077 24157 27111 24191
rect 29561 24157 29595 24191
rect 30021 24157 30055 24191
rect 30757 24157 30791 24191
rect 31309 24157 31343 24191
rect 31585 24157 31619 24191
rect 32229 24157 32263 24191
rect 32413 24157 32447 24191
rect 32505 24157 32539 24191
rect 32965 24157 32999 24191
rect 33149 24157 33183 24191
rect 36185 24157 36219 24191
rect 36961 24157 36995 24191
rect 37662 24157 37696 24191
rect 37841 24157 37875 24191
rect 10241 24089 10275 24123
rect 20361 24089 20395 24123
rect 28641 24089 28675 24123
rect 28857 24089 28891 24123
rect 30481 24089 30515 24123
rect 35909 24089 35943 24123
rect 36093 24089 36127 24123
rect 36645 24089 36679 24123
rect 11713 24021 11747 24055
rect 16865 24021 16899 24055
rect 19717 24021 19751 24055
rect 22477 24021 22511 24055
rect 22937 24021 22971 24055
rect 25697 24021 25731 24055
rect 29929 24021 29963 24055
rect 30665 24021 30699 24055
rect 32321 24021 32355 24055
rect 36185 24021 36219 24055
rect 38025 24021 38059 24055
rect 1961 23817 1995 23851
rect 10149 23817 10183 23851
rect 26341 23817 26375 23851
rect 31309 23817 31343 23851
rect 34713 23817 34747 23851
rect 38485 23817 38519 23851
rect 27077 23749 27111 23783
rect 29837 23749 29871 23783
rect 1869 23681 1903 23715
rect 9781 23681 9815 23715
rect 11529 23681 11563 23715
rect 12449 23681 12483 23715
rect 16681 23681 16715 23715
rect 17693 23681 17727 23715
rect 18429 23681 18463 23715
rect 22477 23681 22511 23715
rect 24041 23681 24075 23715
rect 26249 23681 26283 23715
rect 26433 23681 26467 23715
rect 26985 23681 27019 23715
rect 29561 23681 29595 23715
rect 32137 23681 32171 23715
rect 32321 23681 32355 23715
rect 32413 23681 32447 23715
rect 32689 23681 32723 23715
rect 34713 23681 34747 23715
rect 35449 23681 35483 23715
rect 36369 23681 36403 23715
rect 36553 23681 36587 23715
rect 36737 23681 36771 23715
rect 37565 23681 37599 23715
rect 37657 23681 37691 23715
rect 37749 23681 37783 23715
rect 37933 23681 37967 23715
rect 38393 23681 38427 23715
rect 38577 23681 38611 23715
rect 45201 23681 45235 23715
rect 47593 23681 47627 23715
rect 9873 23613 9907 23647
rect 12541 23613 12575 23647
rect 13461 23613 13495 23647
rect 13737 23613 13771 23647
rect 18705 23613 18739 23647
rect 24133 23613 24167 23647
rect 24409 23613 24443 23647
rect 32505 23613 32539 23647
rect 35541 23613 35575 23647
rect 37289 23613 37323 23647
rect 45385 23613 45419 23647
rect 46857 23613 46891 23647
rect 11713 23477 11747 23511
rect 15209 23477 15243 23511
rect 16773 23477 16807 23511
rect 17877 23477 17911 23511
rect 20177 23477 20211 23511
rect 22293 23477 22327 23511
rect 32873 23477 32907 23511
rect 35725 23477 35759 23511
rect 47685 23477 47719 23511
rect 14657 23273 14691 23307
rect 19349 23273 19383 23307
rect 23765 23273 23799 23307
rect 27077 23273 27111 23307
rect 27537 23273 27571 23307
rect 27997 23273 28031 23307
rect 30297 23273 30331 23307
rect 31217 23273 31251 23307
rect 38485 23273 38519 23307
rect 14381 23137 14415 23171
rect 16773 23137 16807 23171
rect 17049 23137 17083 23171
rect 22017 23137 22051 23171
rect 25329 23137 25363 23171
rect 25605 23137 25639 23171
rect 35265 23137 35299 23171
rect 46489 23137 46523 23171
rect 10425 23069 10459 23103
rect 11529 23069 11563 23103
rect 12357 23069 12391 23103
rect 13277 23069 13311 23103
rect 14289 23069 14323 23103
rect 15117 23069 15151 23103
rect 16589 23069 16623 23103
rect 19257 23069 19291 23103
rect 20637 23069 20671 23103
rect 27721 23069 27755 23103
rect 27813 23069 27847 23103
rect 30297 23069 30331 23103
rect 30481 23069 30515 23103
rect 31125 23069 31159 23103
rect 32965 23069 32999 23103
rect 36737 23069 36771 23103
rect 41429 23069 41463 23103
rect 42165 23069 42199 23103
rect 46305 23069 46339 23103
rect 10793 23001 10827 23035
rect 22293 23001 22327 23035
rect 27537 23001 27571 23035
rect 35173 23001 35207 23035
rect 37013 23001 37047 23035
rect 42441 23001 42475 23035
rect 48145 23001 48179 23035
rect 11713 22933 11747 22967
rect 12449 22933 12483 22967
rect 13461 22933 13495 22967
rect 15301 22933 15335 22967
rect 20453 22933 20487 22967
rect 33057 22933 33091 22967
rect 34713 22933 34747 22967
rect 35081 22933 35115 22967
rect 41613 22933 41647 22967
rect 13277 22729 13311 22763
rect 14289 22729 14323 22763
rect 18429 22729 18463 22763
rect 47685 22729 47719 22763
rect 16957 22661 16991 22695
rect 18981 22661 19015 22695
rect 23397 22661 23431 22695
rect 26341 22661 26375 22695
rect 32413 22661 32447 22695
rect 35173 22661 35207 22695
rect 37381 22661 37415 22695
rect 41521 22661 41555 22695
rect 45385 22661 45419 22695
rect 8033 22593 8067 22627
rect 8677 22593 8711 22627
rect 11529 22593 11563 22627
rect 14197 22593 14231 22627
rect 15853 22593 15887 22627
rect 18889 22593 18923 22627
rect 19717 22593 19751 22627
rect 20545 22593 20579 22627
rect 23305 22593 23339 22627
rect 26249 22593 26283 22627
rect 26985 22593 27019 22627
rect 27077 22593 27111 22627
rect 35081 22593 35115 22627
rect 36093 22593 36127 22627
rect 37289 22593 37323 22627
rect 47593 22593 47627 22627
rect 8861 22525 8895 22559
rect 9137 22525 9171 22559
rect 11805 22525 11839 22559
rect 16681 22525 16715 22559
rect 27261 22525 27295 22559
rect 32137 22525 32171 22559
rect 33885 22525 33919 22559
rect 35357 22525 35391 22559
rect 42441 22525 42475 22559
rect 42625 22525 42659 22559
rect 44005 22525 44039 22559
rect 45201 22525 45235 22559
rect 45661 22525 45695 22559
rect 16037 22457 16071 22491
rect 26985 22457 27019 22491
rect 34713 22457 34747 22491
rect 8125 22389 8159 22423
rect 19993 22389 20027 22423
rect 20729 22389 20763 22423
rect 35909 22389 35943 22423
rect 41613 22389 41647 22423
rect 8309 22185 8343 22219
rect 14841 22185 14875 22219
rect 20802 22185 20836 22219
rect 41429 22185 41463 22219
rect 47961 22185 47995 22219
rect 12633 22117 12667 22151
rect 17049 22117 17083 22151
rect 23121 22117 23155 22151
rect 27997 22117 28031 22151
rect 32781 22117 32815 22151
rect 8953 22049 8987 22083
rect 9137 22049 9171 22083
rect 9413 22049 9447 22083
rect 16129 22049 16163 22083
rect 20545 22049 20579 22083
rect 34713 22049 34747 22083
rect 34989 22049 35023 22083
rect 36461 22049 36495 22083
rect 42717 22049 42751 22083
rect 46673 22049 46707 22083
rect 8217 21981 8251 22015
rect 11345 21981 11379 22015
rect 12357 21981 12391 22015
rect 15853 21981 15887 22015
rect 17785 21981 17819 22015
rect 19901 21981 19935 22015
rect 20085 21981 20119 22015
rect 23029 21981 23063 22015
rect 26157 21981 26191 22015
rect 26341 21981 26375 22015
rect 26801 21981 26835 22015
rect 27721 21981 27755 22015
rect 27813 21981 27847 22015
rect 28457 21981 28491 22015
rect 29837 21981 29871 22015
rect 30021 21981 30055 22015
rect 30113 21981 30147 22015
rect 32597 21981 32631 22015
rect 33425 21981 33459 22015
rect 38853 21981 38887 22015
rect 41337 21981 41371 22015
rect 42165 21981 42199 22015
rect 45477 21981 45511 22015
rect 14657 21913 14691 21947
rect 16681 21913 16715 21947
rect 18337 21913 18371 21947
rect 22569 21913 22603 21947
rect 26985 21913 27019 21947
rect 29653 21913 29687 21947
rect 45661 21913 45695 21947
rect 11437 21845 11471 21879
rect 12817 21845 12851 21879
rect 14857 21845 14891 21879
rect 15025 21845 15059 21879
rect 17141 21845 17175 21879
rect 20085 21845 20119 21879
rect 26341 21845 26375 21879
rect 27169 21845 27203 21879
rect 28549 21845 28583 21879
rect 33517 21845 33551 21879
rect 38945 21845 38979 21879
rect 11805 21641 11839 21675
rect 12633 21641 12667 21675
rect 13001 21641 13035 21675
rect 16773 21641 16807 21675
rect 17417 21641 17451 21675
rect 20821 21641 20855 21675
rect 26341 21641 26375 21675
rect 35633 21641 35667 21675
rect 44925 21641 44959 21675
rect 45661 21641 45695 21675
rect 15577 21573 15611 21607
rect 18429 21573 18463 21607
rect 18629 21573 18663 21607
rect 19809 21573 19843 21607
rect 30113 21573 30147 21607
rect 32229 21573 32263 21607
rect 38945 21573 38979 21607
rect 8861 21505 8895 21539
rect 11989 21505 12023 21539
rect 12817 21505 12851 21539
rect 13737 21505 13771 21539
rect 16957 21505 16991 21539
rect 17693 21505 17727 21539
rect 17877 21505 17911 21539
rect 19625 21505 19659 21539
rect 20453 21505 20487 21539
rect 20637 21505 20671 21539
rect 22385 21505 22419 21539
rect 22569 21505 22603 21539
rect 23029 21505 23063 21539
rect 23673 21505 23707 21539
rect 25329 21505 25363 21539
rect 26433 21505 26467 21539
rect 29837 21505 29871 21539
rect 32137 21505 32171 21539
rect 35541 21505 35575 21539
rect 42625 21505 42659 21539
rect 45109 21505 45143 21539
rect 45569 21505 45603 21539
rect 46213 21505 46247 21539
rect 47593 21505 47627 21539
rect 9045 21437 9079 21471
rect 9321 21437 9355 21471
rect 12909 21437 12943 21471
rect 13185 21437 13219 21471
rect 13277 21437 13311 21471
rect 13921 21437 13955 21471
rect 17601 21437 17635 21471
rect 17785 21437 17819 21471
rect 19993 21437 20027 21471
rect 25973 21437 26007 21471
rect 27537 21437 27571 21471
rect 27813 21437 27847 21471
rect 38761 21437 38795 21471
rect 39221 21437 39255 21471
rect 42809 21437 42843 21471
rect 46489 21437 46523 21471
rect 23121 21369 23155 21403
rect 18613 21301 18647 21335
rect 18797 21301 18831 21335
rect 22385 21301 22419 21335
rect 23765 21301 23799 21335
rect 25421 21301 25455 21335
rect 26157 21301 26191 21335
rect 29285 21301 29319 21335
rect 31585 21301 31619 21335
rect 47685 21301 47719 21335
rect 9137 21097 9171 21131
rect 12725 21097 12759 21131
rect 14289 21097 14323 21131
rect 14473 21097 14507 21131
rect 15025 21097 15059 21131
rect 17233 21097 17267 21131
rect 21925 21097 21959 21131
rect 28273 21097 28307 21131
rect 20545 20961 20579 20995
rect 24869 20961 24903 20995
rect 30389 20961 30423 20995
rect 42073 20961 42107 20995
rect 46489 20961 46523 20995
rect 48145 20961 48179 20995
rect 9045 20893 9079 20927
rect 9689 20893 9723 20927
rect 10333 20893 10367 20927
rect 10425 20893 10459 20927
rect 10977 20893 11011 20927
rect 14933 20893 14967 20927
rect 15577 20893 15611 20927
rect 17417 20893 17451 20927
rect 17601 20893 17635 20927
rect 17693 20893 17727 20927
rect 18153 20893 18187 20927
rect 19901 20893 19935 20927
rect 20821 20893 20855 20927
rect 22109 20893 22143 20927
rect 22201 20893 22235 20927
rect 22661 20893 22695 20927
rect 27629 20893 27663 20927
rect 27722 20893 27756 20927
rect 27905 20893 27939 20927
rect 28094 20893 28128 20927
rect 30481 20893 30515 20927
rect 41889 20893 41923 20927
rect 45845 20893 45879 20927
rect 46305 20893 46339 20927
rect 11253 20825 11287 20859
rect 14105 20825 14139 20859
rect 19717 20825 19751 20859
rect 21925 20825 21959 20859
rect 25145 20825 25179 20859
rect 27997 20825 28031 20859
rect 9781 20757 9815 20791
rect 14305 20757 14339 20791
rect 15669 20757 15703 20791
rect 18245 20757 18279 20791
rect 22845 20757 22879 20791
rect 26617 20757 26651 20791
rect 30849 20757 30883 20791
rect 11713 20553 11747 20587
rect 20821 20553 20855 20587
rect 25513 20553 25547 20587
rect 27537 20553 27571 20587
rect 29469 20553 29503 20587
rect 45569 20553 45603 20587
rect 8217 20485 8251 20519
rect 8953 20485 8987 20519
rect 20913 20485 20947 20519
rect 22753 20485 22787 20519
rect 24501 20485 24535 20519
rect 27353 20485 27387 20519
rect 29101 20485 29135 20519
rect 42901 20485 42935 20519
rect 8125 20417 8159 20451
rect 8769 20417 8803 20451
rect 11621 20417 11655 20451
rect 12449 20417 12483 20451
rect 12633 20417 12667 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 15945 20417 15979 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17601 20417 17635 20451
rect 18337 20417 18371 20451
rect 18521 20417 18555 20451
rect 19717 20417 19751 20451
rect 20729 20417 20763 20451
rect 22477 20417 22511 20451
rect 25697 20417 25731 20451
rect 25789 20417 25823 20451
rect 25973 20417 26007 20451
rect 26065 20417 26099 20451
rect 27169 20417 27203 20451
rect 28917 20417 28951 20451
rect 29193 20417 29227 20451
rect 29285 20417 29319 20451
rect 45477 20417 45511 20451
rect 46029 20417 46063 20451
rect 47593 20417 47627 20451
rect 9229 20349 9263 20383
rect 12542 20349 12576 20383
rect 12725 20349 12759 20383
rect 18245 20349 18279 20383
rect 18429 20349 18463 20383
rect 19993 20349 20027 20383
rect 20453 20349 20487 20383
rect 21189 20349 21223 20383
rect 46305 20349 46339 20383
rect 17509 20281 17543 20315
rect 12265 20213 12299 20247
rect 13369 20213 13403 20247
rect 16037 20213 16071 20247
rect 17049 20213 17083 20247
rect 18061 20213 18095 20247
rect 19533 20213 19567 20247
rect 19901 20213 19935 20247
rect 21097 20213 21131 20247
rect 43177 20213 43211 20247
rect 47685 20213 47719 20247
rect 11897 20009 11931 20043
rect 20913 20009 20947 20043
rect 21097 20009 21131 20043
rect 22017 20009 22051 20043
rect 22201 20009 22235 20043
rect 24869 20009 24903 20043
rect 25697 20009 25731 20043
rect 28181 20009 28215 20043
rect 9597 19873 9631 19907
rect 9781 19873 9815 19907
rect 12357 19873 12391 19907
rect 12817 19873 12851 19907
rect 14197 19873 14231 19907
rect 15301 19873 15335 19907
rect 17693 19873 17727 19907
rect 24501 19873 24535 19907
rect 25329 19873 25363 19907
rect 27813 19873 27847 19907
rect 30205 19873 30239 19907
rect 45845 19873 45879 19907
rect 46489 19873 46523 19907
rect 46949 19873 46983 19907
rect 2053 19805 2087 19839
rect 12081 19805 12115 19839
rect 12265 19805 12299 19839
rect 13001 19805 13035 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 15117 19805 15151 19839
rect 18245 19805 18279 19839
rect 20269 19805 20303 19839
rect 24685 19805 24719 19839
rect 25513 19805 25547 19839
rect 27997 19805 28031 19839
rect 30021 19805 30055 19839
rect 44281 19805 44315 19839
rect 44465 19805 44499 19839
rect 45477 19805 45511 19839
rect 45661 19805 45695 19839
rect 46305 19805 46339 19839
rect 22063 19771 22097 19805
rect 11437 19737 11471 19771
rect 16957 19737 16991 19771
rect 17877 19737 17911 19771
rect 17969 19737 18003 19771
rect 19717 19737 19751 19771
rect 19901 19737 19935 19771
rect 19993 19737 20027 19771
rect 20729 19737 20763 19771
rect 21833 19737 21867 19771
rect 13185 19669 13219 19703
rect 18061 19669 18095 19703
rect 20085 19669 20119 19703
rect 20929 19669 20963 19703
rect 44373 19669 44407 19703
rect 12449 19465 12483 19499
rect 18429 19465 18463 19499
rect 18981 19465 19015 19499
rect 45293 19465 45327 19499
rect 9413 19397 9447 19431
rect 12081 19397 12115 19431
rect 16957 19397 16991 19431
rect 1777 19329 1811 19363
rect 9321 19329 9355 19363
rect 12265 19329 12299 19363
rect 13185 19329 13219 19363
rect 15577 19329 15611 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 22477 19329 22511 19363
rect 24317 19329 24351 19363
rect 27537 19329 27571 19363
rect 42441 19329 42475 19363
rect 45201 19329 45235 19363
rect 45385 19329 45419 19363
rect 45937 19329 45971 19363
rect 46121 19329 46155 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 13461 19261 13495 19295
rect 14933 19261 14967 19295
rect 15853 19261 15887 19295
rect 16681 19261 16715 19295
rect 22569 19261 22603 19295
rect 46857 19261 46891 19295
rect 22845 19125 22879 19159
rect 24501 19125 24535 19159
rect 27629 19125 27663 19159
rect 42533 19125 42567 19159
rect 47777 19125 47811 19159
rect 2237 18921 2271 18955
rect 12633 18921 12667 18955
rect 14105 18921 14139 18955
rect 14933 18921 14967 18955
rect 18337 18921 18371 18955
rect 18521 18921 18555 18955
rect 19993 18921 20027 18955
rect 20729 18921 20763 18955
rect 20913 18921 20947 18955
rect 45661 18921 45695 18955
rect 17509 18853 17543 18887
rect 28457 18853 28491 18887
rect 9229 18785 9263 18819
rect 9413 18785 9447 18819
rect 9689 18785 9723 18819
rect 12265 18785 12299 18819
rect 17693 18785 17727 18819
rect 26157 18785 26191 18819
rect 27537 18785 27571 18819
rect 41429 18785 41463 18819
rect 41705 18785 41739 18819
rect 46305 18785 46339 18819
rect 48145 18785 48179 18819
rect 2145 18717 2179 18751
rect 11713 18717 11747 18751
rect 12357 18717 12391 18751
rect 13369 18717 13403 18751
rect 14289 18717 14323 18751
rect 14841 18717 14875 18751
rect 16773 18717 16807 18751
rect 22385 18717 22419 18751
rect 24409 18717 24443 18751
rect 25973 18717 26007 18751
rect 28273 18717 28307 18751
rect 41245 18717 41279 18751
rect 45569 18717 45603 18751
rect 45753 18717 45787 18751
rect 17233 18649 17267 18683
rect 18153 18649 18187 18683
rect 19717 18649 19751 18683
rect 20545 18649 20579 18683
rect 20745 18649 20779 18683
rect 29653 18649 29687 18683
rect 29745 18649 29779 18683
rect 30665 18649 30699 18683
rect 46489 18649 46523 18683
rect 11529 18581 11563 18615
rect 13369 18581 13403 18615
rect 16589 18581 16623 18615
rect 18363 18581 18397 18615
rect 22569 18581 22603 18615
rect 24501 18581 24535 18615
rect 1593 18377 1627 18411
rect 25697 18377 25731 18411
rect 47685 18377 47719 18411
rect 12909 18309 12943 18343
rect 16957 18309 16991 18343
rect 23029 18309 23063 18343
rect 26249 18309 26283 18343
rect 27445 18309 27479 18343
rect 1409 18241 1443 18275
rect 15669 18241 15703 18275
rect 19349 18241 19383 18275
rect 19533 18241 19567 18275
rect 20177 18241 20211 18275
rect 21005 18241 21039 18275
rect 21833 18241 21867 18275
rect 22753 18241 22787 18275
rect 26065 18241 26099 18275
rect 46397 18241 46431 18275
rect 47593 18241 47627 18275
rect 12633 18173 12667 18207
rect 14381 18173 14415 18207
rect 15945 18173 15979 18207
rect 16681 18173 16715 18207
rect 20269 18173 20303 18207
rect 24777 18173 24811 18207
rect 27261 18173 27295 18207
rect 28181 18173 28215 18207
rect 18429 18037 18463 18071
rect 19349 18037 19383 18071
rect 20545 18037 20579 18071
rect 21005 18037 21039 18071
rect 21925 18037 21959 18071
rect 26433 18037 26467 18071
rect 46213 18037 46247 18071
rect 47041 18037 47075 18071
rect 14197 17833 14231 17867
rect 16957 17833 16991 17867
rect 19809 17833 19843 17867
rect 20545 17697 20579 17731
rect 20821 17697 20855 17731
rect 39957 17697 39991 17731
rect 40233 17697 40267 17731
rect 46489 17697 46523 17731
rect 14105 17629 14139 17663
rect 16865 17629 16899 17663
rect 18245 17629 18279 17663
rect 20085 17629 20119 17663
rect 25513 17629 25547 17663
rect 25697 17629 25731 17663
rect 25881 17629 25915 17663
rect 26433 17629 26467 17663
rect 27077 17629 27111 17663
rect 46305 17629 46339 17663
rect 48145 17629 48179 17663
rect 19809 17561 19843 17595
rect 40049 17561 40083 17595
rect 18429 17493 18463 17527
rect 19993 17493 20027 17527
rect 22293 17493 22327 17527
rect 21281 17289 21315 17323
rect 27353 17289 27387 17323
rect 19809 17221 19843 17255
rect 21925 17221 21959 17255
rect 23673 17221 23707 17255
rect 46765 17221 46799 17255
rect 17141 17153 17175 17187
rect 17693 17153 17727 17187
rect 21833 17153 21867 17187
rect 25421 17153 25455 17187
rect 25697 17153 25731 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 47593 17153 47627 17187
rect 19533 17085 19567 17119
rect 23581 17085 23615 17119
rect 24593 17085 24627 17119
rect 25789 17085 25823 17119
rect 46213 17085 46247 17119
rect 2053 16949 2087 16983
rect 16957 16949 16991 16983
rect 17785 16949 17819 16983
rect 25513 16949 25547 16983
rect 25881 16949 25915 16983
rect 47685 16949 47719 16983
rect 19901 16745 19935 16779
rect 1409 16609 1443 16643
rect 1961 16609 1995 16643
rect 16681 16609 16715 16643
rect 25513 16609 25547 16643
rect 27169 16609 27203 16643
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 14381 16541 14415 16575
rect 19901 16541 19935 16575
rect 23397 16541 23431 16575
rect 25973 16541 26007 16575
rect 26157 16541 26191 16575
rect 26801 16541 26835 16575
rect 26985 16541 27019 16575
rect 1593 16473 1627 16507
rect 14565 16473 14599 16507
rect 16221 16473 16255 16507
rect 16957 16473 16991 16507
rect 18705 16473 18739 16507
rect 25145 16473 25179 16507
rect 25329 16473 25363 16507
rect 46489 16473 46523 16507
rect 23489 16405 23523 16439
rect 26341 16405 26375 16439
rect 2145 16201 2179 16235
rect 15025 16201 15059 16235
rect 17509 16201 17543 16235
rect 26157 16201 26191 16235
rect 26249 16201 26283 16235
rect 23489 16133 23523 16167
rect 26433 16133 26467 16167
rect 27905 16133 27939 16167
rect 46397 16133 46431 16167
rect 47961 16133 47995 16167
rect 2053 16065 2087 16099
rect 14933 16065 14967 16099
rect 17141 16065 17175 16099
rect 19441 16065 19475 16099
rect 19625 16065 19659 16099
rect 20913 16065 20947 16099
rect 23305 16065 23339 16099
rect 26065 16065 26099 16099
rect 27077 16065 27111 16099
rect 27261 16065 27295 16099
rect 27813 16065 27847 16099
rect 27997 16065 28031 16099
rect 40049 16065 40083 16099
rect 43913 16065 43947 16099
rect 46765 16065 46799 16099
rect 47593 16065 47627 16099
rect 47777 16065 47811 16099
rect 17233 15997 17267 16031
rect 25145 15997 25179 16031
rect 25881 15997 25915 16031
rect 40233 15997 40267 16031
rect 41889 15997 41923 16031
rect 44097 15997 44131 16031
rect 45477 15997 45511 16031
rect 46857 15997 46891 16031
rect 27261 15929 27295 15963
rect 47041 15929 47075 15963
rect 19441 15861 19475 15895
rect 21005 15861 21039 15895
rect 19809 15657 19843 15691
rect 20453 15657 20487 15691
rect 25513 15657 25547 15691
rect 27813 15657 27847 15691
rect 40509 15657 40543 15691
rect 44005 15657 44039 15691
rect 45753 15657 45787 15691
rect 47961 15657 47995 15691
rect 19993 15589 20027 15623
rect 2053 15453 2087 15487
rect 15117 15453 15151 15487
rect 17141 15453 17175 15487
rect 17693 15453 17727 15487
rect 20637 15453 20671 15487
rect 20729 15453 20763 15487
rect 21189 15453 21223 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 22201 15453 22235 15487
rect 25421 15453 25455 15487
rect 25605 15453 25639 15487
rect 26525 15453 26559 15487
rect 27169 15453 27203 15487
rect 31217 15453 31251 15487
rect 40417 15453 40451 15487
rect 43913 15453 43947 15487
rect 45661 15453 45695 15487
rect 45845 15453 45879 15487
rect 46673 15453 46707 15487
rect 47041 15453 47075 15487
rect 47869 15453 47903 15487
rect 48053 15453 48087 15487
rect 19625 15385 19659 15419
rect 20453 15385 20487 15419
rect 47409 15385 47443 15419
rect 15209 15317 15243 15351
rect 17141 15317 17175 15351
rect 17785 15317 17819 15351
rect 19835 15317 19869 15351
rect 22017 15317 22051 15351
rect 31309 15317 31343 15351
rect 26157 15113 26191 15147
rect 27077 15113 27111 15147
rect 47685 15113 47719 15147
rect 19533 15045 19567 15079
rect 22109 15045 22143 15079
rect 1777 14977 1811 15011
rect 16681 14977 16715 15011
rect 21833 14977 21867 15011
rect 25973 14977 26007 15011
rect 26157 14977 26191 15011
rect 26985 14977 27019 15011
rect 46305 14977 46339 15011
rect 46489 14977 46523 15011
rect 47593 14977 47627 15011
rect 47777 14977 47811 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 16957 14909 16991 14943
rect 19257 14909 19291 14943
rect 43545 14909 43579 14943
rect 43729 14909 43763 14943
rect 45109 14909 45143 14943
rect 21005 14841 21039 14875
rect 18429 14773 18463 14807
rect 23581 14773 23615 14807
rect 46397 14773 46431 14807
rect 2237 14569 2271 14603
rect 17601 14569 17635 14603
rect 19625 14569 19659 14603
rect 19809 14569 19843 14603
rect 21189 14569 21223 14603
rect 21741 14569 21775 14603
rect 22937 14569 22971 14603
rect 43637 14569 43671 14603
rect 47409 14569 47443 14603
rect 17969 14501 18003 14535
rect 15209 14433 15243 14467
rect 15485 14433 15519 14467
rect 30389 14433 30423 14467
rect 30573 14433 30607 14467
rect 2145 14365 2179 14399
rect 15025 14365 15059 14399
rect 17785 14365 17819 14399
rect 18061 14365 18095 14399
rect 21005 14365 21039 14399
rect 21649 14365 21683 14399
rect 22845 14365 22879 14399
rect 43545 14365 43579 14399
rect 46305 14365 46339 14399
rect 46489 14365 46523 14399
rect 46581 14365 46615 14399
rect 47041 14365 47075 14399
rect 47225 14365 47259 14399
rect 19441 14297 19475 14331
rect 19657 14297 19691 14331
rect 20821 14297 20855 14331
rect 32229 14297 32263 14331
rect 46121 14229 46155 14263
rect 46673 14025 46707 14059
rect 19441 13957 19475 13991
rect 20913 13957 20947 13991
rect 19165 13889 19199 13923
rect 20821 13889 20855 13923
rect 21005 13889 21039 13923
rect 45661 13889 45695 13923
rect 46029 13889 46063 13923
rect 46121 13889 46155 13923
rect 46581 13889 46615 13923
rect 46765 13889 46799 13923
rect 47593 13889 47627 13923
rect 45845 13855 45879 13889
rect 47685 13821 47719 13855
rect 20177 13277 20211 13311
rect 20821 13277 20855 13311
rect 46121 13277 46155 13311
rect 46673 13277 46707 13311
rect 48145 13277 48179 13311
rect 47501 13209 47535 13243
rect 20269 13141 20303 13175
rect 20913 13141 20947 13175
rect 46673 12937 46707 12971
rect 19625 12869 19659 12903
rect 45017 12869 45051 12903
rect 1409 12801 1443 12835
rect 44925 12801 44959 12835
rect 45109 12801 45143 12835
rect 45753 12801 45787 12835
rect 45937 12801 45971 12835
rect 46397 12801 46431 12835
rect 46581 12801 46615 12835
rect 19441 12733 19475 12767
rect 21281 12733 21315 12767
rect 45569 12733 45603 12767
rect 1593 12597 1627 12631
rect 45753 12393 45787 12427
rect 19533 12257 19567 12291
rect 19717 12257 19751 12291
rect 46305 12257 46339 12291
rect 46489 12257 46523 12291
rect 48145 12257 48179 12291
rect 45661 12189 45695 12223
rect 45845 12189 45879 12223
rect 21373 12121 21407 12155
rect 46121 11781 46155 11815
rect 46029 11645 46063 11679
rect 46305 11645 46339 11679
rect 47777 11509 47811 11543
rect 46305 11169 46339 11203
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 47685 10761 47719 10795
rect 47593 10625 47627 10659
rect 47041 10421 47075 10455
rect 19257 10081 19291 10115
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 19441 9945 19475 9979
rect 21097 9945 21131 9979
rect 46489 9945 46523 9979
rect 19257 9605 19291 9639
rect 47685 9605 47719 9639
rect 19165 9537 19199 9571
rect 47041 9537 47075 9571
rect 47593 9537 47627 9571
rect 46857 9401 46891 9435
rect 47317 8925 47351 8959
rect 47593 8925 47627 8959
rect 47777 8517 47811 8551
rect 47961 8313 47995 8347
rect 46305 7905 46339 7939
rect 46489 7905 46523 7939
rect 47961 7905 47995 7939
rect 48145 7361 48179 7395
rect 47961 7157 47995 7191
rect 47133 6817 47167 6851
rect 48053 6817 48087 6851
rect 47225 6681 47259 6715
rect 46489 6273 46523 6307
rect 48145 6273 48179 6307
rect 46213 6205 46247 6239
rect 47961 6069 47995 6103
rect 46305 5729 46339 5763
rect 47869 5729 47903 5763
rect 46489 5593 46523 5627
rect 19625 5253 19659 5287
rect 31217 5253 31251 5287
rect 46029 5253 46063 5287
rect 46121 5253 46155 5287
rect 18245 5185 18279 5219
rect 18889 5185 18923 5219
rect 19533 5185 19567 5219
rect 20269 5185 20303 5219
rect 20913 5185 20947 5219
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 23121 5185 23155 5219
rect 45293 5185 45327 5219
rect 47869 5185 47903 5219
rect 29377 5117 29411 5151
rect 29561 5117 29595 5151
rect 46857 5117 46891 5151
rect 18981 5049 19015 5083
rect 48053 5049 48087 5083
rect 18337 4981 18371 5015
rect 20361 4981 20395 5015
rect 21005 4981 21039 5015
rect 21925 4981 21959 5015
rect 22569 4981 22603 5015
rect 23213 4981 23247 5015
rect 45385 4981 45419 5015
rect 18337 4777 18371 4811
rect 21281 4777 21315 4811
rect 21925 4777 21959 4811
rect 45753 4641 45787 4675
rect 45937 4641 45971 4675
rect 46949 4641 46983 4675
rect 18245 4573 18279 4607
rect 19257 4573 19291 4607
rect 19901 4573 19935 4607
rect 20545 4573 20579 4607
rect 20637 4573 20671 4607
rect 21189 4573 21223 4607
rect 21833 4573 21867 4607
rect 22477 4573 22511 4607
rect 23121 4573 23155 4607
rect 42533 4573 42567 4607
rect 44097 4573 44131 4607
rect 45293 4573 45327 4607
rect 19349 4437 19383 4471
rect 19993 4437 20027 4471
rect 22569 4437 22603 4471
rect 23213 4437 23247 4471
rect 43913 4437 43947 4471
rect 19349 4233 19383 4267
rect 19993 4233 20027 4267
rect 20637 4233 20671 4267
rect 21925 4233 21959 4267
rect 22569 4233 22603 4267
rect 39957 4233 39991 4267
rect 43085 4165 43119 4199
rect 2145 4097 2179 4131
rect 2789 4097 2823 4131
rect 6561 4097 6595 4131
rect 7205 4097 7239 4131
rect 7849 4097 7883 4131
rect 11897 4097 11931 4131
rect 17509 4097 17543 4131
rect 18153 4097 18187 4131
rect 19257 4097 19291 4131
rect 19901 4097 19935 4131
rect 20545 4097 20579 4131
rect 21833 4097 21867 4131
rect 22477 4097 22511 4131
rect 23121 4097 23155 4131
rect 23765 4097 23799 4131
rect 23857 4097 23891 4131
rect 24593 4097 24627 4131
rect 39221 4097 39255 4131
rect 39865 4097 39899 4131
rect 40969 4097 41003 4131
rect 42901 4097 42935 4131
rect 44741 4097 44775 4131
rect 45201 4097 45235 4131
rect 47869 4097 47903 4131
rect 41153 4029 41187 4063
rect 45385 4029 45419 4063
rect 45937 4029 45971 4063
rect 7941 3961 7975 3995
rect 17601 3961 17635 3995
rect 48053 3961 48087 3995
rect 2237 3893 2271 3927
rect 2881 3893 2915 3927
rect 6653 3893 6687 3927
rect 7297 3893 7331 3927
rect 9505 3893 9539 3927
rect 11989 3893 12023 3927
rect 18245 3893 18279 3927
rect 23213 3893 23247 3927
rect 24409 3893 24443 3927
rect 39313 3893 39347 3927
rect 41337 3893 41371 3927
rect 39221 3689 39255 3723
rect 6653 3553 6687 3587
rect 7205 3553 7239 3587
rect 11253 3553 11287 3587
rect 11529 3553 11563 3587
rect 17141 3553 17175 3587
rect 25513 3553 25547 3587
rect 26801 3553 26835 3587
rect 40049 3553 40083 3587
rect 41337 3553 41371 3587
rect 44465 3553 44499 3587
rect 1409 3485 1443 3519
rect 2329 3485 2363 3519
rect 2973 3485 3007 3519
rect 6009 3485 6043 3519
rect 6469 3485 6503 3519
rect 9137 3485 9171 3519
rect 9965 3485 9999 3519
rect 11069 3485 11103 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 15301 3485 15335 3519
rect 18061 3485 18095 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 20729 3485 20763 3519
rect 21557 3485 21591 3519
rect 22753 3485 22787 3519
rect 22845 3485 22879 3519
rect 23397 3485 23431 3519
rect 23489 3485 23523 3519
rect 24685 3485 24719 3519
rect 26525 3485 26559 3519
rect 32965 3485 32999 3519
rect 33057 3485 33091 3519
rect 33793 3485 33827 3519
rect 35909 3485 35943 3519
rect 38485 3485 38519 3519
rect 39129 3485 39163 3519
rect 40325 3485 40359 3519
rect 43637 3485 43671 3519
rect 45017 3485 45051 3519
rect 45661 3487 45695 3521
rect 46305 3485 46339 3519
rect 15485 3417 15519 3451
rect 22109 3417 22143 3451
rect 36093 3417 36127 3451
rect 37749 3417 37783 3451
rect 41521 3417 41555 3451
rect 43177 3417 43211 3451
rect 45753 3417 45787 3451
rect 46489 3417 46523 3451
rect 48145 3417 48179 3451
rect 1593 3349 1627 3383
rect 10057 3349 10091 3383
rect 14197 3349 14231 3383
rect 18153 3349 18187 3383
rect 19533 3349 19567 3383
rect 20821 3349 20855 3383
rect 22201 3349 22235 3383
rect 24777 3349 24811 3383
rect 38577 3349 38611 3383
rect 43729 3349 43763 3383
rect 45109 3349 45143 3383
rect 18429 3145 18463 3179
rect 36185 3145 36219 3179
rect 39129 3145 39163 3179
rect 1961 3077 1995 3111
rect 7297 3077 7331 3111
rect 9689 3077 9723 3111
rect 13921 3077 13955 3111
rect 24777 3077 24811 3111
rect 28273 3077 28307 3111
rect 33057 3077 33091 3111
rect 39773 3077 39807 3111
rect 42625 3077 42659 3111
rect 45385 3077 45419 3111
rect 47777 3077 47811 3111
rect 1777 3009 1811 3043
rect 6653 3009 6687 3043
rect 7113 3009 7147 3043
rect 9505 3009 9539 3043
rect 11713 3009 11747 3043
rect 13737 3009 13771 3043
rect 17509 3009 17543 3043
rect 18337 3009 18371 3043
rect 19349 3009 19383 3043
rect 21833 3009 21867 3043
rect 24593 3009 24627 3043
rect 28089 3009 28123 3043
rect 36369 3009 36403 3043
rect 38485 3009 38519 3043
rect 38669 3009 38703 3043
rect 39589 3009 39623 3043
rect 42441 3009 42475 3043
rect 45201 3009 45235 3043
rect 2237 2941 2271 2975
rect 7757 2941 7791 2975
rect 14197 2941 14231 2975
rect 17417 2941 17451 2975
rect 17877 2941 17911 2975
rect 19533 2941 19567 2975
rect 19993 2941 20027 2975
rect 22017 2941 22051 2975
rect 22569 2941 22603 2975
rect 25145 2941 25179 2975
rect 29929 2941 29963 2975
rect 32873 2941 32907 2975
rect 33517 2941 33551 2975
rect 40049 2941 40083 2975
rect 43177 2941 43211 2975
rect 47041 2941 47075 2975
rect 47869 2805 47903 2839
rect 18613 2601 18647 2635
rect 19349 2601 19383 2635
rect 23029 2601 23063 2635
rect 26157 2601 26191 2635
rect 35771 2601 35805 2635
rect 47869 2601 47903 2635
rect 17325 2533 17359 2567
rect 40509 2533 40543 2567
rect 43085 2533 43119 2567
rect 1409 2465 1443 2499
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 6561 2465 6595 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 9137 2465 9171 2499
rect 9689 2465 9723 2499
rect 15577 2465 15611 2499
rect 20729 2465 20763 2499
rect 24501 2465 24535 2499
rect 25513 2465 25547 2499
rect 28457 2465 28491 2499
rect 30021 2465 30055 2499
rect 38393 2465 38427 2499
rect 41337 2465 41371 2499
rect 43637 2465 43671 2499
rect 46213 2465 46247 2499
rect 4997 2397 5031 2431
rect 15301 2397 15335 2431
rect 18521 2397 18555 2431
rect 19257 2397 19291 2431
rect 20453 2397 20487 2431
rect 22201 2397 22235 2431
rect 23121 2397 23155 2431
rect 28181 2397 28215 2431
rect 29745 2397 29779 2431
rect 35541 2397 35575 2431
rect 41061 2397 41095 2431
rect 43913 2397 43947 2431
rect 45477 2397 45511 2431
rect 46489 2397 46523 2431
rect 1593 2329 1627 2363
rect 4169 2329 4203 2363
rect 9321 2329 9355 2363
rect 17141 2329 17175 2363
rect 24593 2329 24627 2363
rect 26065 2329 26099 2363
rect 27445 2329 27479 2363
rect 27629 2329 27663 2363
rect 38209 2329 38243 2363
rect 40325 2329 40359 2363
rect 42901 2329 42935 2363
rect 47777 2329 47811 2363
rect 4445 2261 4479 2295
rect 45661 2261 45695 2295
<< metal1 >>
rect 15286 47404 15292 47456
rect 15344 47444 15350 47456
rect 16482 47444 16488 47456
rect 15344 47416 16488 47444
rect 15344 47404 15350 47416
rect 16482 47404 16488 47416
rect 16540 47404 16546 47456
rect 40034 47404 40040 47456
rect 40092 47444 40098 47456
rect 41230 47444 41236 47456
rect 40092 47416 41236 47444
rect 40092 47404 40098 47416
rect 41230 47404 41236 47416
rect 41288 47404 41294 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 12437 47175 12495 47181
rect 12437 47141 12449 47175
rect 12483 47172 12495 47175
rect 12802 47172 12808 47184
rect 12483 47144 12808 47172
rect 12483 47141 12495 47144
rect 12437 47135 12495 47141
rect 12802 47132 12808 47144
rect 12860 47132 12866 47184
rect 19426 47172 19432 47184
rect 19387 47144 19432 47172
rect 19426 47132 19432 47144
rect 19484 47132 19490 47184
rect 29086 47132 29092 47184
rect 29144 47172 29150 47184
rect 29917 47175 29975 47181
rect 29917 47172 29929 47175
rect 29144 47144 29929 47172
rect 29144 47132 29150 47144
rect 29917 47141 29929 47144
rect 29963 47141 29975 47175
rect 29917 47135 29975 47141
rect 19978 47064 19984 47116
rect 20036 47104 20042 47116
rect 20073 47107 20131 47113
rect 20073 47104 20085 47107
rect 20036 47076 20085 47104
rect 20036 47064 20042 47076
rect 20073 47073 20085 47076
rect 20119 47073 20131 47107
rect 30742 47104 30748 47116
rect 30703 47076 30748 47104
rect 20073 47067 20131 47073
rect 30742 47064 30748 47076
rect 30800 47064 30806 47116
rect 43162 47104 43168 47116
rect 43123 47076 43168 47104
rect 43162 47064 43168 47076
rect 43220 47064 43226 47116
rect 47029 47107 47087 47113
rect 47029 47073 47041 47107
rect 47075 47104 47087 47107
rect 48314 47104 48320 47116
rect 47075 47076 48320 47104
rect 47075 47073 47087 47076
rect 47029 47067 47087 47073
rect 48314 47064 48320 47076
rect 48372 47064 48378 47116
rect 1946 47036 1952 47048
rect 1907 47008 1952 47036
rect 1946 46996 1952 47008
rect 2004 46996 2010 47048
rect 2590 46996 2596 47048
rect 2648 47036 2654 47048
rect 2685 47039 2743 47045
rect 2685 47036 2697 47039
rect 2648 47008 2697 47036
rect 2648 46996 2654 47008
rect 2685 47005 2697 47008
rect 2731 47005 2743 47039
rect 2685 46999 2743 47005
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3292 47008 3801 47036
rect 3292 46996 3298 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 4706 47036 4712 47048
rect 4667 47008 4712 47036
rect 3789 46999 3847 47005
rect 4706 46996 4712 47008
rect 4764 46996 4770 47048
rect 5810 46996 5816 47048
rect 5868 47036 5874 47048
rect 6825 47039 6883 47045
rect 6825 47036 6837 47039
rect 5868 47008 6837 47036
rect 5868 46996 5874 47008
rect 6825 47005 6837 47008
rect 6871 47005 6883 47039
rect 6825 46999 6883 47005
rect 7098 46996 7104 47048
rect 7156 47036 7162 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7156 47008 7757 47036
rect 7156 46996 7162 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 7745 46999 7803 47005
rect 9030 46996 9036 47048
rect 9088 47036 9094 47048
rect 9125 47039 9183 47045
rect 9125 47036 9137 47039
rect 9088 47008 9137 47036
rect 9088 46996 9094 47008
rect 9125 47005 9137 47008
rect 9171 47005 9183 47039
rect 11606 47036 11612 47048
rect 11567 47008 11612 47036
rect 9125 46999 9183 47005
rect 11606 46996 11612 47008
rect 11664 46996 11670 47048
rect 12250 47036 12256 47048
rect 12211 47008 12256 47036
rect 12250 46996 12256 47008
rect 12308 46996 12314 47048
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 13081 47039 13139 47045
rect 13081 47036 13093 47039
rect 12952 47008 13093 47036
rect 12952 46996 12958 47008
rect 13081 47005 13093 47008
rect 13127 47005 13139 47039
rect 13081 46999 13139 47005
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 14553 47039 14611 47045
rect 14553 47036 14565 47039
rect 13872 47008 14565 47036
rect 13872 46996 13878 47008
rect 14553 47005 14565 47008
rect 14599 47005 14611 47039
rect 14553 46999 14611 47005
rect 18690 46996 18696 47048
rect 18748 47036 18754 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18748 47008 19257 47036
rect 18748 46996 18754 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 19245 46999 19303 47005
rect 20349 47039 20407 47045
rect 20349 47005 20361 47039
rect 20395 47036 20407 47039
rect 22738 47036 22744 47048
rect 20395 47008 22744 47036
rect 20395 47005 20407 47008
rect 20349 46999 20407 47005
rect 22738 46996 22744 47008
rect 22796 46996 22802 47048
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 28350 46996 28356 47048
rect 28408 47036 28414 47048
rect 28629 47039 28687 47045
rect 28629 47036 28641 47039
rect 28408 47008 28641 47036
rect 28408 46996 28414 47008
rect 28629 47005 28641 47008
rect 28675 47005 28687 47039
rect 28629 46999 28687 47005
rect 29638 46996 29644 47048
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 31021 47039 31079 47045
rect 31021 47005 31033 47039
rect 31067 47036 31079 47039
rect 31110 47036 31116 47048
rect 31067 47008 31116 47036
rect 31067 47005 31079 47008
rect 31021 46999 31079 47005
rect 31110 46996 31116 47008
rect 31168 46996 31174 47048
rect 38102 46996 38108 47048
rect 38160 47036 38166 47048
rect 38289 47039 38347 47045
rect 38289 47036 38301 47039
rect 38160 47008 38301 47036
rect 38160 46996 38166 47008
rect 38289 47005 38301 47008
rect 38335 47005 38347 47039
rect 42610 47036 42616 47048
rect 42571 47008 42616 47036
rect 38289 46999 38347 47005
rect 42610 46996 42616 47008
rect 42668 46996 42674 47048
rect 44450 46996 44456 47048
rect 44508 47036 44514 47048
rect 45189 47039 45247 47045
rect 45189 47036 45201 47039
rect 44508 47008 45201 47036
rect 44508 46996 44514 47008
rect 45189 47005 45201 47008
rect 45235 47005 45247 47039
rect 45189 46999 45247 47005
rect 47670 46996 47676 47048
rect 47728 47036 47734 47048
rect 47765 47039 47823 47045
rect 47765 47036 47777 47039
rect 47728 47008 47777 47036
rect 47728 46996 47734 47008
rect 47765 47005 47777 47008
rect 47811 47005 47823 47039
rect 47765 46999 47823 47005
rect 4062 46968 4068 46980
rect 4023 46940 4068 46968
rect 4062 46928 4068 46940
rect 4120 46928 4126 46980
rect 4982 46968 4988 46980
rect 4943 46940 4988 46968
rect 4982 46928 4988 46940
rect 5040 46928 5046 46980
rect 7834 46928 7840 46980
rect 7892 46968 7898 46980
rect 7929 46971 7987 46977
rect 7929 46968 7941 46971
rect 7892 46940 7941 46968
rect 7892 46928 7898 46940
rect 7929 46937 7941 46940
rect 7975 46937 7987 46971
rect 7929 46931 7987 46937
rect 11698 46928 11704 46980
rect 11756 46968 11762 46980
rect 11793 46971 11851 46977
rect 11793 46968 11805 46971
rect 11756 46940 11805 46968
rect 11756 46928 11762 46940
rect 11793 46937 11805 46940
rect 11839 46937 11851 46971
rect 11793 46931 11851 46937
rect 13354 46928 13360 46980
rect 13412 46968 13418 46980
rect 13449 46971 13507 46977
rect 13449 46968 13461 46971
rect 13412 46940 13461 46968
rect 13412 46928 13418 46940
rect 13449 46937 13461 46940
rect 13495 46937 13507 46971
rect 13449 46931 13507 46937
rect 14642 46928 14648 46980
rect 14700 46968 14706 46980
rect 14737 46971 14795 46977
rect 14737 46968 14749 46971
rect 14700 46940 14749 46968
rect 14700 46928 14706 46940
rect 14737 46937 14749 46940
rect 14783 46937 14795 46971
rect 17129 46971 17187 46977
rect 17129 46968 17141 46971
rect 14737 46931 14795 46937
rect 16546 46940 17141 46968
rect 2130 46900 2136 46912
rect 2091 46872 2136 46900
rect 2130 46860 2136 46872
rect 2188 46860 2194 46912
rect 2866 46900 2872 46912
rect 2827 46872 2872 46900
rect 2866 46860 2872 46872
rect 2924 46860 2930 46912
rect 6914 46860 6920 46912
rect 6972 46900 6978 46912
rect 9306 46900 9312 46912
rect 6972 46872 7017 46900
rect 9267 46872 9312 46900
rect 6972 46860 6978 46872
rect 9306 46860 9312 46872
rect 9364 46860 9370 46912
rect 16114 46860 16120 46912
rect 16172 46900 16178 46912
rect 16546 46900 16574 46940
rect 17129 46937 17141 46940
rect 17175 46937 17187 46971
rect 17129 46931 17187 46937
rect 17313 46971 17371 46977
rect 17313 46937 17325 46971
rect 17359 46968 17371 46971
rect 17586 46968 17592 46980
rect 17359 46940 17592 46968
rect 17359 46937 17371 46940
rect 17313 46931 17371 46937
rect 17586 46928 17592 46940
rect 17644 46928 17650 46980
rect 40313 46971 40371 46977
rect 40313 46937 40325 46971
rect 40359 46937 40371 46971
rect 40313 46931 40371 46937
rect 16172 46872 16574 46900
rect 16172 46860 16178 46872
rect 28166 46860 28172 46912
rect 28224 46900 28230 46912
rect 28445 46903 28503 46909
rect 28445 46900 28457 46903
rect 28224 46872 28457 46900
rect 28224 46860 28230 46872
rect 28445 46869 28457 46872
rect 28491 46869 28503 46903
rect 28445 46863 28503 46869
rect 39298 46860 39304 46912
rect 39356 46900 39362 46912
rect 40328 46900 40356 46931
rect 40402 46928 40408 46980
rect 40460 46968 40466 46980
rect 40497 46971 40555 46977
rect 40497 46968 40509 46971
rect 40460 46940 40509 46968
rect 40460 46928 40466 46940
rect 40497 46937 40509 46940
rect 40543 46937 40555 46971
rect 40497 46931 40555 46937
rect 42797 46971 42855 46977
rect 42797 46937 42809 46971
rect 42843 46968 42855 46971
rect 43162 46968 43168 46980
rect 42843 46940 43168 46968
rect 42843 46937 42855 46940
rect 42797 46931 42855 46937
rect 43162 46928 43168 46940
rect 43220 46928 43226 46980
rect 45370 46968 45376 46980
rect 45331 46940 45376 46968
rect 45370 46928 45376 46940
rect 45428 46928 45434 46980
rect 47946 46900 47952 46912
rect 39356 46872 40356 46900
rect 47907 46872 47952 46900
rect 39356 46860 39362 46872
rect 47946 46860 47952 46872
rect 48004 46860 48010 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 6886 46668 26234 46696
rect 2866 46588 2872 46640
rect 2924 46628 2930 46640
rect 6886 46628 6914 46668
rect 24854 46628 24860 46640
rect 2924 46600 6914 46628
rect 24596 46600 24860 46628
rect 2924 46588 2930 46600
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 24596 46569 24624 46600
rect 24854 46588 24860 46600
rect 24912 46588 24918 46640
rect 26206 46628 26234 46668
rect 28353 46631 28411 46637
rect 28353 46628 28365 46631
rect 26206 46600 28365 46628
rect 28353 46597 28365 46600
rect 28399 46597 28411 46631
rect 28353 46591 28411 46597
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 28166 46560 28172 46572
rect 28127 46532 28172 46560
rect 24581 46523 24639 46529
rect 28166 46520 28172 46532
rect 28224 46520 28230 46572
rect 38102 46560 38108 46572
rect 38063 46532 38108 46560
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 47854 46560 47860 46572
rect 47815 46532 47860 46560
rect 47854 46520 47860 46532
rect 47912 46520 47918 46572
rect 3970 46492 3976 46504
rect 3931 46464 3976 46492
rect 3970 46452 3976 46464
rect 4028 46452 4034 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46492 4215 46495
rect 5074 46492 5080 46504
rect 4203 46464 5080 46492
rect 4203 46461 4215 46464
rect 4157 46455 4215 46461
rect 5074 46452 5080 46464
rect 5132 46452 5138 46504
rect 5169 46495 5227 46501
rect 5169 46461 5181 46495
rect 5215 46461 5227 46495
rect 5169 46455 5227 46461
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11517 46455 11575 46461
rect 11701 46495 11759 46501
rect 11701 46461 11713 46495
rect 11747 46492 11759 46495
rect 12158 46492 12164 46504
rect 11747 46464 12164 46492
rect 11747 46461 11759 46464
rect 11701 46455 11759 46461
rect 3878 46384 3884 46436
rect 3936 46424 3942 46436
rect 5184 46424 5212 46455
rect 12158 46452 12164 46464
rect 12216 46452 12222 46504
rect 12437 46495 12495 46501
rect 12437 46461 12449 46495
rect 12483 46461 12495 46495
rect 12437 46455 12495 46461
rect 3936 46396 5212 46424
rect 3936 46384 3942 46396
rect 1581 46359 1639 46365
rect 1581 46325 1593 46359
rect 1627 46356 1639 46359
rect 1670 46356 1676 46368
rect 1627 46328 1676 46356
rect 1627 46325 1639 46328
rect 1581 46319 1639 46325
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 10962 46316 10968 46368
rect 11020 46356 11026 46368
rect 12452 46356 12480 46455
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13817 46495 13875 46501
rect 13817 46492 13829 46495
rect 13596 46464 13829 46492
rect 13596 46452 13602 46464
rect 13817 46461 13829 46464
rect 13863 46461 13875 46495
rect 13817 46455 13875 46461
rect 14001 46495 14059 46501
rect 14001 46461 14013 46495
rect 14047 46492 14059 46495
rect 14182 46492 14188 46504
rect 14047 46464 14188 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 14182 46452 14188 46464
rect 14240 46452 14246 46504
rect 14274 46452 14280 46504
rect 14332 46492 14338 46504
rect 19242 46492 19248 46504
rect 14332 46464 14377 46492
rect 19203 46464 19248 46492
rect 14332 46452 14338 46464
rect 19242 46452 19248 46464
rect 19300 46452 19306 46504
rect 19429 46495 19487 46501
rect 19429 46461 19441 46495
rect 19475 46461 19487 46495
rect 20622 46492 20628 46504
rect 20583 46464 20628 46492
rect 19429 46455 19487 46461
rect 18598 46384 18604 46436
rect 18656 46424 18662 46436
rect 19444 46424 19472 46455
rect 20622 46452 20628 46464
rect 20680 46452 20686 46504
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 25130 46492 25136 46504
rect 25091 46464 25136 46492
rect 25130 46452 25136 46464
rect 25188 46452 25194 46504
rect 29362 46492 29368 46504
rect 29323 46464 29368 46492
rect 29362 46452 29368 46464
rect 29420 46452 29426 46504
rect 31573 46495 31631 46501
rect 31573 46461 31585 46495
rect 31619 46492 31631 46495
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 31619 46464 32137 46492
rect 31619 46461 31631 46464
rect 31573 46455 31631 46461
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32306 46492 32312 46504
rect 32267 46464 32312 46492
rect 32125 46455 32183 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 38286 46492 38292 46504
rect 38247 46464 38292 46492
rect 32585 46455 32643 46461
rect 18656 46396 19472 46424
rect 18656 46384 18662 46396
rect 32214 46384 32220 46436
rect 32272 46424 32278 46436
rect 32600 46424 32628 46455
rect 38286 46452 38292 46464
rect 38344 46452 38350 46504
rect 38654 46492 38660 46504
rect 38615 46464 38660 46492
rect 38654 46452 38660 46464
rect 38712 46452 38718 46504
rect 41877 46495 41935 46501
rect 41877 46461 41889 46495
rect 41923 46492 41935 46495
rect 42429 46495 42487 46501
rect 42429 46492 42441 46495
rect 41923 46464 42441 46492
rect 41923 46461 41935 46464
rect 41877 46455 41935 46461
rect 42429 46461 42441 46464
rect 42475 46461 42487 46495
rect 42610 46492 42616 46504
rect 42571 46464 42616 46492
rect 42429 46455 42487 46461
rect 42610 46452 42616 46464
rect 42668 46452 42674 46504
rect 42889 46495 42947 46501
rect 42889 46461 42901 46495
rect 42935 46461 42947 46495
rect 42889 46455 42947 46461
rect 45189 46495 45247 46501
rect 45189 46461 45201 46495
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46658 46492 46664 46504
rect 45419 46464 46664 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 32272 46396 32628 46424
rect 32272 46384 32278 46396
rect 42518 46384 42524 46436
rect 42576 46424 42582 46436
rect 42904 46424 42932 46455
rect 42576 46396 42932 46424
rect 45204 46424 45232 46455
rect 46658 46452 46664 46464
rect 46716 46452 46722 46504
rect 46842 46492 46848 46504
rect 46803 46464 46848 46492
rect 46842 46452 46848 46464
rect 46900 46452 46906 46504
rect 47762 46424 47768 46436
rect 45204 46396 47768 46424
rect 42576 46384 42582 46396
rect 47762 46384 47768 46396
rect 47820 46384 47826 46436
rect 11020 46328 12480 46356
rect 11020 46316 11026 46328
rect 20714 46316 20720 46368
rect 20772 46356 20778 46368
rect 22005 46359 22063 46365
rect 22005 46356 22017 46359
rect 20772 46328 22017 46356
rect 20772 46316 20778 46328
rect 22005 46325 22017 46328
rect 22051 46325 22063 46359
rect 41230 46356 41236 46368
rect 41191 46328 41236 46356
rect 22005 46319 22063 46325
rect 41230 46316 41236 46328
rect 41288 46316 41294 46368
rect 48038 46356 48044 46368
rect 47999 46328 48044 46356
rect 48038 46316 48044 46328
rect 48096 46316 48102 46368
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 3970 46112 3976 46164
rect 4028 46152 4034 46164
rect 4433 46155 4491 46161
rect 4433 46152 4445 46155
rect 4028 46124 4445 46152
rect 4028 46112 4034 46124
rect 4433 46121 4445 46124
rect 4479 46121 4491 46155
rect 5074 46152 5080 46164
rect 5035 46124 5080 46152
rect 4433 46115 4491 46121
rect 5074 46112 5080 46124
rect 5132 46112 5138 46164
rect 12158 46152 12164 46164
rect 12119 46124 12164 46152
rect 12158 46112 12164 46124
rect 12216 46112 12222 46164
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14182 46152 14188 46164
rect 14143 46124 14188 46152
rect 14182 46112 14188 46124
rect 14240 46112 14246 46164
rect 18598 46152 18604 46164
rect 18559 46124 18604 46152
rect 18598 46112 18604 46124
rect 18656 46112 18662 46164
rect 19242 46112 19248 46164
rect 19300 46152 19306 46164
rect 19429 46155 19487 46161
rect 19429 46152 19441 46155
rect 19300 46124 19441 46152
rect 19300 46112 19306 46124
rect 19429 46121 19441 46124
rect 19475 46121 19487 46155
rect 19429 46115 19487 46121
rect 24673 46155 24731 46161
rect 24673 46121 24685 46155
rect 24719 46152 24731 46155
rect 24762 46152 24768 46164
rect 24719 46124 24768 46152
rect 24719 46121 24731 46124
rect 24673 46115 24731 46121
rect 24762 46112 24768 46124
rect 24820 46112 24826 46164
rect 31849 46155 31907 46161
rect 31849 46121 31861 46155
rect 31895 46152 31907 46155
rect 32306 46152 32312 46164
rect 31895 46124 32312 46152
rect 31895 46121 31907 46124
rect 31849 46115 31907 46121
rect 32306 46112 32312 46124
rect 32364 46112 32370 46164
rect 38286 46152 38292 46164
rect 38247 46124 38292 46152
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 45002 46084 45008 46096
rect 35866 46056 45008 46084
rect 20714 46016 20720 46028
rect 12084 45988 18644 46016
rect 20675 45988 20720 46016
rect 1762 45908 1768 45960
rect 1820 45948 1826 45960
rect 2041 45951 2099 45957
rect 2041 45948 2053 45951
rect 1820 45920 2053 45948
rect 1820 45908 1826 45920
rect 2041 45917 2053 45920
rect 2087 45917 2099 45951
rect 2041 45911 2099 45917
rect 4985 45951 5043 45957
rect 4985 45917 4997 45951
rect 5031 45948 5043 45951
rect 11606 45948 11612 45960
rect 5031 45920 11612 45948
rect 5031 45917 5043 45920
rect 4985 45911 5043 45917
rect 11606 45908 11612 45920
rect 11664 45908 11670 45960
rect 12084 45957 12112 45988
rect 12069 45951 12127 45957
rect 12069 45917 12081 45951
rect 12115 45917 12127 45951
rect 14090 45948 14096 45960
rect 14003 45920 14096 45948
rect 12069 45911 12127 45917
rect 14090 45908 14096 45920
rect 14148 45948 14154 45960
rect 18506 45948 18512 45960
rect 14148 45920 18512 45948
rect 14148 45908 14154 45920
rect 18506 45908 18512 45920
rect 18564 45908 18570 45960
rect 18616 45880 18644 45988
rect 20714 45976 20720 45988
rect 20772 45976 20778 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 25225 46019 25283 46025
rect 25225 45985 25237 46019
rect 25271 46016 25283 46019
rect 25498 46016 25504 46028
rect 25271 45988 25504 46016
rect 25271 45985 25283 45988
rect 25225 45979 25283 45985
rect 25498 45976 25504 45988
rect 25556 45976 25562 46028
rect 25774 46016 25780 46028
rect 25735 45988 25780 46016
rect 25774 45976 25780 45988
rect 25832 45976 25838 46028
rect 24578 45948 24584 45960
rect 24539 45920 24584 45948
rect 24578 45908 24584 45920
rect 24636 45908 24642 45960
rect 31754 45948 31760 45960
rect 31667 45920 31760 45948
rect 31754 45908 31760 45920
rect 31812 45948 31818 45960
rect 35866 45948 35894 46056
rect 45002 46044 45008 46056
rect 45060 46044 45066 46096
rect 41230 46016 41236 46028
rect 41191 45988 41236 46016
rect 41230 45976 41236 45988
rect 41288 45976 41294 46028
rect 41874 46016 41880 46028
rect 41835 45988 41880 46016
rect 41874 45976 41880 45988
rect 41932 45976 41938 46028
rect 47026 46016 47032 46028
rect 46987 45988 47032 46016
rect 47026 45976 47032 45988
rect 47084 45976 47090 46028
rect 31812 45920 35894 45948
rect 38197 45951 38255 45957
rect 31812 45908 31818 45920
rect 38197 45917 38209 45951
rect 38243 45948 38255 45951
rect 38243 45920 40816 45948
rect 38243 45917 38255 45920
rect 38197 45911 38255 45917
rect 20714 45880 20720 45892
rect 18616 45852 20720 45880
rect 20714 45840 20720 45852
rect 20772 45840 20778 45892
rect 20898 45880 20904 45892
rect 20859 45852 20904 45880
rect 20898 45840 20904 45852
rect 20956 45840 20962 45892
rect 25406 45880 25412 45892
rect 25367 45852 25412 45880
rect 25406 45840 25412 45852
rect 25464 45840 25470 45892
rect 40788 45824 40816 45920
rect 43806 45908 43812 45960
rect 43864 45948 43870 45960
rect 43993 45951 44051 45957
rect 43993 45948 44005 45951
rect 43864 45920 44005 45948
rect 43864 45908 43870 45920
rect 43993 45917 44005 45920
rect 44039 45917 44051 45951
rect 43993 45911 44051 45917
rect 45557 45951 45615 45957
rect 45557 45917 45569 45951
rect 45603 45948 45615 45951
rect 45738 45948 45744 45960
rect 45603 45920 45744 45948
rect 45603 45917 45615 45920
rect 45557 45911 45615 45917
rect 45738 45908 45744 45920
rect 45796 45908 45802 45960
rect 45830 45908 45836 45960
rect 45888 45948 45894 45960
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45888 45920 46305 45948
rect 45888 45908 45894 45920
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 41414 45880 41420 45892
rect 41375 45852 41420 45880
rect 41414 45840 41420 45852
rect 41472 45840 41478 45892
rect 44177 45883 44235 45889
rect 44177 45849 44189 45883
rect 44223 45880 44235 45883
rect 44266 45880 44272 45892
rect 44223 45852 44272 45880
rect 44223 45849 44235 45852
rect 44177 45843 44235 45849
rect 44266 45840 44272 45852
rect 44324 45840 44330 45892
rect 46474 45880 46480 45892
rect 45526 45852 45876 45880
rect 46435 45852 46480 45880
rect 40770 45772 40776 45824
rect 40828 45812 40834 45824
rect 45526 45812 45554 45852
rect 40828 45784 45554 45812
rect 40828 45772 40834 45784
rect 45646 45772 45652 45824
rect 45704 45812 45710 45824
rect 45741 45815 45799 45821
rect 45741 45812 45753 45815
rect 45704 45784 45753 45812
rect 45704 45772 45710 45784
rect 45741 45781 45753 45784
rect 45787 45781 45799 45815
rect 45848 45812 45876 45852
rect 46474 45840 46480 45852
rect 46532 45840 46538 45892
rect 46842 45812 46848 45824
rect 45848 45784 46848 45812
rect 45741 45775 45799 45781
rect 46842 45772 46848 45784
rect 46900 45772 46906 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 11606 45568 11612 45620
rect 11664 45608 11670 45620
rect 20898 45608 20904 45620
rect 11664 45580 20760 45608
rect 20859 45580 20904 45608
rect 11664 45568 11670 45580
rect 20732 45540 20760 45580
rect 20898 45568 20904 45580
rect 20956 45568 20962 45620
rect 24578 45608 24584 45620
rect 21008 45580 24584 45608
rect 21008 45540 21036 45580
rect 24578 45568 24584 45580
rect 24636 45568 24642 45620
rect 25406 45608 25412 45620
rect 25367 45580 25412 45608
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 41414 45608 41420 45620
rect 41375 45580 41420 45608
rect 41414 45568 41420 45580
rect 41472 45568 41478 45620
rect 42521 45611 42579 45617
rect 42521 45577 42533 45611
rect 42567 45608 42579 45611
rect 42610 45608 42616 45620
rect 42567 45580 42616 45608
rect 42567 45577 42579 45580
rect 42521 45571 42579 45577
rect 42610 45568 42616 45580
rect 42668 45568 42674 45620
rect 45094 45568 45100 45620
rect 45152 45608 45158 45620
rect 45554 45608 45560 45620
rect 45152 45580 45560 45608
rect 45152 45568 45158 45580
rect 45554 45568 45560 45580
rect 45612 45568 45618 45620
rect 46382 45568 46388 45620
rect 46440 45608 46446 45620
rect 46440 45580 47624 45608
rect 46440 45568 46446 45580
rect 43162 45540 43168 45552
rect 20732 45512 21036 45540
rect 43123 45512 43168 45540
rect 43162 45500 43168 45512
rect 43220 45500 43226 45552
rect 43901 45543 43959 45549
rect 43901 45509 43913 45543
rect 43947 45540 43959 45543
rect 44174 45540 44180 45552
rect 43947 45512 44180 45540
rect 43947 45509 43959 45512
rect 43901 45503 43959 45509
rect 44174 45500 44180 45512
rect 44232 45500 44238 45552
rect 44284 45512 46612 45540
rect 1762 45472 1768 45484
rect 1723 45444 1768 45472
rect 1762 45432 1768 45444
rect 1820 45432 1826 45484
rect 20714 45432 20720 45484
rect 20772 45472 20778 45484
rect 20809 45475 20867 45481
rect 20809 45472 20821 45475
rect 20772 45444 20821 45472
rect 20772 45432 20778 45444
rect 20809 45441 20821 45444
rect 20855 45441 20867 45475
rect 25314 45472 25320 45484
rect 25275 45444 25320 45472
rect 20809 45435 20867 45441
rect 25314 45432 25320 45444
rect 25372 45432 25378 45484
rect 41046 45432 41052 45484
rect 41104 45472 41110 45484
rect 41325 45475 41383 45481
rect 41325 45472 41337 45475
rect 41104 45444 41337 45472
rect 41104 45432 41110 45444
rect 41325 45441 41337 45444
rect 41371 45441 41383 45475
rect 41325 45435 41383 45441
rect 42429 45475 42487 45481
rect 42429 45441 42441 45475
rect 42475 45441 42487 45475
rect 42429 45435 42487 45441
rect 43073 45475 43131 45481
rect 43073 45441 43085 45475
rect 43119 45472 43131 45475
rect 44284 45472 44312 45512
rect 43119 45444 44312 45472
rect 43119 45441 43131 45444
rect 43073 45435 43131 45441
rect 1949 45407 2007 45413
rect 1949 45373 1961 45407
rect 1995 45404 2007 45407
rect 2222 45404 2228 45416
rect 1995 45376 2228 45404
rect 1995 45373 2007 45376
rect 1949 45367 2007 45373
rect 2222 45364 2228 45376
rect 2280 45364 2286 45416
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 42444 45336 42472 45435
rect 44542 45404 44548 45416
rect 44503 45376 44548 45404
rect 44542 45364 44548 45376
rect 44600 45364 44606 45416
rect 44729 45407 44787 45413
rect 44729 45373 44741 45407
rect 44775 45404 44787 45407
rect 45094 45404 45100 45416
rect 44775 45376 45100 45404
rect 44775 45373 44787 45376
rect 44729 45367 44787 45373
rect 45094 45364 45100 45376
rect 45152 45364 45158 45416
rect 45554 45364 45560 45416
rect 45612 45404 45618 45416
rect 46584 45404 46612 45512
rect 46658 45500 46664 45552
rect 46716 45540 46722 45552
rect 46937 45543 46995 45549
rect 46937 45540 46949 45543
rect 46716 45512 46949 45540
rect 46716 45500 46722 45512
rect 46937 45509 46949 45512
rect 46983 45509 46995 45543
rect 46937 45503 46995 45509
rect 46842 45472 46848 45484
rect 46803 45444 46848 45472
rect 46842 45432 46848 45444
rect 46900 45432 46906 45484
rect 47596 45481 47624 45580
rect 47581 45475 47639 45481
rect 47581 45441 47593 45475
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 47118 45404 47124 45416
rect 45612 45376 45657 45404
rect 46584 45376 47124 45404
rect 45612 45364 45618 45376
rect 47118 45364 47124 45376
rect 47176 45364 47182 45416
rect 46382 45336 46388 45348
rect 42444 45308 46388 45336
rect 46382 45296 46388 45308
rect 46440 45296 46446 45348
rect 38470 45228 38476 45280
rect 38528 45268 38534 45280
rect 43993 45271 44051 45277
rect 43993 45268 44005 45271
rect 38528 45240 44005 45268
rect 38528 45228 38534 45240
rect 43993 45237 44005 45240
rect 44039 45237 44051 45271
rect 43993 45231 44051 45237
rect 47302 45228 47308 45280
rect 47360 45268 47366 45280
rect 47765 45271 47823 45277
rect 47765 45268 47777 45271
rect 47360 45240 47777 45268
rect 47360 45228 47366 45240
rect 47765 45237 47777 45240
rect 47811 45237 47823 45271
rect 47765 45231 47823 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 2222 45064 2228 45076
rect 2183 45036 2228 45064
rect 2222 45024 2228 45036
rect 2280 45024 2286 45076
rect 42702 45024 42708 45076
rect 42760 45064 42766 45076
rect 42981 45067 43039 45073
rect 42981 45064 42993 45067
rect 42760 45036 42993 45064
rect 42760 45024 42766 45036
rect 42981 45033 42993 45036
rect 43027 45033 43039 45067
rect 44450 45064 44456 45076
rect 44411 45036 44456 45064
rect 42981 45027 43039 45033
rect 44450 45024 44456 45036
rect 44508 45024 44514 45076
rect 45094 45064 45100 45076
rect 45055 45036 45100 45064
rect 45094 45024 45100 45036
rect 45152 45024 45158 45076
rect 45370 45024 45376 45076
rect 45428 45064 45434 45076
rect 45741 45067 45799 45073
rect 45741 45064 45753 45067
rect 45428 45036 45753 45064
rect 45428 45024 45434 45036
rect 45741 45033 45753 45036
rect 45787 45033 45799 45067
rect 45741 45027 45799 45033
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 47026 44928 47032 44940
rect 46339 44900 47032 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 47026 44888 47032 44900
rect 47084 44888 47090 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 2133 44863 2191 44869
rect 2133 44829 2145 44863
rect 2179 44860 2191 44863
rect 2406 44860 2412 44872
rect 2179 44832 2412 44860
rect 2179 44829 2191 44832
rect 2133 44823 2191 44829
rect 2406 44820 2412 44832
rect 2464 44820 2470 44872
rect 45002 44860 45008 44872
rect 44963 44832 45008 44860
rect 45002 44820 45008 44832
rect 45060 44860 45066 44872
rect 45554 44860 45560 44872
rect 45060 44832 45560 44860
rect 45060 44820 45066 44832
rect 45554 44820 45560 44832
rect 45612 44820 45618 44872
rect 45649 44863 45707 44869
rect 45649 44829 45661 44863
rect 45695 44860 45707 44863
rect 46198 44860 46204 44872
rect 45695 44832 46204 44860
rect 45695 44829 45707 44832
rect 45649 44823 45707 44829
rect 46198 44820 46204 44832
rect 46256 44820 46262 44872
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 47670 44792 47676 44804
rect 46523 44764 47676 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 47670 44752 47676 44764
rect 47728 44752 47734 44804
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 46293 44523 46351 44529
rect 46293 44489 46305 44523
rect 46339 44520 46351 44523
rect 46474 44520 46480 44532
rect 46339 44492 46480 44520
rect 46339 44489 46351 44492
rect 46293 44483 46351 44489
rect 46474 44480 46480 44492
rect 46532 44480 46538 44532
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 26206 44424 46244 44452
rect 24578 44344 24584 44396
rect 24636 44384 24642 44396
rect 26206 44384 26234 44424
rect 24636 44356 26234 44384
rect 24636 44344 24642 44356
rect 44542 44344 44548 44396
rect 44600 44384 44606 44396
rect 44821 44387 44879 44393
rect 44821 44384 44833 44387
rect 44600 44356 44833 44384
rect 44600 44344 44606 44356
rect 44821 44353 44833 44356
rect 44867 44353 44879 44387
rect 45738 44384 45744 44396
rect 45699 44356 45744 44384
rect 44821 44347 44879 44353
rect 45738 44344 45744 44356
rect 45796 44344 45802 44396
rect 46216 44393 46244 44424
rect 46201 44387 46259 44393
rect 46201 44353 46213 44387
rect 46247 44384 46259 44387
rect 46566 44384 46572 44396
rect 46247 44356 46572 44384
rect 46247 44353 46259 44356
rect 46201 44347 46259 44353
rect 46566 44344 46572 44356
rect 46624 44344 46630 44396
rect 46658 44344 46664 44396
rect 46716 44384 46722 44396
rect 46845 44387 46903 44393
rect 46845 44384 46857 44387
rect 46716 44356 46857 44384
rect 46716 44344 46722 44356
rect 46845 44353 46857 44356
rect 46891 44384 46903 44387
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 46891 44356 47593 44384
rect 46891 44353 46903 44356
rect 46845 44347 46903 44353
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 41046 44208 41052 44260
rect 41104 44248 41110 44260
rect 47578 44248 47584 44260
rect 41104 44220 47584 44248
rect 41104 44208 41110 44220
rect 47578 44208 47584 44220
rect 47636 44208 47642 44260
rect 20714 44140 20720 44192
rect 20772 44180 20778 44192
rect 21358 44180 21364 44192
rect 20772 44152 21364 44180
rect 20772 44140 20778 44152
rect 21358 44140 21364 44152
rect 21416 44140 21422 44192
rect 46934 44180 46940 44192
rect 46895 44152 46940 44180
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 46477 43843 46535 43849
rect 46477 43809 46489 43843
rect 46523 43840 46535 43843
rect 46934 43840 46940 43852
rect 46523 43812 46940 43840
rect 46523 43809 46535 43812
rect 46477 43803 46535 43809
rect 46934 43800 46940 43812
rect 46992 43800 46998 43852
rect 48133 43843 48191 43849
rect 48133 43809 48145 43843
rect 48179 43840 48191 43843
rect 48222 43840 48228 43852
rect 48179 43812 48228 43840
rect 48179 43809 48191 43812
rect 48133 43803 48191 43809
rect 48222 43800 48228 43812
rect 48280 43800 48286 43852
rect 45833 43775 45891 43781
rect 45833 43741 45845 43775
rect 45879 43772 45891 43775
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 45879 43744 46305 43772
rect 45879 43741 45891 43744
rect 45833 43735 45891 43741
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 47026 43296 47032 43308
rect 46987 43268 47032 43296
rect 47026 43256 47032 43268
rect 47084 43256 47090 43308
rect 47762 43296 47768 43308
rect 47723 43268 47768 43296
rect 47762 43256 47768 43268
rect 47820 43256 47826 43308
rect 1673 43231 1731 43237
rect 1673 43197 1685 43231
rect 1719 43228 1731 43231
rect 1946 43228 1952 43240
rect 1719 43200 1952 43228
rect 1719 43197 1731 43200
rect 1673 43191 1731 43197
rect 1946 43188 1952 43200
rect 2004 43188 2010 43240
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46290 42684 46296 42696
rect 46251 42656 46296 42684
rect 46290 42644 46296 42656
rect 46348 42644 46354 42696
rect 46477 42619 46535 42625
rect 46477 42585 46489 42619
rect 46523 42616 46535 42619
rect 47670 42616 47676 42628
rect 46523 42588 47676 42616
rect 46523 42585 46535 42588
rect 46477 42579 46535 42585
rect 47670 42576 47676 42588
rect 47728 42576 47734 42628
rect 48130 42616 48136 42628
rect 48091 42588 48136 42616
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 47670 42344 47676 42356
rect 47631 42316 47676 42344
rect 47670 42304 47676 42316
rect 47728 42304 47734 42356
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 47029 42211 47087 42217
rect 47029 42208 47041 42211
rect 46348 42180 47041 42208
rect 46348 42168 46354 42180
rect 47029 42177 47041 42180
rect 47075 42177 47087 42211
rect 47029 42171 47087 42177
rect 47581 42211 47639 42217
rect 47581 42177 47593 42211
rect 47627 42177 47639 42211
rect 47581 42171 47639 42177
rect 46934 42100 46940 42152
rect 46992 42140 46998 42152
rect 47118 42140 47124 42152
rect 46992 42112 47124 42140
rect 46992 42100 46998 42112
rect 47118 42100 47124 42112
rect 47176 42140 47182 42152
rect 47596 42140 47624 42171
rect 47176 42112 47624 42140
rect 47176 42100 47182 42112
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47762 41664 47768 41676
rect 46339 41636 47768 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47762 41624 47768 41636
rect 47820 41624 47826 41676
rect 27341 41599 27399 41605
rect 27341 41565 27353 41599
rect 27387 41596 27399 41599
rect 31754 41596 31760 41608
rect 27387 41568 31760 41596
rect 27387 41565 27399 41568
rect 27341 41559 27399 41565
rect 31754 41556 31760 41568
rect 31812 41556 31818 41608
rect 48130 41596 48136 41608
rect 48091 41568 48136 41596
rect 48130 41556 48136 41568
rect 48188 41556 48194 41608
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 46474 41528 46480 41540
rect 46435 41500 46480 41528
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 27154 41420 27160 41472
rect 27212 41460 27218 41472
rect 27433 41463 27491 41469
rect 27433 41460 27445 41463
rect 27212 41432 27445 41460
rect 27212 41420 27218 41432
rect 27433 41429 27445 41432
rect 27479 41429 27491 41463
rect 27433 41423 27491 41429
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2133 41259 2191 41265
rect 2133 41256 2145 41259
rect 1636 41228 2145 41256
rect 1636 41216 1642 41228
rect 2133 41225 2145 41228
rect 2179 41225 2191 41259
rect 2133 41219 2191 41225
rect 26234 41216 26240 41268
rect 26292 41256 26298 41268
rect 26292 41228 28856 41256
rect 26292 41216 26298 41228
rect 27154 41188 27160 41200
rect 27115 41160 27160 41188
rect 27154 41148 27160 41160
rect 27212 41148 27218 41200
rect 28828 41197 28856 41228
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46753 41259 46811 41265
rect 46753 41256 46765 41259
rect 46532 41228 46765 41256
rect 46532 41216 46538 41228
rect 46753 41225 46765 41228
rect 46799 41225 46811 41259
rect 46753 41219 46811 41225
rect 28813 41191 28871 41197
rect 28813 41157 28825 41191
rect 28859 41157 28871 41191
rect 28813 41151 28871 41157
rect 2041 41123 2099 41129
rect 2041 41089 2053 41123
rect 2087 41120 2099 41123
rect 14090 41120 14096 41132
rect 2087 41092 14096 41120
rect 2087 41089 2099 41092
rect 2041 41083 2099 41089
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 46382 41080 46388 41132
rect 46440 41120 46446 41132
rect 46661 41123 46719 41129
rect 46661 41120 46673 41123
rect 46440 41092 46673 41120
rect 46440 41080 46446 41092
rect 46661 41089 46673 41092
rect 46707 41089 46719 41123
rect 47762 41120 47768 41132
rect 47723 41092 47768 41120
rect 46661 41083 46719 41089
rect 47762 41080 47768 41092
rect 47820 41080 47826 41132
rect 26050 41012 26056 41064
rect 26108 41052 26114 41064
rect 26973 41055 27031 41061
rect 26973 41052 26985 41055
rect 26108 41024 26985 41052
rect 26108 41012 26114 41024
rect 26973 41021 26985 41024
rect 27019 41052 27031 41055
rect 42794 41052 42800 41064
rect 27019 41024 31754 41052
rect 27019 41021 27031 41024
rect 26973 41015 27031 41021
rect 31726 40984 31754 41024
rect 35866 41024 42800 41052
rect 35866 40984 35894 41024
rect 42794 41012 42800 41024
rect 42852 41012 42858 41064
rect 31726 40956 35894 40984
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 46845 40647 46903 40653
rect 46845 40644 46857 40647
rect 45526 40616 46857 40644
rect 26050 40576 26056 40588
rect 26011 40548 26056 40576
rect 26050 40536 26056 40548
rect 26108 40536 26114 40588
rect 45526 40576 45554 40616
rect 46845 40613 46857 40616
rect 46891 40613 46903 40647
rect 46845 40607 46903 40613
rect 45480 40548 45554 40576
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 45094 40508 45100 40520
rect 45055 40480 45100 40508
rect 45094 40468 45100 40480
rect 45152 40468 45158 40520
rect 45480 40517 45508 40548
rect 45465 40511 45523 40517
rect 45465 40477 45477 40511
rect 45511 40477 45523 40511
rect 45465 40471 45523 40477
rect 46842 40468 46848 40520
rect 46900 40508 46906 40520
rect 47029 40511 47087 40517
rect 47029 40508 47041 40511
rect 46900 40480 47041 40508
rect 46900 40468 46906 40480
rect 47029 40477 47041 40480
rect 47075 40477 47087 40511
rect 47670 40508 47676 40520
rect 47631 40480 47676 40508
rect 47029 40471 47087 40477
rect 47670 40468 47676 40480
rect 47728 40468 47734 40520
rect 2130 40400 2136 40452
rect 2188 40440 2194 40452
rect 26237 40443 26295 40449
rect 26237 40440 26249 40443
rect 2188 40412 26249 40440
rect 2188 40400 2194 40412
rect 26237 40409 26249 40412
rect 26283 40409 26295 40443
rect 26237 40403 26295 40409
rect 27893 40443 27951 40449
rect 27893 40409 27905 40443
rect 27939 40440 27951 40443
rect 28074 40440 28080 40452
rect 27939 40412 28080 40440
rect 27939 40409 27951 40412
rect 27893 40403 27951 40409
rect 28074 40400 28080 40412
rect 28132 40400 28138 40452
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40372 1639 40375
rect 1854 40372 1860 40384
rect 1627 40344 1860 40372
rect 1627 40341 1639 40344
rect 1581 40335 1639 40341
rect 1854 40332 1860 40344
rect 1912 40332 1918 40384
rect 46106 40372 46112 40384
rect 46067 40344 46112 40372
rect 46106 40332 46112 40344
rect 46164 40332 46170 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 45922 40100 45928 40112
rect 45848 40072 45928 40100
rect 45848 40041 45876 40072
rect 45922 40060 45928 40072
rect 45980 40060 45986 40112
rect 45833 40035 45891 40041
rect 45833 40001 45845 40035
rect 45879 40001 45891 40035
rect 46106 40032 46112 40044
rect 46067 40004 46112 40032
rect 45833 39995 45891 40001
rect 46106 39992 46112 40004
rect 46164 39992 46170 40044
rect 47578 40032 47584 40044
rect 47539 40004 47584 40032
rect 47578 39992 47584 40004
rect 47636 39992 47642 40044
rect 42794 39856 42800 39908
rect 42852 39896 42858 39908
rect 46109 39899 46167 39905
rect 46109 39896 46121 39899
rect 42852 39868 46121 39896
rect 42852 39856 42858 39868
rect 46109 39865 46121 39868
rect 46155 39865 46167 39899
rect 46109 39859 46167 39865
rect 46474 39788 46480 39840
rect 46532 39828 46538 39840
rect 47673 39831 47731 39837
rect 47673 39828 47685 39831
rect 46532 39800 47685 39828
rect 46532 39788 46538 39800
rect 47673 39797 47685 39800
rect 47719 39797 47731 39831
rect 47673 39791 47731 39797
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 47670 39556 47676 39568
rect 46308 39528 47676 39556
rect 46308 39497 46336 39528
rect 47670 39516 47676 39528
rect 47728 39516 47734 39568
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39457 46351 39491
rect 46474 39488 46480 39500
rect 46435 39460 46480 39488
rect 46293 39451 46351 39457
rect 46474 39448 46480 39460
rect 46532 39448 46538 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 45189 39083 45247 39089
rect 45189 39049 45201 39083
rect 45235 39080 45247 39083
rect 45235 39052 45876 39080
rect 45235 39049 45247 39052
rect 45189 39043 45247 39049
rect 45848 38956 45876 39052
rect 42058 38904 42064 38956
rect 42116 38944 42122 38956
rect 45005 38947 45063 38953
rect 45005 38944 45017 38947
rect 42116 38916 45017 38944
rect 42116 38904 42122 38916
rect 45005 38913 45017 38916
rect 45051 38913 45063 38947
rect 45830 38944 45836 38956
rect 45791 38916 45836 38944
rect 45005 38907 45063 38913
rect 45020 38808 45048 38907
rect 45830 38904 45836 38916
rect 45888 38904 45894 38956
rect 47854 38944 47860 38956
rect 47815 38916 47860 38944
rect 47854 38904 47860 38916
rect 47912 38904 47918 38956
rect 46385 38879 46443 38885
rect 46385 38845 46397 38879
rect 46431 38876 46443 38879
rect 46658 38876 46664 38888
rect 46431 38848 46664 38876
rect 46431 38845 46443 38848
rect 46385 38839 46443 38845
rect 46658 38836 46664 38848
rect 46716 38836 46722 38888
rect 48041 38811 48099 38817
rect 48041 38808 48053 38811
rect 45020 38780 48053 38808
rect 48041 38777 48053 38780
rect 48087 38777 48099 38811
rect 48041 38771 48099 38777
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 45554 38360 45560 38412
rect 45612 38400 45618 38412
rect 46014 38400 46020 38412
rect 45612 38372 46020 38400
rect 45612 38360 45618 38372
rect 46014 38360 46020 38372
rect 46072 38360 46078 38412
rect 45189 38335 45247 38341
rect 45189 38301 45201 38335
rect 45235 38332 45247 38335
rect 45830 38332 45836 38344
rect 45235 38304 45836 38332
rect 45235 38301 45247 38304
rect 45189 38295 45247 38301
rect 45830 38292 45836 38304
rect 45888 38292 45894 38344
rect 46290 38332 46296 38344
rect 46251 38304 46296 38332
rect 46290 38292 46296 38304
rect 46348 38292 46354 38344
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 47670 38264 47676 38276
rect 46523 38236 47676 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 47670 38224 47676 38236
rect 47728 38224 47734 38276
rect 48130 38264 48136 38276
rect 48091 38236 48136 38264
rect 48130 38224 48136 38236
rect 48188 38224 48194 38276
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 47670 37992 47676 38004
rect 47631 37964 47676 37992
rect 47670 37952 47676 37964
rect 47728 37952 47734 38004
rect 25314 37884 25320 37936
rect 25372 37924 25378 37936
rect 25372 37896 47532 37924
rect 25372 37884 25378 37896
rect 47504 37868 47532 37896
rect 45830 37856 45836 37868
rect 45791 37828 45836 37856
rect 45830 37816 45836 37828
rect 45888 37816 45894 37868
rect 47486 37816 47492 37868
rect 47544 37856 47550 37868
rect 47581 37859 47639 37865
rect 47581 37856 47593 37859
rect 47544 37828 47593 37856
rect 47544 37816 47550 37828
rect 47581 37825 47593 37828
rect 47627 37825 47639 37859
rect 47581 37819 47639 37825
rect 46198 37788 46204 37800
rect 46159 37760 46204 37788
rect 46198 37748 46204 37760
rect 46256 37748 46262 37800
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 46290 37408 46296 37460
rect 46348 37448 46354 37460
rect 47673 37451 47731 37457
rect 47673 37448 47685 37451
rect 46348 37420 47685 37448
rect 46348 37408 46354 37420
rect 47673 37417 47685 37420
rect 47719 37417 47731 37451
rect 47673 37411 47731 37417
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 1820 37216 2053 37244
rect 1820 37204 1826 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 45830 37244 45836 37256
rect 45791 37216 45836 37244
rect 2041 37207 2099 37213
rect 45830 37204 45836 37216
rect 45888 37204 45894 37256
rect 46385 37179 46443 37185
rect 46385 37145 46397 37179
rect 46431 37176 46443 37179
rect 46566 37176 46572 37188
rect 46431 37148 46572 37176
rect 46431 37145 46443 37148
rect 46385 37139 46443 37145
rect 46566 37136 46572 37148
rect 46624 37136 46630 37188
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 46382 36836 46388 36848
rect 46343 36808 46388 36836
rect 46382 36796 46388 36808
rect 46440 36796 46446 36848
rect 1762 36768 1768 36780
rect 1723 36740 1768 36768
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 45830 36768 45836 36780
rect 45791 36740 45836 36768
rect 45830 36728 45836 36740
rect 45888 36728 45894 36780
rect 1949 36703 2007 36709
rect 1949 36669 1961 36703
rect 1995 36700 2007 36703
rect 2222 36700 2228 36712
rect 1995 36672 2228 36700
rect 1995 36669 2007 36672
rect 1949 36663 2007 36669
rect 2222 36660 2228 36672
rect 2280 36660 2286 36712
rect 2774 36700 2780 36712
rect 2735 36672 2780 36700
rect 2774 36660 2780 36672
rect 2832 36660 2838 36712
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 2130 36156 2136 36168
rect 2043 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36156 2194 36168
rect 46198 36156 46204 36168
rect 2188 36128 46204 36156
rect 2188 36116 2194 36128
rect 46198 36116 46204 36128
rect 46256 36116 46262 36168
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 1486 35476 1492 35488
rect 1443 35448 1492 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 1486 35436 1492 35448
rect 1544 35436 1550 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 48130 35068 48136 35080
rect 48091 35040 48136 35068
rect 48130 35028 48136 35040
rect 48188 35028 48194 35080
rect 47118 34892 47124 34944
rect 47176 34932 47182 34944
rect 47949 34935 48007 34941
rect 47949 34932 47961 34935
rect 47176 34904 47961 34932
rect 47176 34892 47182 34904
rect 47949 34901 47961 34904
rect 47995 34901 48007 34935
rect 47949 34895 48007 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34592 29607 34595
rect 30558 34592 30564 34604
rect 29595 34564 30420 34592
rect 30519 34564 30564 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 29638 34524 29644 34536
rect 29599 34496 29644 34524
rect 29638 34484 29644 34496
rect 29696 34484 29702 34536
rect 30392 34524 30420 34564
rect 30558 34552 30564 34564
rect 30616 34552 30622 34604
rect 48130 34592 48136 34604
rect 48091 34564 48136 34592
rect 48130 34552 48136 34564
rect 48188 34552 48194 34604
rect 31754 34524 31760 34536
rect 30392 34496 31760 34524
rect 31754 34484 31760 34496
rect 31812 34484 31818 34536
rect 30374 34388 30380 34400
rect 30335 34360 30380 34388
rect 30374 34348 30380 34360
rect 30432 34348 30438 34400
rect 47210 34348 47216 34400
rect 47268 34388 47274 34400
rect 47949 34391 48007 34397
rect 47949 34388 47961 34391
rect 47268 34360 47961 34388
rect 47268 34348 47274 34360
rect 47949 34357 47961 34360
rect 47995 34357 48007 34391
rect 47949 34351 48007 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 45830 34076 45836 34128
rect 45888 34116 45894 34128
rect 45888 34088 47440 34116
rect 45888 34076 45894 34088
rect 24670 34008 24676 34060
rect 24728 34048 24734 34060
rect 24949 34051 25007 34057
rect 24949 34048 24961 34051
rect 24728 34020 24961 34048
rect 24728 34008 24734 34020
rect 24949 34017 24961 34020
rect 24995 34017 25007 34051
rect 24949 34011 25007 34017
rect 30009 34051 30067 34057
rect 30009 34017 30021 34051
rect 30055 34048 30067 34051
rect 32214 34048 32220 34060
rect 30055 34020 32220 34048
rect 30055 34017 30067 34020
rect 30009 34011 30067 34017
rect 32214 34008 32220 34020
rect 32272 34008 32278 34060
rect 47118 34048 47124 34060
rect 47079 34020 47124 34048
rect 47118 34008 47124 34020
rect 47176 34008 47182 34060
rect 47412 34057 47440 34088
rect 47397 34051 47455 34057
rect 47397 34017 47409 34051
rect 47443 34017 47455 34051
rect 47397 34011 47455 34017
rect 1302 33940 1308 33992
rect 1360 33980 1366 33992
rect 1581 33983 1639 33989
rect 1581 33980 1593 33983
rect 1360 33952 1593 33980
rect 1360 33940 1366 33952
rect 1581 33949 1593 33952
rect 1627 33949 1639 33983
rect 1581 33943 1639 33949
rect 20438 33940 20444 33992
rect 20496 33980 20502 33992
rect 20533 33983 20591 33989
rect 20533 33980 20545 33983
rect 20496 33952 20545 33980
rect 20496 33940 20502 33952
rect 20533 33949 20545 33952
rect 20579 33949 20591 33983
rect 20533 33943 20591 33949
rect 20809 33915 20867 33921
rect 20809 33881 20821 33915
rect 20855 33912 20867 33915
rect 21082 33912 21088 33924
rect 20855 33884 21088 33912
rect 20855 33881 20867 33884
rect 20809 33875 20867 33881
rect 21082 33872 21088 33884
rect 21140 33872 21146 33924
rect 21542 33872 21548 33924
rect 21600 33872 21606 33924
rect 24486 33872 24492 33924
rect 24544 33912 24550 33924
rect 24857 33915 24915 33921
rect 24857 33912 24869 33915
rect 24544 33884 24869 33912
rect 24544 33872 24550 33884
rect 24857 33881 24869 33884
rect 24903 33881 24915 33915
rect 24857 33875 24915 33881
rect 30285 33915 30343 33921
rect 30285 33881 30297 33915
rect 30331 33912 30343 33915
rect 30374 33912 30380 33924
rect 30331 33884 30380 33912
rect 30331 33881 30343 33884
rect 30285 33875 30343 33881
rect 30374 33872 30380 33884
rect 30432 33872 30438 33924
rect 31846 33912 31852 33924
rect 31510 33884 31852 33912
rect 31846 33872 31852 33884
rect 31904 33872 31910 33924
rect 47210 33872 47216 33924
rect 47268 33912 47274 33924
rect 47268 33884 47313 33912
rect 47268 33872 47274 33884
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 1578 33844 1584 33856
rect 1443 33816 1584 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 22278 33844 22284 33856
rect 22239 33816 22284 33844
rect 22278 33804 22284 33816
rect 22336 33804 22342 33856
rect 23474 33804 23480 33856
rect 23532 33844 23538 33856
rect 24397 33847 24455 33853
rect 24397 33844 24409 33847
rect 23532 33816 24409 33844
rect 23532 33804 23538 33816
rect 24397 33813 24409 33816
rect 24443 33813 24455 33847
rect 24762 33844 24768 33856
rect 24723 33816 24768 33844
rect 24397 33807 24455 33813
rect 24762 33804 24768 33816
rect 24820 33804 24826 33856
rect 31662 33804 31668 33856
rect 31720 33844 31726 33856
rect 31757 33847 31815 33853
rect 31757 33844 31769 33847
rect 31720 33816 31769 33844
rect 31720 33804 31726 33816
rect 31757 33813 31769 33816
rect 31803 33813 31815 33847
rect 31757 33807 31815 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 11698 33600 11704 33652
rect 11756 33640 11762 33652
rect 30469 33643 30527 33649
rect 30469 33640 30481 33643
rect 11756 33612 23244 33640
rect 11756 33600 11762 33612
rect 14642 33532 14648 33584
rect 14700 33572 14706 33584
rect 22373 33575 22431 33581
rect 22373 33572 22385 33575
rect 14700 33544 22385 33572
rect 14700 33532 14706 33544
rect 22373 33541 22385 33544
rect 22419 33541 22431 33575
rect 23216 33572 23244 33612
rect 24596 33612 30481 33640
rect 24596 33572 24624 33612
rect 30469 33609 30481 33612
rect 30515 33640 30527 33643
rect 31205 33643 31263 33649
rect 31205 33640 31217 33643
rect 30515 33612 31217 33640
rect 30515 33609 30527 33612
rect 30469 33603 30527 33609
rect 31205 33609 31217 33612
rect 31251 33609 31263 33643
rect 31205 33603 31263 33609
rect 31297 33643 31355 33649
rect 31297 33609 31309 33643
rect 31343 33640 31355 33643
rect 32677 33643 32735 33649
rect 32677 33640 32689 33643
rect 31343 33612 32689 33640
rect 31343 33609 31355 33612
rect 31297 33603 31355 33609
rect 32677 33609 32689 33612
rect 32723 33609 32735 33643
rect 32677 33603 32735 33609
rect 25682 33572 25688 33584
rect 23216 33544 24624 33572
rect 25438 33544 25688 33572
rect 22373 33535 22431 33541
rect 25682 33532 25688 33544
rect 25740 33532 25746 33584
rect 29638 33572 29644 33584
rect 29394 33544 29644 33572
rect 29638 33532 29644 33544
rect 29696 33532 29702 33584
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33504 19395 33507
rect 19426 33504 19432 33516
rect 19383 33476 19432 33504
rect 19383 33473 19395 33476
rect 19337 33467 19395 33473
rect 19426 33464 19432 33476
rect 19484 33464 19490 33516
rect 21266 33504 21272 33516
rect 21227 33476 21272 33504
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 23474 33504 23480 33516
rect 23435 33476 23480 33504
rect 23474 33464 23480 33476
rect 23532 33464 23538 33516
rect 29914 33464 29920 33516
rect 29972 33504 29978 33516
rect 30009 33507 30067 33513
rect 30009 33504 30021 33507
rect 29972 33476 30021 33504
rect 29972 33464 29978 33476
rect 30009 33473 30021 33476
rect 30055 33473 30067 33507
rect 30009 33467 30067 33473
rect 30193 33507 30251 33513
rect 30193 33473 30205 33507
rect 30239 33473 30251 33507
rect 30193 33467 30251 33473
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2314 33436 2320 33448
rect 1719 33408 2320 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2314 33396 2320 33408
rect 2372 33396 2378 33448
rect 22462 33436 22468 33448
rect 22423 33408 22468 33436
rect 22462 33396 22468 33408
rect 22520 33396 22526 33448
rect 22649 33439 22707 33445
rect 22649 33405 22661 33439
rect 22695 33436 22707 33439
rect 23566 33436 23572 33448
rect 22695 33408 23572 33436
rect 22695 33405 22707 33408
rect 22649 33399 22707 33405
rect 23566 33396 23572 33408
rect 23624 33396 23630 33448
rect 23934 33436 23940 33448
rect 23895 33408 23940 33436
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 24213 33439 24271 33445
rect 24213 33436 24225 33439
rect 24044 33408 24225 33436
rect 20438 33328 20444 33380
rect 20496 33368 20502 33380
rect 23952 33368 23980 33396
rect 20496 33340 23980 33368
rect 20496 33328 20502 33340
rect 19334 33260 19340 33312
rect 19392 33300 19398 33312
rect 19429 33303 19487 33309
rect 19429 33300 19441 33303
rect 19392 33272 19441 33300
rect 19392 33260 19398 33272
rect 19429 33269 19441 33272
rect 19475 33269 19487 33303
rect 21082 33300 21088 33312
rect 21043 33272 21088 33300
rect 19429 33263 19487 33269
rect 21082 33260 21088 33272
rect 21140 33260 21146 33312
rect 22002 33300 22008 33312
rect 21963 33272 22008 33300
rect 22002 33260 22008 33272
rect 22060 33260 22066 33312
rect 23293 33303 23351 33309
rect 23293 33269 23305 33303
rect 23339 33300 23351 33303
rect 24044 33300 24072 33408
rect 24213 33405 24225 33408
rect 24259 33405 24271 33439
rect 24213 33399 24271 33405
rect 27246 33396 27252 33448
rect 27304 33436 27310 33448
rect 27893 33439 27951 33445
rect 27893 33436 27905 33439
rect 27304 33408 27905 33436
rect 27304 33396 27310 33408
rect 27893 33405 27905 33408
rect 27939 33405 27951 33439
rect 28166 33436 28172 33448
rect 28127 33408 28172 33436
rect 27893 33399 27951 33405
rect 28166 33396 28172 33408
rect 28224 33396 28230 33448
rect 29822 33396 29828 33448
rect 29880 33436 29886 33448
rect 30208 33436 30236 33467
rect 31662 33464 31668 33516
rect 31720 33504 31726 33516
rect 32309 33507 32367 33513
rect 32309 33504 32321 33507
rect 31720 33476 32321 33504
rect 31720 33464 31726 33476
rect 32309 33473 32321 33476
rect 32355 33473 32367 33507
rect 47762 33504 47768 33516
rect 47723 33476 47768 33504
rect 32309 33467 32367 33473
rect 47762 33464 47768 33476
rect 47820 33464 47826 33516
rect 29880 33408 30236 33436
rect 29880 33396 29886 33408
rect 30208 33368 30236 33408
rect 31481 33439 31539 33445
rect 31481 33405 31493 33439
rect 31527 33436 31539 33439
rect 32122 33436 32128 33448
rect 31527 33408 32128 33436
rect 31527 33405 31539 33408
rect 31481 33399 31539 33405
rect 32122 33396 32128 33408
rect 32180 33396 32186 33448
rect 32217 33439 32275 33445
rect 32217 33405 32229 33439
rect 32263 33405 32275 33439
rect 32217 33399 32275 33405
rect 32232 33368 32260 33399
rect 30208 33340 32260 33368
rect 23339 33272 24072 33300
rect 23339 33269 23351 33272
rect 23293 33263 23351 33269
rect 24762 33260 24768 33312
rect 24820 33300 24826 33312
rect 25685 33303 25743 33309
rect 25685 33300 25697 33303
rect 24820 33272 25697 33300
rect 24820 33260 24826 33272
rect 25685 33269 25697 33272
rect 25731 33269 25743 33303
rect 29638 33300 29644 33312
rect 29599 33272 29644 33300
rect 25685 33263 25743 33269
rect 29638 33260 29644 33272
rect 29696 33260 29702 33312
rect 29730 33260 29736 33312
rect 29788 33300 29794 33312
rect 30009 33303 30067 33309
rect 30009 33300 30021 33303
rect 29788 33272 30021 33300
rect 29788 33260 29794 33272
rect 30009 33269 30021 33272
rect 30055 33269 30067 33303
rect 30834 33300 30840 33312
rect 30795 33272 30840 33300
rect 30009 33263 30067 33269
rect 30834 33260 30840 33272
rect 30892 33260 30898 33312
rect 47854 33300 47860 33312
rect 47815 33272 47860 33300
rect 47854 33260 47860 33272
rect 47912 33260 47918 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 18601 33099 18659 33105
rect 18601 33065 18613 33099
rect 18647 33096 18659 33099
rect 19150 33096 19156 33108
rect 18647 33068 19156 33096
rect 18647 33065 18659 33068
rect 18601 33059 18659 33065
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 21266 33056 21272 33108
rect 21324 33096 21330 33108
rect 21637 33099 21695 33105
rect 21637 33096 21649 33099
rect 21324 33068 21649 33096
rect 21324 33056 21330 33068
rect 21637 33065 21649 33068
rect 21683 33065 21695 33099
rect 21637 33059 21695 33065
rect 24397 33099 24455 33105
rect 24397 33065 24409 33099
rect 24443 33096 24455 33099
rect 24486 33096 24492 33108
rect 24443 33068 24492 33096
rect 24443 33065 24455 33068
rect 24397 33059 24455 33065
rect 24486 33056 24492 33068
rect 24544 33056 24550 33108
rect 24578 33056 24584 33108
rect 24636 33096 24642 33108
rect 25682 33096 25688 33108
rect 24636 33068 24992 33096
rect 25643 33068 25688 33096
rect 24636 33056 24642 33068
rect 1486 33028 1492 33040
rect 1412 33000 1492 33028
rect 1412 32969 1440 33000
rect 1486 32988 1492 33000
rect 1544 32988 1550 33040
rect 1854 32988 1860 33040
rect 1912 33028 1918 33040
rect 24854 33028 24860 33040
rect 1912 33000 24860 33028
rect 1912 32988 1918 33000
rect 24854 32988 24860 33000
rect 24912 32988 24918 33040
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32929 1455 32963
rect 1578 32960 1584 32972
rect 1539 32932 1584 32960
rect 1397 32923 1455 32929
rect 1578 32920 1584 32932
rect 1636 32920 1642 32972
rect 19426 32960 19432 32972
rect 18524 32932 19432 32960
rect 12437 32895 12495 32901
rect 12437 32861 12449 32895
rect 12483 32892 12495 32895
rect 12526 32892 12532 32904
rect 12483 32864 12532 32892
rect 12483 32861 12495 32864
rect 12437 32855 12495 32861
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 12618 32852 12624 32904
rect 12676 32892 12682 32904
rect 18524 32901 18552 32932
rect 19426 32920 19432 32932
rect 19484 32920 19490 32972
rect 22002 32920 22008 32972
rect 22060 32960 22066 32972
rect 22097 32963 22155 32969
rect 22097 32960 22109 32963
rect 22060 32932 22109 32960
rect 22060 32920 22066 32932
rect 22097 32929 22109 32932
rect 22143 32929 22155 32963
rect 22097 32923 22155 32929
rect 22281 32963 22339 32969
rect 22281 32929 22293 32963
rect 22327 32929 22339 32963
rect 22281 32923 22339 32929
rect 18509 32895 18567 32901
rect 12676 32864 12721 32892
rect 12676 32852 12682 32864
rect 18509 32861 18521 32895
rect 18555 32861 18567 32895
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18509 32855 18567 32861
rect 18800 32864 19257 32892
rect 3234 32824 3240 32836
rect 3195 32796 3240 32824
rect 3234 32784 3240 32796
rect 3292 32784 3298 32836
rect 11974 32716 11980 32768
rect 12032 32756 12038 32768
rect 12529 32759 12587 32765
rect 12529 32756 12541 32759
rect 12032 32728 12541 32756
rect 12032 32716 12038 32728
rect 12529 32725 12541 32728
rect 12575 32725 12587 32759
rect 12529 32719 12587 32725
rect 17770 32716 17776 32768
rect 17828 32756 17834 32768
rect 18800 32756 18828 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 22296 32892 22324 32923
rect 22738 32920 22744 32972
rect 22796 32960 22802 32972
rect 24964 32969 24992 33068
rect 25682 33056 25688 33068
rect 25740 33056 25746 33108
rect 28166 33056 28172 33108
rect 28224 33096 28230 33108
rect 28629 33099 28687 33105
rect 28629 33096 28641 33099
rect 28224 33068 28641 33096
rect 28224 33056 28230 33068
rect 28629 33065 28641 33068
rect 28675 33065 28687 33099
rect 30558 33096 30564 33108
rect 30519 33068 30564 33096
rect 28629 33059 28687 33065
rect 30558 33056 30564 33068
rect 30616 33056 30622 33108
rect 31846 33096 31852 33108
rect 31807 33068 31852 33096
rect 31846 33056 31852 33068
rect 31904 33056 31910 33108
rect 31938 33056 31944 33108
rect 31996 33096 32002 33108
rect 37274 33096 37280 33108
rect 31996 33068 37280 33096
rect 31996 33056 32002 33068
rect 37274 33056 37280 33068
rect 37332 33056 37338 33108
rect 25038 32988 25044 33040
rect 25096 32988 25102 33040
rect 31110 32988 31116 33040
rect 31168 33028 31174 33040
rect 35066 33028 35072 33040
rect 31168 33000 35072 33028
rect 31168 32988 31174 33000
rect 35066 32988 35072 33000
rect 35124 32988 35130 33040
rect 35713 33031 35771 33037
rect 35713 32997 35725 33031
rect 35759 33028 35771 33031
rect 37458 33028 37464 33040
rect 35759 33000 37464 33028
rect 35759 32997 35771 33000
rect 35713 32991 35771 32997
rect 37458 32988 37464 33000
rect 37516 32988 37522 33040
rect 24949 32963 25007 32969
rect 22796 32932 24808 32960
rect 22796 32920 22802 32932
rect 22833 32895 22891 32901
rect 22833 32892 22845 32895
rect 22296 32864 22845 32892
rect 19245 32855 19303 32861
rect 22833 32861 22845 32864
rect 22879 32892 22891 32895
rect 23382 32892 23388 32904
rect 22879 32864 23388 32892
rect 22879 32861 22891 32864
rect 22833 32855 22891 32861
rect 23382 32852 23388 32864
rect 23440 32852 23446 32904
rect 23566 32892 23572 32904
rect 23527 32864 23572 32892
rect 23566 32852 23572 32864
rect 23624 32892 23630 32904
rect 24026 32892 24032 32904
rect 23624 32864 24032 32892
rect 23624 32852 23630 32864
rect 24026 32852 24032 32864
rect 24084 32892 24090 32904
rect 24578 32892 24584 32904
rect 24084 32864 24584 32892
rect 24084 32852 24090 32864
rect 24578 32852 24584 32864
rect 24636 32852 24642 32904
rect 24780 32901 24808 32932
rect 24949 32929 24961 32963
rect 24995 32929 25007 32963
rect 25056 32960 25084 32988
rect 28261 32963 28319 32969
rect 28261 32960 28273 32963
rect 25056 32932 28273 32960
rect 24949 32923 25007 32929
rect 28261 32929 28273 32932
rect 28307 32929 28319 32963
rect 29638 32960 29644 32972
rect 28261 32923 28319 32929
rect 28368 32932 29644 32960
rect 24765 32895 24823 32901
rect 24765 32861 24777 32895
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25038 32892 25044 32904
rect 24903 32864 25044 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 25593 32895 25651 32901
rect 25593 32861 25605 32895
rect 25639 32892 25651 32895
rect 26326 32892 26332 32904
rect 25639 32864 26332 32892
rect 25639 32861 25651 32864
rect 25593 32855 25651 32861
rect 26326 32852 26332 32864
rect 26384 32852 26390 32904
rect 27890 32892 27896 32904
rect 27851 32864 27896 32892
rect 27890 32852 27896 32864
rect 27948 32852 27954 32904
rect 27982 32852 27988 32904
rect 28040 32892 28046 32904
rect 28077 32895 28135 32901
rect 28077 32892 28089 32895
rect 28040 32864 28089 32892
rect 28040 32852 28046 32864
rect 28077 32861 28089 32864
rect 28123 32861 28135 32895
rect 28077 32855 28135 32861
rect 28169 32895 28227 32901
rect 28169 32861 28181 32895
rect 28215 32892 28227 32895
rect 28368 32892 28396 32932
rect 29638 32920 29644 32932
rect 29696 32960 29702 32972
rect 29696 32932 29776 32960
rect 29696 32920 29702 32932
rect 28215 32864 28396 32892
rect 28215 32861 28227 32864
rect 28169 32855 28227 32861
rect 28442 32852 28448 32904
rect 28500 32892 28506 32904
rect 29748 32901 29776 32932
rect 30834 32920 30840 32972
rect 30892 32960 30898 32972
rect 31021 32963 31079 32969
rect 31021 32960 31033 32963
rect 30892 32932 31033 32960
rect 30892 32920 30898 32932
rect 31021 32929 31033 32932
rect 31067 32929 31079 32963
rect 31021 32923 31079 32929
rect 31205 32963 31263 32969
rect 31205 32929 31217 32963
rect 31251 32960 31263 32963
rect 36357 32963 36415 32969
rect 36357 32960 36369 32963
rect 31251 32932 36369 32960
rect 31251 32929 31263 32932
rect 31205 32923 31263 32929
rect 29733 32895 29791 32901
rect 28500 32864 28545 32892
rect 28500 32852 28506 32864
rect 29733 32861 29745 32895
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29822 32852 29828 32904
rect 29880 32892 29886 32904
rect 29917 32895 29975 32901
rect 29917 32892 29929 32895
rect 29880 32864 29929 32892
rect 29880 32852 29886 32864
rect 29917 32861 29929 32864
rect 29963 32861 29975 32895
rect 29917 32855 29975 32861
rect 30006 32852 30012 32904
rect 30064 32892 30070 32904
rect 30929 32895 30987 32901
rect 30929 32892 30941 32895
rect 30064 32864 30941 32892
rect 30064 32852 30070 32864
rect 30929 32861 30941 32864
rect 30975 32892 30987 32895
rect 31662 32892 31668 32904
rect 30975 32864 31668 32892
rect 30975 32861 30987 32864
rect 30929 32855 30987 32861
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 31754 32852 31760 32904
rect 31812 32892 31818 32904
rect 32692 32901 32720 32932
rect 36357 32929 36369 32932
rect 36403 32960 36415 32963
rect 36538 32960 36544 32972
rect 36403 32932 36544 32960
rect 36403 32929 36415 32932
rect 36357 32923 36415 32929
rect 36538 32920 36544 32932
rect 36596 32920 36602 32972
rect 32677 32895 32735 32901
rect 31812 32864 31857 32892
rect 31812 32852 31818 32864
rect 32677 32861 32689 32895
rect 32723 32861 32735 32895
rect 32677 32855 32735 32861
rect 32766 32852 32772 32904
rect 32824 32892 32830 32904
rect 33597 32895 33655 32901
rect 33597 32892 33609 32895
rect 32824 32864 33609 32892
rect 32824 32852 32830 32864
rect 33597 32861 33609 32864
rect 33643 32861 33655 32895
rect 33597 32855 33655 32861
rect 36081 32895 36139 32901
rect 36081 32861 36093 32895
rect 36127 32892 36139 32895
rect 36170 32892 36176 32904
rect 36127 32864 36176 32892
rect 36127 32861 36139 32864
rect 36081 32855 36139 32861
rect 36170 32852 36176 32864
rect 36228 32852 36234 32904
rect 46290 32892 46296 32904
rect 46251 32864 46296 32892
rect 46290 32852 46296 32864
rect 46348 32852 46354 32904
rect 19150 32784 19156 32836
rect 19208 32824 19214 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 19208 32796 19441 32824
rect 19208 32784 19214 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 21082 32824 21088 32836
rect 21043 32796 21088 32824
rect 19429 32787 19487 32793
rect 21082 32784 21088 32796
rect 21140 32784 21146 32836
rect 24946 32784 24952 32836
rect 25004 32824 25010 32836
rect 40034 32824 40040 32836
rect 25004 32796 40040 32824
rect 25004 32784 25010 32796
rect 40034 32784 40040 32796
rect 40092 32784 40098 32836
rect 46477 32827 46535 32833
rect 46477 32793 46489 32827
rect 46523 32824 46535 32827
rect 47670 32824 47676 32836
rect 46523 32796 47676 32824
rect 46523 32793 46535 32796
rect 46477 32787 46535 32793
rect 47670 32784 47676 32796
rect 47728 32784 47734 32836
rect 48130 32824 48136 32836
rect 48091 32796 48136 32824
rect 48130 32784 48136 32796
rect 48188 32784 48194 32836
rect 17828 32728 18828 32756
rect 22005 32759 22063 32765
rect 17828 32716 17834 32728
rect 22005 32725 22017 32759
rect 22051 32756 22063 32759
rect 22278 32756 22284 32768
rect 22051 32728 22284 32756
rect 22051 32725 22063 32728
rect 22005 32719 22063 32725
rect 22278 32716 22284 32728
rect 22336 32716 22342 32768
rect 22738 32716 22744 32768
rect 22796 32756 22802 32768
rect 23017 32759 23075 32765
rect 23017 32756 23029 32759
rect 22796 32728 23029 32756
rect 22796 32716 22802 32728
rect 23017 32725 23029 32728
rect 23063 32725 23075 32759
rect 23017 32719 23075 32725
rect 23753 32759 23811 32765
rect 23753 32725 23765 32759
rect 23799 32756 23811 32759
rect 28442 32756 28448 32768
rect 23799 32728 28448 32756
rect 23799 32725 23811 32728
rect 23753 32719 23811 32725
rect 28442 32716 28448 32728
rect 28500 32716 28506 32768
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 29549 32759 29607 32765
rect 29549 32756 29561 32759
rect 28868 32728 29561 32756
rect 28868 32716 28874 32728
rect 29549 32725 29561 32728
rect 29595 32725 29607 32759
rect 29549 32719 29607 32725
rect 32030 32716 32036 32768
rect 32088 32756 32094 32768
rect 32861 32759 32919 32765
rect 32861 32756 32873 32759
rect 32088 32728 32873 32756
rect 32088 32716 32094 32728
rect 32861 32725 32873 32728
rect 32907 32725 32919 32759
rect 33410 32756 33416 32768
rect 33371 32728 33416 32756
rect 32861 32719 32919 32725
rect 33410 32716 33416 32728
rect 33468 32716 33474 32768
rect 36170 32716 36176 32768
rect 36228 32756 36234 32768
rect 36228 32728 36273 32756
rect 36228 32716 36234 32728
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 22373 32555 22431 32561
rect 22373 32521 22385 32555
rect 22419 32552 22431 32555
rect 22462 32552 22468 32564
rect 22419 32524 22468 32552
rect 22419 32521 22431 32524
rect 22373 32515 22431 32521
rect 22462 32512 22468 32524
rect 22520 32512 22526 32564
rect 24857 32555 24915 32561
rect 24857 32521 24869 32555
rect 24903 32552 24915 32555
rect 25038 32552 25044 32564
rect 24903 32524 25044 32552
rect 24903 32521 24915 32524
rect 24857 32515 24915 32521
rect 25038 32512 25044 32524
rect 25096 32512 25102 32564
rect 27890 32512 27896 32564
rect 27948 32552 27954 32564
rect 28997 32555 29055 32561
rect 28997 32552 29009 32555
rect 27948 32524 29009 32552
rect 27948 32512 27954 32524
rect 28997 32521 29009 32524
rect 29043 32521 29055 32555
rect 31938 32552 31944 32564
rect 28997 32515 29055 32521
rect 31726 32524 31944 32552
rect 2314 32484 2320 32496
rect 2275 32456 2320 32484
rect 2314 32444 2320 32456
rect 2372 32444 2378 32496
rect 12710 32484 12716 32496
rect 11716 32456 12716 32484
rect 11716 32425 11744 32456
rect 12710 32444 12716 32456
rect 12768 32484 12774 32496
rect 19334 32484 19340 32496
rect 12768 32456 14688 32484
rect 19295 32456 19340 32484
rect 12768 32444 12774 32456
rect 11701 32419 11759 32425
rect 11701 32385 11713 32419
rect 11747 32385 11759 32419
rect 11701 32379 11759 32385
rect 12805 32419 12863 32425
rect 12805 32385 12817 32419
rect 12851 32416 12863 32419
rect 14550 32416 14556 32428
rect 12851 32388 14556 32416
rect 12851 32385 12863 32388
rect 12805 32379 12863 32385
rect 14550 32376 14556 32388
rect 14608 32376 14614 32428
rect 14660 32425 14688 32456
rect 19334 32444 19340 32456
rect 19392 32444 19398 32496
rect 20993 32487 21051 32493
rect 20993 32453 21005 32487
rect 21039 32484 21051 32487
rect 31726 32484 31754 32524
rect 31938 32512 31944 32524
rect 31996 32512 32002 32564
rect 33410 32552 33416 32564
rect 32508 32524 33416 32552
rect 32508 32493 32536 32524
rect 33410 32512 33416 32524
rect 33468 32512 33474 32564
rect 35713 32555 35771 32561
rect 35713 32521 35725 32555
rect 35759 32552 35771 32555
rect 36170 32552 36176 32564
rect 35759 32524 36176 32552
rect 35759 32521 35771 32524
rect 35713 32515 35771 32521
rect 36170 32512 36176 32524
rect 36228 32512 36234 32564
rect 46845 32555 46903 32561
rect 46845 32552 46857 32555
rect 45526 32524 46857 32552
rect 21039 32456 31754 32484
rect 32493 32487 32551 32493
rect 21039 32453 21051 32456
rect 20993 32447 21051 32453
rect 32493 32453 32505 32487
rect 32539 32453 32551 32487
rect 34054 32484 34060 32496
rect 33718 32456 34060 32484
rect 32493 32447 32551 32453
rect 34054 32444 34060 32456
rect 34112 32444 34118 32496
rect 34793 32487 34851 32493
rect 34793 32453 34805 32487
rect 34839 32484 34851 32487
rect 45526 32484 45554 32524
rect 46845 32521 46857 32524
rect 46891 32521 46903 32555
rect 47670 32552 47676 32564
rect 47631 32524 47676 32552
rect 46845 32515 46903 32521
rect 47670 32512 47676 32524
rect 47728 32512 47734 32564
rect 34839 32456 45554 32484
rect 34839 32453 34851 32456
rect 34793 32447 34851 32453
rect 46658 32444 46664 32496
rect 46716 32484 46722 32496
rect 46716 32456 47256 32484
rect 46716 32444 46722 32456
rect 47228 32428 47256 32456
rect 14645 32419 14703 32425
rect 14645 32385 14657 32419
rect 14691 32385 14703 32419
rect 15654 32416 15660 32428
rect 15615 32388 15660 32416
rect 14645 32379 14703 32385
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 16390 32376 16396 32428
rect 16448 32416 16454 32428
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 16448 32388 16681 32416
rect 16448 32376 16454 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 22005 32419 22063 32425
rect 22005 32385 22017 32419
rect 22051 32416 22063 32419
rect 22278 32416 22284 32428
rect 22051 32388 22284 32416
rect 22051 32385 22063 32388
rect 22005 32379 22063 32385
rect 22278 32376 22284 32388
rect 22336 32416 22342 32428
rect 22554 32416 22560 32428
rect 22336 32388 22560 32416
rect 22336 32376 22342 32388
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 24210 32376 24216 32428
rect 24268 32416 24274 32428
rect 24489 32419 24547 32425
rect 24489 32416 24501 32419
rect 24268 32388 24501 32416
rect 24268 32376 24274 32388
rect 24489 32385 24501 32388
rect 24535 32416 24547 32419
rect 24762 32416 24768 32428
rect 24535 32388 24768 32416
rect 24535 32385 24547 32388
rect 24489 32379 24547 32385
rect 24762 32376 24768 32388
rect 24820 32376 24826 32428
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 28445 32419 28503 32425
rect 28445 32385 28457 32419
rect 28491 32416 28503 32419
rect 28626 32416 28632 32428
rect 28491 32388 28632 32416
rect 28491 32385 28503 32388
rect 28445 32379 28503 32385
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 28813 32419 28871 32425
rect 28813 32385 28825 32419
rect 28859 32416 28871 32419
rect 29730 32416 29736 32428
rect 28859 32388 29736 32416
rect 28859 32385 28871 32388
rect 28813 32379 28871 32385
rect 29730 32376 29736 32388
rect 29788 32376 29794 32428
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32416 29975 32419
rect 30006 32416 30012 32428
rect 29963 32388 30012 32416
rect 29963 32385 29975 32388
rect 29917 32379 29975 32385
rect 30006 32376 30012 32388
rect 30064 32376 30070 32428
rect 30101 32419 30159 32425
rect 30101 32385 30113 32419
rect 30147 32385 30159 32419
rect 32214 32416 32220 32428
rect 32175 32388 32220 32416
rect 30101 32379 30159 32385
rect 2133 32351 2191 32357
rect 2133 32317 2145 32351
rect 2179 32348 2191 32351
rect 2406 32348 2412 32360
rect 2179 32320 2412 32348
rect 2179 32317 2191 32320
rect 2133 32311 2191 32317
rect 2406 32308 2412 32320
rect 2464 32308 2470 32360
rect 3234 32348 3240 32360
rect 3195 32320 3240 32348
rect 3234 32308 3240 32320
rect 3292 32308 3298 32360
rect 12618 32308 12624 32360
rect 12676 32348 12682 32360
rect 12897 32351 12955 32357
rect 12897 32348 12909 32351
rect 12676 32320 12909 32348
rect 12676 32308 12682 32320
rect 12897 32317 12909 32320
rect 12943 32348 12955 32351
rect 14458 32348 14464 32360
rect 12943 32320 14464 32348
rect 12943 32317 12955 32320
rect 12897 32311 12955 32317
rect 14458 32308 14464 32320
rect 14516 32308 14522 32360
rect 17586 32308 17592 32360
rect 17644 32348 17650 32360
rect 19153 32351 19211 32357
rect 19153 32348 19165 32351
rect 17644 32320 19165 32348
rect 17644 32308 17650 32320
rect 19153 32317 19165 32320
rect 19199 32317 19211 32351
rect 19153 32311 19211 32317
rect 21913 32351 21971 32357
rect 21913 32317 21925 32351
rect 21959 32348 21971 32351
rect 22462 32348 22468 32360
rect 21959 32320 22468 32348
rect 21959 32317 21971 32320
rect 21913 32311 21971 32317
rect 22462 32308 22468 32320
rect 22520 32308 22526 32360
rect 24581 32351 24639 32357
rect 24581 32317 24593 32351
rect 24627 32348 24639 32351
rect 25130 32348 25136 32360
rect 24627 32320 25136 32348
rect 24627 32317 24639 32320
rect 24581 32311 24639 32317
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 25240 32320 28396 32348
rect 14182 32240 14188 32292
rect 14240 32280 14246 32292
rect 17770 32280 17776 32292
rect 14240 32252 17776 32280
rect 14240 32240 14246 32252
rect 17770 32240 17776 32252
rect 17828 32240 17834 32292
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1673 32215 1731 32221
rect 1673 32212 1685 32215
rect 1452 32184 1685 32212
rect 1452 32172 1458 32184
rect 1673 32181 1685 32184
rect 1719 32181 1731 32215
rect 11698 32212 11704 32224
rect 11659 32184 11704 32212
rect 1673 32175 1731 32181
rect 11698 32172 11704 32184
rect 11756 32172 11762 32224
rect 13170 32212 13176 32224
rect 13131 32184 13176 32212
rect 13170 32172 13176 32184
rect 13228 32172 13234 32224
rect 14737 32215 14795 32221
rect 14737 32181 14749 32215
rect 14783 32212 14795 32215
rect 15194 32212 15200 32224
rect 14783 32184 15200 32212
rect 14783 32181 14795 32184
rect 14737 32175 14795 32181
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 15470 32212 15476 32224
rect 15431 32184 15476 32212
rect 15470 32172 15476 32184
rect 15528 32172 15534 32224
rect 16758 32212 16764 32224
rect 16719 32184 16764 32212
rect 16758 32172 16764 32184
rect 16816 32172 16822 32224
rect 23474 32172 23480 32224
rect 23532 32212 23538 32224
rect 24670 32212 24676 32224
rect 23532 32184 24676 32212
rect 23532 32172 23538 32184
rect 24670 32172 24676 32184
rect 24728 32212 24734 32224
rect 25240 32212 25268 32320
rect 28368 32280 28396 32320
rect 29638 32308 29644 32360
rect 29696 32348 29702 32360
rect 30116 32348 30144 32379
rect 32214 32376 32220 32388
rect 32272 32376 32278 32428
rect 34440 32388 35020 32416
rect 29696 32320 30144 32348
rect 29696 32308 29702 32320
rect 32122 32308 32128 32360
rect 32180 32348 32186 32360
rect 34440 32348 34468 32388
rect 32180 32320 34468 32348
rect 32180 32308 32186 32320
rect 34514 32308 34520 32360
rect 34572 32348 34578 32360
rect 34992 32357 35020 32388
rect 35066 32376 35072 32428
rect 35124 32416 35130 32428
rect 36081 32419 36139 32425
rect 36081 32416 36093 32419
rect 35124 32388 36093 32416
rect 35124 32376 35130 32388
rect 36081 32385 36093 32388
rect 36127 32385 36139 32419
rect 37458 32416 37464 32428
rect 37419 32388 37464 32416
rect 36081 32379 36139 32385
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 46842 32376 46848 32428
rect 46900 32416 46906 32428
rect 47029 32419 47087 32425
rect 47029 32416 47041 32419
rect 46900 32388 47041 32416
rect 46900 32376 46906 32388
rect 47029 32385 47041 32388
rect 47075 32385 47087 32419
rect 47029 32379 47087 32385
rect 47210 32376 47216 32428
rect 47268 32416 47274 32428
rect 47581 32419 47639 32425
rect 47581 32416 47593 32419
rect 47268 32388 47593 32416
rect 47268 32376 47274 32388
rect 47581 32385 47593 32388
rect 47627 32385 47639 32419
rect 47581 32379 47639 32385
rect 34885 32351 34943 32357
rect 34885 32348 34897 32351
rect 34572 32320 34897 32348
rect 34572 32308 34578 32320
rect 34885 32317 34897 32320
rect 34931 32317 34943 32351
rect 34885 32311 34943 32317
rect 34977 32351 35035 32357
rect 34977 32317 34989 32351
rect 35023 32348 35035 32351
rect 36170 32348 36176 32360
rect 35023 32320 35894 32348
rect 36131 32320 36176 32348
rect 35023 32317 35035 32320
rect 34977 32311 35035 32317
rect 32030 32280 32036 32292
rect 28368 32252 32036 32280
rect 32030 32240 32036 32252
rect 32088 32240 32094 32292
rect 34425 32283 34483 32289
rect 34425 32280 34437 32283
rect 33520 32252 34437 32280
rect 24728 32184 25268 32212
rect 25501 32215 25559 32221
rect 24728 32172 24734 32184
rect 25501 32181 25513 32215
rect 25547 32212 25559 32215
rect 26326 32212 26332 32224
rect 25547 32184 26332 32212
rect 25547 32181 25559 32184
rect 25501 32175 25559 32181
rect 26326 32172 26332 32184
rect 26384 32172 26390 32224
rect 28810 32212 28816 32224
rect 28771 32184 28816 32212
rect 28810 32172 28816 32184
rect 28868 32172 28874 32224
rect 29914 32172 29920 32224
rect 29972 32212 29978 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 29972 32184 30297 32212
rect 29972 32172 29978 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 30285 32175 30343 32181
rect 33226 32172 33232 32224
rect 33284 32212 33290 32224
rect 33520 32212 33548 32252
rect 34425 32249 34437 32252
rect 34471 32249 34483 32283
rect 35866 32280 35894 32320
rect 36170 32308 36176 32320
rect 36228 32308 36234 32360
rect 36354 32348 36360 32360
rect 36315 32320 36360 32348
rect 36354 32308 36360 32320
rect 36412 32308 36418 32360
rect 36372 32280 36400 32308
rect 35866 32252 36400 32280
rect 34425 32243 34483 32249
rect 33284 32184 33548 32212
rect 33284 32172 33290 32184
rect 33870 32172 33876 32224
rect 33928 32212 33934 32224
rect 33965 32215 34023 32221
rect 33965 32212 33977 32215
rect 33928 32184 33977 32212
rect 33928 32172 33934 32184
rect 33965 32181 33977 32184
rect 34011 32181 34023 32215
rect 33965 32175 34023 32181
rect 36078 32172 36084 32224
rect 36136 32212 36142 32224
rect 37277 32215 37335 32221
rect 37277 32212 37289 32215
rect 36136 32184 37289 32212
rect 36136 32172 36142 32184
rect 37277 32181 37289 32184
rect 37323 32181 37335 32215
rect 37277 32175 37335 32181
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 14277 32011 14335 32017
rect 14277 31977 14289 32011
rect 14323 31977 14335 32011
rect 14458 32008 14464 32020
rect 14419 31980 14464 32008
rect 14277 31971 14335 31977
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 11698 31872 11704 31884
rect 11659 31844 11704 31872
rect 11698 31832 11704 31844
rect 11756 31832 11762 31884
rect 11974 31872 11980 31884
rect 11935 31844 11980 31872
rect 11974 31832 11980 31844
rect 12032 31832 12038 31884
rect 12618 31832 12624 31884
rect 12676 31872 12682 31884
rect 14292 31872 14320 31971
rect 14458 31968 14464 31980
rect 14516 31968 14522 32020
rect 14550 31968 14556 32020
rect 14608 32008 14614 32020
rect 16850 32008 16856 32020
rect 14608 31980 16856 32008
rect 14608 31968 14614 31980
rect 16850 31968 16856 31980
rect 16908 32008 16914 32020
rect 17678 32008 17684 32020
rect 16908 31980 17684 32008
rect 16908 31968 16914 31980
rect 17678 31968 17684 31980
rect 17736 31968 17742 32020
rect 21542 31968 21548 32020
rect 21600 32008 21606 32020
rect 21637 32011 21695 32017
rect 21637 32008 21649 32011
rect 21600 31980 21649 32008
rect 21600 31968 21606 31980
rect 21637 31977 21649 31980
rect 21683 31977 21695 32011
rect 32766 32008 32772 32020
rect 32727 31980 32772 32008
rect 21637 31971 21695 31977
rect 32766 31968 32772 31980
rect 32824 31968 32830 32020
rect 34054 32008 34060 32020
rect 34015 31980 34060 32008
rect 34054 31968 34060 31980
rect 34112 31968 34118 32020
rect 36262 31968 36268 32020
rect 36320 32008 36326 32020
rect 37553 32011 37611 32017
rect 37553 32008 37565 32011
rect 36320 31980 37565 32008
rect 36320 31968 36326 31980
rect 37553 31977 37565 31980
rect 37599 31977 37611 32011
rect 37553 31971 37611 31977
rect 46290 31968 46296 32020
rect 46348 32008 46354 32020
rect 47673 32011 47731 32017
rect 47673 32008 47685 32011
rect 46348 31980 47685 32008
rect 46348 31968 46354 31980
rect 47673 31977 47685 31980
rect 47719 31977 47731 32011
rect 47673 31971 47731 31977
rect 18156 31912 19748 31940
rect 14366 31872 14372 31884
rect 12676 31844 14372 31872
rect 12676 31832 12682 31844
rect 14366 31832 14372 31844
rect 14424 31832 14430 31884
rect 15194 31872 15200 31884
rect 15155 31844 15200 31872
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 15470 31872 15476 31884
rect 15431 31844 15476 31872
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 16666 31832 16672 31884
rect 16724 31872 16730 31884
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 16724 31844 16957 31872
rect 16724 31832 16730 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 14182 31806 14188 31816
rect 14108 31804 14188 31806
rect 13464 31778 14188 31804
rect 13464 31776 14136 31778
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 9306 31696 9312 31748
rect 9364 31736 9370 31748
rect 10778 31736 10784 31748
rect 9364 31708 10784 31736
rect 9364 31696 9370 31708
rect 10778 31696 10784 31708
rect 10836 31696 10842 31748
rect 12434 31696 12440 31748
rect 12492 31696 12498 31748
rect 3970 31628 3976 31680
rect 4028 31668 4034 31680
rect 12802 31668 12808 31680
rect 4028 31640 12808 31668
rect 4028 31628 4034 31640
rect 12802 31628 12808 31640
rect 12860 31628 12866 31680
rect 12894 31628 12900 31680
rect 12952 31668 12958 31680
rect 13464 31677 13492 31776
rect 14108 31745 14136 31776
rect 14182 31764 14188 31778
rect 14240 31764 14246 31816
rect 16758 31804 16764 31816
rect 16606 31776 16764 31804
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 16960 31804 16988 31835
rect 17310 31832 17316 31884
rect 17368 31872 17374 31884
rect 18049 31875 18107 31881
rect 18049 31872 18061 31875
rect 17368 31844 18061 31872
rect 17368 31832 17374 31844
rect 18049 31841 18061 31844
rect 18095 31841 18107 31875
rect 18049 31835 18107 31841
rect 17586 31804 17592 31816
rect 16960 31776 17592 31804
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 17678 31764 17684 31816
rect 17736 31804 17742 31816
rect 17736 31776 17781 31804
rect 17736 31764 17742 31776
rect 18156 31748 18184 31912
rect 19720 31881 19748 31912
rect 32214 31900 32220 31952
rect 32272 31940 32278 31952
rect 32272 31912 35848 31940
rect 32272 31900 32278 31912
rect 18601 31875 18659 31881
rect 18601 31841 18613 31875
rect 18647 31872 18659 31875
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 18647 31844 19441 31872
rect 18647 31841 18659 31844
rect 18601 31835 18659 31841
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 19429 31835 19487 31841
rect 19705 31875 19763 31881
rect 19705 31841 19717 31875
rect 19751 31841 19763 31875
rect 19705 31835 19763 31841
rect 20990 31832 20996 31884
rect 21048 31872 21054 31884
rect 27246 31872 27252 31884
rect 21048 31844 21588 31872
rect 27207 31844 27252 31872
rect 21048 31832 21054 31844
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18555 31776 19104 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 14093 31739 14151 31745
rect 14093 31705 14105 31739
rect 14139 31736 14151 31739
rect 14309 31739 14367 31745
rect 14139 31708 14171 31736
rect 14139 31705 14151 31708
rect 14093 31699 14151 31705
rect 14309 31705 14321 31739
rect 14355 31736 14367 31739
rect 14642 31736 14648 31748
rect 14355 31708 14648 31736
rect 14355 31705 14367 31708
rect 14309 31699 14367 31705
rect 14642 31696 14648 31708
rect 14700 31696 14706 31748
rect 17034 31736 17040 31748
rect 16868 31708 17040 31736
rect 13449 31671 13507 31677
rect 13449 31668 13461 31671
rect 12952 31640 13461 31668
rect 12952 31628 12958 31640
rect 13449 31637 13461 31640
rect 13495 31637 13507 31671
rect 13449 31631 13507 31637
rect 14458 31628 14464 31680
rect 14516 31668 14522 31680
rect 16868 31668 16896 31708
rect 17034 31696 17040 31708
rect 17092 31736 17098 31748
rect 17957 31739 18015 31745
rect 17957 31736 17969 31739
rect 17092 31708 17969 31736
rect 17092 31696 17098 31708
rect 17957 31705 17969 31708
rect 18003 31705 18015 31739
rect 17957 31699 18015 31705
rect 18138 31696 18144 31748
rect 18196 31696 18202 31748
rect 19076 31736 19104 31776
rect 19150 31764 19156 31816
rect 19208 31804 19214 31816
rect 21560 31813 21588 31844
rect 27246 31832 27252 31844
rect 27304 31832 27310 31884
rect 27525 31875 27583 31881
rect 27525 31841 27537 31875
rect 27571 31872 27583 31875
rect 28534 31872 28540 31884
rect 27571 31844 28540 31872
rect 27571 31841 27583 31844
rect 27525 31835 27583 31841
rect 28534 31832 28540 31844
rect 28592 31832 28598 31884
rect 32030 31832 32036 31884
rect 32088 31872 32094 31884
rect 32490 31872 32496 31884
rect 32088 31844 32496 31872
rect 32088 31832 32094 31844
rect 32490 31832 32496 31844
rect 32548 31872 32554 31884
rect 35820 31881 35848 31912
rect 33321 31875 33379 31881
rect 33321 31872 33333 31875
rect 32548 31844 33333 31872
rect 32548 31832 32554 31844
rect 33321 31841 33333 31844
rect 33367 31841 33379 31875
rect 33321 31835 33379 31841
rect 35805 31875 35863 31881
rect 35805 31841 35817 31875
rect 35851 31841 35863 31875
rect 36078 31872 36084 31884
rect 36039 31844 36084 31872
rect 35805 31835 35863 31841
rect 36078 31832 36084 31844
rect 36136 31832 36142 31884
rect 19245 31807 19303 31813
rect 19245 31804 19257 31807
rect 19208 31776 19257 31804
rect 19208 31764 19214 31776
rect 19245 31773 19257 31776
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 21545 31807 21603 31813
rect 21545 31773 21557 31807
rect 21591 31773 21603 31807
rect 21545 31767 21603 31773
rect 25593 31807 25651 31813
rect 25593 31773 25605 31807
rect 25639 31804 25651 31807
rect 26326 31804 26332 31816
rect 25639 31776 26332 31804
rect 25639 31773 25651 31776
rect 25593 31767 25651 31773
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 19426 31736 19432 31748
rect 19076 31708 19432 31736
rect 19426 31696 19432 31708
rect 19484 31696 19490 31748
rect 26234 31696 26240 31748
rect 26292 31736 26298 31748
rect 27264 31736 27292 31832
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 33962 31804 33968 31816
rect 31812 31776 33364 31804
rect 33923 31776 33968 31804
rect 31812 31764 31818 31776
rect 33336 31748 33364 31776
rect 33962 31764 33968 31776
rect 34020 31764 34026 31816
rect 26292 31708 27292 31736
rect 26292 31696 26298 31708
rect 27982 31696 27988 31748
rect 28040 31696 28046 31748
rect 33226 31736 33232 31748
rect 33187 31708 33232 31736
rect 33226 31696 33232 31708
rect 33284 31696 33290 31748
rect 33318 31696 33324 31748
rect 33376 31696 33382 31748
rect 37366 31736 37372 31748
rect 37306 31708 37372 31736
rect 37366 31696 37372 31708
rect 37424 31696 37430 31748
rect 14516 31640 16896 31668
rect 14516 31628 14522 31640
rect 16942 31628 16948 31680
rect 17000 31668 17006 31680
rect 17405 31671 17463 31677
rect 17405 31668 17417 31671
rect 17000 31640 17417 31668
rect 17000 31628 17006 31640
rect 17405 31637 17417 31640
rect 17451 31637 17463 31671
rect 17770 31668 17776 31680
rect 17731 31640 17776 31668
rect 17405 31631 17463 31637
rect 17770 31628 17776 31640
rect 17828 31628 17834 31680
rect 25590 31628 25596 31680
rect 25648 31668 25654 31680
rect 25685 31671 25743 31677
rect 25685 31668 25697 31671
rect 25648 31640 25697 31668
rect 25648 31628 25654 31640
rect 25685 31637 25697 31640
rect 25731 31637 25743 31671
rect 25685 31631 25743 31637
rect 28997 31671 29055 31677
rect 28997 31637 29009 31671
rect 29043 31668 29055 31671
rect 29178 31668 29184 31680
rect 29043 31640 29184 31668
rect 29043 31637 29055 31640
rect 28997 31631 29055 31637
rect 29178 31628 29184 31640
rect 29236 31628 29242 31680
rect 31018 31628 31024 31680
rect 31076 31668 31082 31680
rect 33137 31671 33195 31677
rect 33137 31668 33149 31671
rect 31076 31640 33149 31668
rect 31076 31628 31082 31640
rect 33137 31637 33149 31640
rect 33183 31668 33195 31671
rect 33594 31668 33600 31680
rect 33183 31640 33600 31668
rect 33183 31637 33195 31640
rect 33137 31631 33195 31637
rect 33594 31628 33600 31640
rect 33652 31668 33658 31680
rect 33870 31668 33876 31680
rect 33652 31640 33876 31668
rect 33652 31628 33658 31640
rect 33870 31628 33876 31640
rect 33928 31628 33934 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 1636 31436 2237 31464
rect 1636 31424 1642 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 9398 31464 9404 31476
rect 2225 31427 2283 31433
rect 9140 31436 9404 31464
rect 2133 31331 2191 31337
rect 2133 31297 2145 31331
rect 2179 31328 2191 31331
rect 2222 31328 2228 31340
rect 2179 31300 2228 31328
rect 2179 31297 2191 31300
rect 2133 31291 2191 31297
rect 2222 31288 2228 31300
rect 2280 31328 2286 31340
rect 7190 31328 7196 31340
rect 2280 31300 7196 31328
rect 2280 31288 2286 31300
rect 7190 31288 7196 31300
rect 7248 31288 7254 31340
rect 9140 31337 9168 31436
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 11609 31467 11667 31473
rect 11609 31433 11621 31467
rect 11655 31464 11667 31467
rect 12250 31464 12256 31476
rect 11655 31436 12256 31464
rect 11655 31433 11667 31436
rect 11609 31427 11667 31433
rect 12250 31424 12256 31436
rect 12308 31424 12314 31476
rect 12345 31467 12403 31473
rect 12345 31433 12357 31467
rect 12391 31464 12403 31467
rect 12618 31464 12624 31476
rect 12391 31436 12624 31464
rect 12391 31433 12403 31436
rect 12345 31427 12403 31433
rect 12618 31424 12624 31436
rect 12676 31424 12682 31476
rect 12802 31424 12808 31476
rect 12860 31464 12866 31476
rect 12860 31436 14504 31464
rect 12860 31424 12866 31436
rect 12161 31399 12219 31405
rect 9324 31368 11652 31396
rect 9125 31331 9183 31337
rect 9125 31297 9137 31331
rect 9171 31297 9183 31331
rect 9324 31328 9352 31368
rect 9125 31291 9183 31297
rect 9232 31300 9352 31328
rect 10045 31331 10103 31337
rect 8754 31220 8760 31272
rect 8812 31260 8818 31272
rect 9232 31269 9260 31300
rect 10045 31297 10057 31331
rect 10091 31328 10103 31331
rect 10689 31331 10747 31337
rect 10091 31300 10548 31328
rect 10091 31297 10103 31300
rect 10045 31291 10103 31297
rect 9217 31263 9275 31269
rect 9217 31260 9229 31263
rect 8812 31232 9229 31260
rect 8812 31220 8818 31232
rect 9217 31229 9229 31232
rect 9263 31229 9275 31263
rect 9217 31223 9275 31229
rect 10520 31192 10548 31300
rect 10689 31297 10701 31331
rect 10735 31328 10747 31331
rect 11514 31328 11520 31340
rect 10735 31300 11520 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 11624 31328 11652 31368
rect 12161 31365 12173 31399
rect 12207 31396 12219 31399
rect 12894 31396 12900 31408
rect 12207 31368 12900 31396
rect 12207 31365 12219 31368
rect 12161 31359 12219 31365
rect 12894 31356 12900 31368
rect 12952 31356 12958 31408
rect 13170 31396 13176 31408
rect 13131 31368 13176 31396
rect 13170 31356 13176 31368
rect 13228 31356 13234 31408
rect 14182 31356 14188 31408
rect 14240 31356 14246 31408
rect 14476 31396 14504 31436
rect 14550 31424 14556 31476
rect 14608 31464 14614 31476
rect 14645 31467 14703 31473
rect 14645 31464 14657 31467
rect 14608 31436 14657 31464
rect 14608 31424 14614 31436
rect 14645 31433 14657 31436
rect 14691 31433 14703 31467
rect 14645 31427 14703 31433
rect 15654 31424 15660 31476
rect 15712 31464 15718 31476
rect 15749 31467 15807 31473
rect 15749 31464 15761 31467
rect 15712 31436 15761 31464
rect 15712 31424 15718 31436
rect 15749 31433 15761 31436
rect 15795 31433 15807 31467
rect 16945 31467 17003 31473
rect 15749 31427 15807 31433
rect 15856 31436 16896 31464
rect 15856 31396 15884 31436
rect 16666 31396 16672 31408
rect 14476 31368 15884 31396
rect 16627 31368 16672 31396
rect 16666 31356 16672 31368
rect 16724 31356 16730 31408
rect 16868 31396 16896 31436
rect 16945 31433 16957 31467
rect 16991 31464 17003 31467
rect 17770 31464 17776 31476
rect 16991 31436 17776 31464
rect 16991 31433 17003 31436
rect 16945 31427 17003 31433
rect 17770 31424 17776 31436
rect 17828 31424 17834 31476
rect 23934 31424 23940 31476
rect 23992 31464 23998 31476
rect 26234 31464 26240 31476
rect 23992 31436 26240 31464
rect 23992 31424 23998 31436
rect 18138 31396 18144 31408
rect 16868 31368 18144 31396
rect 18138 31356 18144 31368
rect 18196 31356 18202 31408
rect 24688 31396 24716 31436
rect 26234 31424 26240 31436
rect 26292 31424 26298 31476
rect 27341 31467 27399 31473
rect 27341 31433 27353 31467
rect 27387 31464 27399 31467
rect 27982 31464 27988 31476
rect 27387 31436 27988 31464
rect 27387 31433 27399 31436
rect 27341 31427 27399 31433
rect 27982 31424 27988 31436
rect 28040 31424 28046 31476
rect 28534 31424 28540 31476
rect 28592 31464 28598 31476
rect 28629 31467 28687 31473
rect 28629 31464 28641 31467
rect 28592 31436 28641 31464
rect 28592 31424 28598 31436
rect 28629 31433 28641 31436
rect 28675 31433 28687 31467
rect 28629 31427 28687 31433
rect 36170 31424 36176 31476
rect 36228 31464 36234 31476
rect 36633 31467 36691 31473
rect 36633 31464 36645 31467
rect 36228 31436 36645 31464
rect 36228 31424 36234 31436
rect 36633 31433 36645 31436
rect 36679 31433 36691 31467
rect 37366 31464 37372 31476
rect 37327 31436 37372 31464
rect 36633 31427 36691 31433
rect 37366 31424 37372 31436
rect 37424 31424 37430 31476
rect 24596 31368 24716 31396
rect 12437 31331 12495 31337
rect 12437 31328 12449 31331
rect 11624 31300 12449 31328
rect 12437 31297 12449 31300
rect 12483 31328 12495 31331
rect 12802 31328 12808 31340
rect 12483 31300 12808 31328
rect 12483 31297 12495 31300
rect 12437 31291 12495 31297
rect 12802 31288 12808 31300
rect 12860 31288 12866 31340
rect 15565 31331 15623 31337
rect 15565 31297 15577 31331
rect 15611 31328 15623 31331
rect 16758 31328 16764 31340
rect 15611 31300 16764 31328
rect 15611 31297 15623 31300
rect 15565 31291 15623 31297
rect 16758 31288 16764 31300
rect 16816 31288 16822 31340
rect 16850 31288 16856 31340
rect 16908 31328 16914 31340
rect 16908 31300 16953 31328
rect 16908 31288 16914 31300
rect 17034 31288 17040 31340
rect 17092 31328 17098 31340
rect 17092 31300 17137 31328
rect 17092 31288 17098 31300
rect 19242 31288 19248 31340
rect 19300 31288 19306 31340
rect 22278 31328 22284 31340
rect 22239 31300 22284 31328
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22462 31328 22468 31340
rect 22423 31300 22468 31328
rect 22462 31288 22468 31300
rect 22520 31288 22526 31340
rect 24596 31337 24624 31368
rect 25590 31356 25596 31408
rect 25648 31356 25654 31408
rect 29457 31399 29515 31405
rect 29457 31396 29469 31399
rect 28092 31368 29469 31396
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31328 27307 31331
rect 27614 31328 27620 31340
rect 27295 31300 27620 31328
rect 27295 31297 27307 31300
rect 27249 31291 27307 31297
rect 27614 31288 27620 31300
rect 27672 31288 27678 31340
rect 27890 31328 27896 31340
rect 27851 31300 27896 31328
rect 27890 31288 27896 31300
rect 27948 31288 27954 31340
rect 28092 31337 28120 31368
rect 29457 31365 29469 31368
rect 29503 31365 29515 31399
rect 29457 31359 29515 31365
rect 28077 31331 28135 31337
rect 28077 31297 28089 31331
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 28169 31331 28227 31337
rect 28169 31297 28181 31331
rect 28215 31328 28227 31331
rect 28350 31328 28356 31340
rect 28215 31300 28356 31328
rect 28215 31297 28227 31300
rect 28169 31291 28227 31297
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 28442 31288 28448 31340
rect 28500 31328 28506 31340
rect 29270 31328 29276 31340
rect 28500 31300 28545 31328
rect 29231 31300 29276 31328
rect 28500 31288 28506 31300
rect 29270 31288 29276 31300
rect 29328 31288 29334 31340
rect 33594 31328 33600 31340
rect 33555 31300 33600 31328
rect 33594 31288 33600 31300
rect 33652 31288 33658 31340
rect 36170 31288 36176 31340
rect 36228 31328 36234 31340
rect 36541 31331 36599 31337
rect 36541 31328 36553 31331
rect 36228 31300 36553 31328
rect 36228 31288 36234 31300
rect 36541 31297 36553 31300
rect 36587 31297 36599 31331
rect 36541 31291 36599 31297
rect 36725 31331 36783 31337
rect 36725 31297 36737 31331
rect 36771 31328 36783 31331
rect 37090 31328 37096 31340
rect 36771 31300 37096 31328
rect 36771 31297 36783 31300
rect 36725 31291 36783 31297
rect 37090 31288 37096 31300
rect 37148 31288 37154 31340
rect 37274 31328 37280 31340
rect 37235 31300 37280 31328
rect 37274 31288 37280 31300
rect 37332 31288 37338 31340
rect 10778 31220 10784 31272
rect 10836 31260 10842 31272
rect 12894 31260 12900 31272
rect 10836 31232 12756 31260
rect 12855 31232 12900 31260
rect 10836 31220 10842 31232
rect 12161 31195 12219 31201
rect 10520 31164 11284 31192
rect 9490 31124 9496 31136
rect 9451 31096 9496 31124
rect 9490 31084 9496 31096
rect 9548 31084 9554 31136
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 10137 31127 10195 31133
rect 10137 31124 10149 31127
rect 9732 31096 10149 31124
rect 9732 31084 9738 31096
rect 10137 31093 10149 31096
rect 10183 31093 10195 31127
rect 10137 31087 10195 31093
rect 10686 31084 10692 31136
rect 10744 31124 10750 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 10744 31096 10793 31124
rect 10744 31084 10750 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 11256 31124 11284 31164
rect 12161 31161 12173 31195
rect 12207 31192 12219 31195
rect 12526 31192 12532 31204
rect 12207 31164 12532 31192
rect 12207 31161 12219 31164
rect 12161 31155 12219 31161
rect 12526 31152 12532 31164
rect 12584 31152 12590 31204
rect 12434 31124 12440 31136
rect 11256 31096 12440 31124
rect 10781 31087 10839 31093
rect 12434 31084 12440 31096
rect 12492 31084 12498 31136
rect 12728 31124 12756 31232
rect 12894 31220 12900 31232
rect 12952 31220 12958 31272
rect 14642 31260 14648 31272
rect 13004 31232 14648 31260
rect 12802 31152 12808 31204
rect 12860 31192 12866 31204
rect 13004 31192 13032 31232
rect 14642 31220 14648 31232
rect 14700 31220 14706 31272
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31260 15439 31263
rect 16206 31260 16212 31272
rect 15427 31232 16212 31260
rect 15427 31229 15439 31232
rect 15381 31223 15439 31229
rect 16206 31220 16212 31232
rect 16264 31220 16270 31272
rect 17862 31260 17868 31272
rect 17823 31232 17868 31260
rect 17862 31220 17868 31232
rect 17920 31220 17926 31272
rect 18138 31260 18144 31272
rect 18099 31232 18144 31260
rect 18138 31220 18144 31232
rect 18196 31220 18202 31272
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 19150 31260 19156 31272
rect 18288 31232 19156 31260
rect 18288 31220 18294 31232
rect 19150 31220 19156 31232
rect 19208 31260 19214 31272
rect 19613 31263 19671 31269
rect 19613 31260 19625 31263
rect 19208 31232 19625 31260
rect 19208 31220 19214 31232
rect 19613 31229 19625 31232
rect 19659 31229 19671 31263
rect 22554 31260 22560 31272
rect 22467 31232 22560 31260
rect 19613 31223 19671 31229
rect 22554 31220 22560 31232
rect 22612 31260 22618 31272
rect 23014 31260 23020 31272
rect 22612 31232 23020 31260
rect 22612 31220 22618 31232
rect 23014 31220 23020 31232
rect 23072 31220 23078 31272
rect 24854 31260 24860 31272
rect 24815 31232 24860 31260
rect 24854 31220 24860 31232
rect 24912 31220 24918 31272
rect 28261 31263 28319 31269
rect 28261 31229 28273 31263
rect 28307 31229 28319 31263
rect 28261 31223 28319 31229
rect 29089 31263 29147 31269
rect 29089 31229 29101 31263
rect 29135 31260 29147 31263
rect 29178 31260 29184 31272
rect 29135 31232 29184 31260
rect 29135 31229 29147 31232
rect 29089 31223 29147 31229
rect 28276 31192 28304 31223
rect 29178 31220 29184 31232
rect 29236 31220 29242 31272
rect 33502 31260 33508 31272
rect 33463 31232 33508 31260
rect 33502 31220 33508 31232
rect 33560 31220 33566 31272
rect 33965 31263 34023 31269
rect 33965 31229 33977 31263
rect 34011 31260 34023 31263
rect 34514 31260 34520 31272
rect 34011 31232 34520 31260
rect 34011 31229 34023 31232
rect 33965 31223 34023 31229
rect 34514 31220 34520 31232
rect 34572 31220 34578 31272
rect 12860 31164 13032 31192
rect 14200 31164 17356 31192
rect 12860 31152 12866 31164
rect 14200 31124 14228 31164
rect 12728 31096 14228 31124
rect 17034 31084 17040 31136
rect 17092 31124 17098 31136
rect 17221 31127 17279 31133
rect 17221 31124 17233 31127
rect 17092 31096 17233 31124
rect 17092 31084 17098 31096
rect 17221 31093 17233 31096
rect 17267 31093 17279 31127
rect 17328 31124 17356 31164
rect 19168 31164 24716 31192
rect 19168 31124 19196 31164
rect 17328 31096 19196 31124
rect 17221 31087 17279 31093
rect 22094 31084 22100 31136
rect 22152 31124 22158 31136
rect 24688 31124 24716 31164
rect 25884 31164 28304 31192
rect 25884 31124 25912 31164
rect 45554 31152 45560 31204
rect 45612 31192 45618 31204
rect 46014 31192 46020 31204
rect 45612 31164 46020 31192
rect 45612 31152 45618 31164
rect 46014 31152 46020 31164
rect 46072 31152 46078 31204
rect 22152 31096 22197 31124
rect 24688 31096 25912 31124
rect 22152 31084 22158 31096
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 26329 31127 26387 31133
rect 26329 31124 26341 31127
rect 26016 31096 26341 31124
rect 26016 31084 26022 31096
rect 26329 31093 26341 31096
rect 26375 31093 26387 31127
rect 26329 31087 26387 31093
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 29638 31124 29644 31136
rect 29052 31096 29644 31124
rect 29052 31084 29058 31096
rect 29638 31084 29644 31096
rect 29696 31084 29702 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 7834 30880 7840 30932
rect 7892 30920 7898 30932
rect 12894 30920 12900 30932
rect 7892 30892 12434 30920
rect 12855 30892 12900 30920
rect 7892 30880 7898 30892
rect 9490 30812 9496 30864
rect 9548 30852 9554 30864
rect 12406 30852 12434 30892
rect 12894 30880 12900 30892
rect 12952 30880 12958 30932
rect 14182 30920 14188 30932
rect 14143 30892 14188 30920
rect 14182 30880 14188 30892
rect 14240 30880 14246 30932
rect 18049 30923 18107 30929
rect 18049 30889 18061 30923
rect 18095 30920 18107 30923
rect 18138 30920 18144 30932
rect 18095 30892 18144 30920
rect 18095 30889 18107 30892
rect 18049 30883 18107 30889
rect 18138 30880 18144 30892
rect 18196 30880 18202 30932
rect 19242 30880 19248 30932
rect 19300 30920 19306 30932
rect 19337 30923 19395 30929
rect 19337 30920 19349 30923
rect 19300 30892 19349 30920
rect 19300 30880 19306 30892
rect 19337 30889 19349 30892
rect 19383 30889 19395 30923
rect 23385 30923 23443 30929
rect 23385 30920 23397 30923
rect 19337 30883 19395 30889
rect 22066 30892 23397 30920
rect 9548 30824 9812 30852
rect 12406 30824 17264 30852
rect 9548 30812 9554 30824
rect 9674 30784 9680 30796
rect 9635 30756 9680 30784
rect 9674 30744 9680 30756
rect 9732 30744 9738 30796
rect 9784 30784 9812 30824
rect 9953 30787 10011 30793
rect 9953 30784 9965 30787
rect 9784 30756 9965 30784
rect 9953 30753 9965 30756
rect 9999 30753 10011 30787
rect 9953 30747 10011 30753
rect 12434 30676 12440 30728
rect 12492 30716 12498 30728
rect 12710 30716 12716 30728
rect 12492 30688 12716 30716
rect 12492 30676 12498 30688
rect 12710 30676 12716 30688
rect 12768 30716 12774 30728
rect 12897 30719 12955 30725
rect 12897 30716 12909 30719
rect 12768 30688 12909 30716
rect 12768 30676 12774 30688
rect 12897 30685 12909 30688
rect 12943 30685 12955 30719
rect 12897 30679 12955 30685
rect 10686 30608 10692 30660
rect 10744 30608 10750 30660
rect 11701 30651 11759 30657
rect 11701 30617 11713 30651
rect 11747 30648 11759 30651
rect 12618 30648 12624 30660
rect 11747 30620 12624 30648
rect 11747 30617 11759 30620
rect 11701 30611 11759 30617
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 11716 30580 11744 30611
rect 12618 30608 12624 30620
rect 12676 30608 12682 30660
rect 12912 30648 12940 30679
rect 13262 30676 13268 30728
rect 13320 30716 13326 30728
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13320 30688 14105 30716
rect 13320 30676 13326 30688
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 14642 30676 14648 30728
rect 14700 30716 14706 30728
rect 15657 30719 15715 30725
rect 15657 30716 15669 30719
rect 14700 30688 15669 30716
rect 14700 30676 14706 30688
rect 15657 30685 15669 30688
rect 15703 30716 15715 30719
rect 16117 30719 16175 30725
rect 16117 30716 16129 30719
rect 15703 30688 16129 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 16117 30685 16129 30688
rect 16163 30685 16175 30719
rect 16117 30679 16175 30685
rect 16301 30719 16359 30725
rect 16301 30685 16313 30719
rect 16347 30716 16359 30719
rect 17034 30716 17040 30728
rect 16347 30688 17040 30716
rect 16347 30685 16359 30688
rect 16301 30679 16359 30685
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 13354 30648 13360 30660
rect 12912 30620 13360 30648
rect 13354 30608 13360 30620
rect 13412 30608 13418 30660
rect 15473 30651 15531 30657
rect 15473 30617 15485 30651
rect 15519 30648 15531 30651
rect 16850 30648 16856 30660
rect 15519 30620 16856 30648
rect 15519 30617 15531 30620
rect 15473 30611 15531 30617
rect 16850 30608 16856 30620
rect 16908 30608 16914 30660
rect 16206 30580 16212 30592
rect 9456 30552 11744 30580
rect 16167 30552 16212 30580
rect 9456 30540 9462 30552
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 17236 30580 17264 30824
rect 17862 30812 17868 30864
rect 17920 30852 17926 30864
rect 18601 30855 18659 30861
rect 18601 30852 18613 30855
rect 17920 30824 18613 30852
rect 17920 30812 17926 30824
rect 18601 30821 18613 30824
rect 18647 30821 18659 30855
rect 18601 30815 18659 30821
rect 17586 30784 17592 30796
rect 17547 30756 17592 30784
rect 17586 30744 17592 30756
rect 17644 30744 17650 30796
rect 20438 30784 20444 30796
rect 20399 30756 20444 30784
rect 20438 30744 20444 30756
rect 20496 30744 20502 30796
rect 20717 30787 20775 30793
rect 20717 30753 20729 30787
rect 20763 30784 20775 30787
rect 22066 30784 22094 30892
rect 23385 30889 23397 30892
rect 23431 30889 23443 30923
rect 23385 30883 23443 30889
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 25685 30923 25743 30929
rect 25685 30920 25697 30923
rect 24912 30892 25697 30920
rect 24912 30880 24918 30892
rect 25685 30889 25697 30892
rect 25731 30889 25743 30923
rect 25685 30883 25743 30889
rect 26513 30923 26571 30929
rect 26513 30889 26525 30923
rect 26559 30920 26571 30923
rect 27614 30920 27620 30932
rect 26559 30892 27620 30920
rect 26559 30889 26571 30892
rect 26513 30883 26571 30889
rect 27614 30880 27620 30892
rect 27672 30880 27678 30932
rect 27801 30923 27859 30929
rect 27801 30889 27813 30923
rect 27847 30889 27859 30923
rect 27801 30883 27859 30889
rect 23198 30852 23204 30864
rect 22940 30824 23204 30852
rect 22940 30793 22968 30824
rect 23198 30812 23204 30824
rect 23256 30812 23262 30864
rect 25222 30812 25228 30864
rect 25280 30812 25286 30864
rect 26142 30812 26148 30864
rect 26200 30852 26206 30864
rect 27816 30852 27844 30883
rect 27890 30880 27896 30932
rect 27948 30920 27954 30932
rect 28169 30923 28227 30929
rect 28169 30920 28181 30923
rect 27948 30892 28181 30920
rect 27948 30880 27954 30892
rect 28169 30889 28181 30892
rect 28215 30889 28227 30923
rect 28169 30883 28227 30889
rect 28350 30880 28356 30932
rect 28408 30920 28414 30932
rect 29641 30923 29699 30929
rect 29641 30920 29653 30923
rect 28408 30892 29653 30920
rect 28408 30880 28414 30892
rect 29641 30889 29653 30892
rect 29687 30889 29699 30923
rect 29641 30883 29699 30889
rect 30098 30880 30104 30932
rect 30156 30920 30162 30932
rect 31021 30923 31079 30929
rect 31021 30920 31033 30923
rect 30156 30892 31033 30920
rect 30156 30880 30162 30892
rect 31021 30889 31033 30892
rect 31067 30920 31079 30923
rect 32953 30923 33011 30929
rect 31067 30892 32536 30920
rect 31067 30889 31079 30892
rect 31021 30883 31079 30889
rect 28994 30852 29000 30864
rect 26200 30824 29000 30852
rect 26200 30812 26206 30824
rect 28994 30812 29000 30824
rect 29052 30812 29058 30864
rect 29270 30812 29276 30864
rect 29328 30852 29334 30864
rect 31205 30855 31263 30861
rect 31205 30852 31217 30855
rect 29328 30824 31217 30852
rect 29328 30812 29334 30824
rect 31205 30821 31217 30824
rect 31251 30821 31263 30855
rect 31205 30815 31263 30821
rect 20763 30756 22094 30784
rect 22919 30787 22977 30793
rect 20763 30753 20775 30756
rect 20717 30747 20775 30753
rect 22919 30753 22931 30787
rect 22965 30753 22977 30787
rect 22919 30747 22977 30753
rect 17681 30719 17739 30725
rect 17681 30685 17693 30719
rect 17727 30716 17739 30719
rect 18230 30716 18236 30728
rect 17727 30688 18236 30716
rect 17727 30685 17739 30688
rect 17681 30679 17739 30685
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30685 18567 30719
rect 19242 30716 19248 30728
rect 19203 30688 19248 30716
rect 18509 30679 18567 30685
rect 18138 30608 18144 30660
rect 18196 30648 18202 30660
rect 18524 30648 18552 30679
rect 19242 30676 19248 30688
rect 19300 30676 19306 30728
rect 22646 30716 22652 30728
rect 22607 30688 22652 30716
rect 22646 30676 22652 30688
rect 22704 30676 22710 30728
rect 22738 30676 22744 30728
rect 22796 30716 22802 30728
rect 22833 30719 22891 30725
rect 22833 30716 22845 30719
rect 22796 30688 22845 30716
rect 22796 30676 22802 30688
rect 22833 30685 22845 30688
rect 22879 30685 22891 30719
rect 22833 30679 22891 30685
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30716 23259 30719
rect 23474 30716 23480 30728
rect 23247 30688 23480 30716
rect 23247 30685 23259 30688
rect 23201 30679 23259 30685
rect 18196 30620 18552 30648
rect 18196 30608 18202 30620
rect 21174 30608 21180 30660
rect 21232 30608 21238 30660
rect 23032 30648 23060 30679
rect 23474 30676 23480 30688
rect 23532 30676 23538 30728
rect 24946 30716 24952 30728
rect 24907 30688 24952 30716
rect 24946 30676 24952 30688
rect 25004 30676 25010 30728
rect 25038 30676 25044 30728
rect 25096 30716 25102 30728
rect 25240 30725 25268 30812
rect 25406 30744 25412 30796
rect 25464 30784 25470 30796
rect 29288 30784 29316 30812
rect 31662 30784 31668 30796
rect 25464 30756 25636 30784
rect 25464 30744 25470 30756
rect 25133 30719 25191 30725
rect 25133 30716 25145 30719
rect 25096 30688 25145 30716
rect 25096 30676 25102 30688
rect 25133 30685 25145 30688
rect 25179 30685 25191 30719
rect 25133 30679 25191 30685
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30685 25283 30719
rect 25225 30679 25283 30685
rect 25314 30676 25320 30728
rect 25372 30716 25378 30728
rect 25501 30719 25559 30725
rect 25372 30688 25417 30716
rect 25372 30676 25378 30688
rect 25501 30685 25513 30719
rect 25547 30685 25559 30719
rect 25501 30679 25559 30685
rect 22020 30620 23060 30648
rect 22020 30580 22048 30620
rect 24762 30608 24768 30660
rect 24820 30648 24826 30660
rect 25406 30648 25412 30660
rect 24820 30620 25412 30648
rect 24820 30608 24826 30620
rect 25406 30608 25412 30620
rect 25464 30608 25470 30660
rect 17236 30552 22048 30580
rect 22189 30583 22247 30589
rect 22189 30549 22201 30583
rect 22235 30580 22247 30583
rect 22278 30580 22284 30592
rect 22235 30552 22284 30580
rect 22235 30549 22247 30552
rect 22189 30543 22247 30549
rect 22278 30540 22284 30552
rect 22336 30580 22342 30592
rect 23198 30580 23204 30592
rect 22336 30552 23204 30580
rect 22336 30540 22342 30552
rect 23198 30540 23204 30552
rect 23256 30540 23262 30592
rect 23474 30540 23480 30592
rect 23532 30580 23538 30592
rect 25516 30580 25544 30679
rect 25608 30648 25636 30756
rect 28644 30756 29316 30784
rect 30852 30756 31668 30784
rect 25682 30676 25688 30728
rect 25740 30716 25746 30728
rect 28644 30725 28672 30756
rect 27801 30719 27859 30725
rect 27801 30716 27813 30719
rect 25740 30688 27813 30716
rect 25740 30676 25746 30688
rect 27801 30685 27813 30688
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 28629 30719 28687 30725
rect 28629 30685 28641 30719
rect 28675 30685 28687 30719
rect 28629 30679 28687 30685
rect 26237 30651 26295 30657
rect 26237 30648 26249 30651
rect 25608 30620 26249 30648
rect 26237 30617 26249 30620
rect 26283 30617 26295 30651
rect 28000 30648 28028 30679
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 29549 30719 29607 30725
rect 29549 30716 29561 30719
rect 29052 30688 29561 30716
rect 29052 30676 29058 30688
rect 29549 30685 29561 30688
rect 29595 30685 29607 30719
rect 29730 30716 29736 30728
rect 29691 30688 29736 30716
rect 29549 30679 29607 30685
rect 29730 30676 29736 30688
rect 29788 30676 29794 30728
rect 30852 30725 30880 30756
rect 31662 30744 31668 30756
rect 31720 30784 31726 30796
rect 32508 30784 32536 30892
rect 32953 30889 32965 30923
rect 32999 30920 33011 30923
rect 33502 30920 33508 30932
rect 32999 30892 33508 30920
rect 32999 30889 33011 30892
rect 32953 30883 33011 30889
rect 33502 30880 33508 30892
rect 33560 30920 33566 30932
rect 33689 30923 33747 30929
rect 33689 30920 33701 30923
rect 33560 30892 33701 30920
rect 33560 30880 33566 30892
rect 33689 30889 33701 30892
rect 33735 30889 33747 30923
rect 36170 30920 36176 30932
rect 36131 30892 36176 30920
rect 33689 30883 33747 30889
rect 36170 30880 36176 30892
rect 36228 30880 36234 30932
rect 34514 30784 34520 30796
rect 31720 30756 32352 30784
rect 31720 30744 31726 30756
rect 30837 30719 30895 30725
rect 30837 30685 30849 30719
rect 30883 30685 30895 30719
rect 31018 30716 31024 30728
rect 30979 30688 31024 30716
rect 30837 30679 30895 30685
rect 31018 30676 31024 30688
rect 31076 30676 31082 30728
rect 32324 30725 32352 30756
rect 32508 30756 34520 30784
rect 32508 30725 32536 30756
rect 32309 30719 32367 30725
rect 32309 30685 32321 30719
rect 32355 30685 32367 30719
rect 32309 30679 32367 30685
rect 32493 30719 32551 30725
rect 32493 30685 32505 30719
rect 32539 30685 32551 30719
rect 32950 30716 32956 30728
rect 32911 30688 32956 30716
rect 32493 30679 32551 30685
rect 28813 30651 28871 30657
rect 28813 30648 28825 30651
rect 28000 30620 28825 30648
rect 26237 30611 26295 30617
rect 28813 30617 28825 30620
rect 28859 30648 28871 30651
rect 29178 30648 29184 30660
rect 28859 30620 29184 30648
rect 28859 30617 28871 30620
rect 28813 30611 28871 30617
rect 29178 30608 29184 30620
rect 29236 30648 29242 30660
rect 30006 30648 30012 30660
rect 29236 30620 30012 30648
rect 29236 30608 29242 30620
rect 30006 30608 30012 30620
rect 30064 30608 30070 30660
rect 28994 30580 29000 30592
rect 23532 30552 25544 30580
rect 28955 30552 29000 30580
rect 23532 30540 23538 30552
rect 28994 30540 29000 30552
rect 29052 30540 29058 30592
rect 32324 30580 32352 30679
rect 32950 30676 32956 30688
rect 33008 30676 33014 30728
rect 33152 30725 33180 30756
rect 34514 30744 34520 30756
rect 34572 30744 34578 30796
rect 33137 30719 33195 30725
rect 33137 30685 33149 30719
rect 33183 30685 33195 30719
rect 33137 30679 33195 30685
rect 33597 30719 33655 30725
rect 33597 30685 33609 30719
rect 33643 30685 33655 30719
rect 33597 30679 33655 30685
rect 36081 30719 36139 30725
rect 36081 30685 36093 30719
rect 36127 30685 36139 30719
rect 36262 30716 36268 30728
rect 36223 30688 36268 30716
rect 36081 30679 36139 30685
rect 32401 30651 32459 30657
rect 32401 30617 32413 30651
rect 32447 30648 32459 30651
rect 33612 30648 33640 30679
rect 32447 30620 33640 30648
rect 36096 30648 36124 30679
rect 36262 30676 36268 30688
rect 36320 30716 36326 30728
rect 36814 30716 36820 30728
rect 36320 30688 36820 30716
rect 36320 30676 36326 30688
rect 36814 30676 36820 30688
rect 36872 30716 36878 30728
rect 36909 30719 36967 30725
rect 36909 30716 36921 30719
rect 36872 30688 36921 30716
rect 36872 30676 36878 30688
rect 36909 30685 36921 30688
rect 36955 30685 36967 30719
rect 36909 30679 36967 30685
rect 36725 30651 36783 30657
rect 36725 30648 36737 30651
rect 36096 30620 36737 30648
rect 32447 30617 32459 30620
rect 32401 30611 32459 30617
rect 36725 30617 36737 30620
rect 36771 30648 36783 30651
rect 36998 30648 37004 30660
rect 36771 30620 37004 30648
rect 36771 30617 36783 30620
rect 36725 30611 36783 30617
rect 36998 30608 37004 30620
rect 37056 30608 37062 30660
rect 32950 30580 32956 30592
rect 32324 30552 32956 30580
rect 32950 30540 32956 30552
rect 33008 30540 33014 30592
rect 34057 30583 34115 30589
rect 34057 30549 34069 30583
rect 34103 30580 34115 30583
rect 34790 30580 34796 30592
rect 34103 30552 34796 30580
rect 34103 30549 34115 30552
rect 34057 30543 34115 30549
rect 34790 30540 34796 30552
rect 34848 30540 34854 30592
rect 37090 30580 37096 30592
rect 37051 30552 37096 30580
rect 37090 30540 37096 30552
rect 37148 30540 37154 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 17497 30379 17555 30385
rect 17497 30345 17509 30379
rect 17543 30376 17555 30379
rect 17586 30376 17592 30388
rect 17543 30348 17592 30376
rect 17543 30345 17555 30348
rect 17497 30339 17555 30345
rect 17586 30336 17592 30348
rect 17644 30336 17650 30388
rect 22557 30379 22615 30385
rect 22557 30345 22569 30379
rect 22603 30376 22615 30379
rect 22646 30376 22652 30388
rect 22603 30348 22652 30376
rect 22603 30345 22615 30348
rect 22557 30339 22615 30345
rect 22646 30336 22652 30348
rect 22704 30336 22710 30388
rect 24946 30336 24952 30388
rect 25004 30376 25010 30388
rect 26053 30379 26111 30385
rect 26053 30376 26065 30379
rect 25004 30348 26065 30376
rect 25004 30336 25010 30348
rect 26053 30345 26065 30348
rect 26099 30345 26111 30379
rect 26053 30339 26111 30345
rect 13004 30280 16804 30308
rect 9861 30243 9919 30249
rect 9861 30209 9873 30243
rect 9907 30240 9919 30243
rect 11514 30240 11520 30252
rect 9907 30212 11520 30240
rect 9907 30209 9919 30212
rect 9861 30203 9919 30209
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 13004 30249 13032 30280
rect 12989 30243 13047 30249
rect 12989 30209 13001 30243
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 13170 30172 13176 30184
rect 13131 30144 13176 30172
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 13449 30175 13507 30181
rect 13449 30141 13461 30175
rect 13495 30141 13507 30175
rect 13449 30135 13507 30141
rect 3694 30064 3700 30116
rect 3752 30104 3758 30116
rect 13464 30104 13492 30135
rect 3752 30076 13492 30104
rect 16776 30104 16804 30280
rect 17034 30268 17040 30320
rect 17092 30308 17098 30320
rect 17221 30311 17279 30317
rect 17221 30308 17233 30311
rect 17092 30280 17233 30308
rect 17092 30268 17098 30280
rect 17221 30277 17233 30280
rect 17267 30277 17279 30311
rect 21174 30308 21180 30320
rect 21135 30280 21180 30308
rect 17221 30271 17279 30277
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 23014 30308 23020 30320
rect 22975 30280 23020 30308
rect 23014 30268 23020 30280
rect 23072 30268 23078 30320
rect 24670 30308 24676 30320
rect 23860 30280 24676 30308
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 17129 30243 17187 30249
rect 17129 30240 17141 30243
rect 17000 30212 17141 30240
rect 17000 30200 17006 30212
rect 17129 30209 17141 30212
rect 17175 30209 17187 30243
rect 17129 30203 17187 30209
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17368 30212 17461 30240
rect 17368 30200 17374 30212
rect 20990 30200 20996 30252
rect 21048 30240 21054 30252
rect 21085 30243 21143 30249
rect 21085 30240 21097 30243
rect 21048 30212 21097 30240
rect 21048 30200 21054 30212
rect 21085 30209 21097 30212
rect 21131 30209 21143 30243
rect 21085 30203 21143 30209
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22373 30243 22431 30249
rect 22373 30209 22385 30243
rect 22419 30240 22431 30243
rect 22462 30240 22468 30252
rect 22419 30212 22468 30240
rect 22419 30209 22431 30212
rect 22373 30203 22431 30209
rect 16850 30132 16856 30184
rect 16908 30172 16914 30184
rect 17328 30172 17356 30200
rect 16908 30144 17356 30172
rect 16908 30132 16914 30144
rect 16945 30107 17003 30113
rect 16945 30104 16957 30107
rect 16776 30076 16957 30104
rect 3752 30064 3758 30076
rect 16945 30073 16957 30076
rect 16991 30104 17003 30107
rect 17310 30104 17316 30116
rect 16991 30076 17316 30104
rect 16991 30073 17003 30076
rect 16945 30067 17003 30073
rect 17310 30064 17316 30076
rect 17368 30064 17374 30116
rect 22020 30104 22048 30203
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 23198 30240 23204 30252
rect 23159 30212 23204 30240
rect 23198 30200 23204 30212
rect 23256 30200 23262 30252
rect 23860 30104 23888 30280
rect 24670 30268 24676 30280
rect 24728 30268 24734 30320
rect 24765 30311 24823 30317
rect 24765 30277 24777 30311
rect 24811 30308 24823 30311
rect 25038 30308 25044 30320
rect 24811 30280 25044 30308
rect 24811 30277 24823 30280
rect 24765 30271 24823 30277
rect 25038 30268 25044 30280
rect 25096 30268 25102 30320
rect 30009 30311 30067 30317
rect 25240 30280 25912 30308
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 24121 30243 24179 30249
rect 24121 30209 24133 30243
rect 24167 30240 24179 30243
rect 24949 30243 25007 30249
rect 24949 30240 24961 30243
rect 24167 30212 24961 30240
rect 24167 30209 24179 30212
rect 24121 30203 24179 30209
rect 24949 30209 24961 30212
rect 24995 30240 25007 30243
rect 25240 30240 25268 30280
rect 25682 30240 25688 30252
rect 24995 30212 25268 30240
rect 25643 30212 25688 30240
rect 24995 30209 25007 30212
rect 24949 30203 25007 30209
rect 22020 30076 23888 30104
rect 23952 30104 23980 30203
rect 25682 30200 25688 30212
rect 25740 30200 25746 30252
rect 25884 30249 25912 30280
rect 30009 30277 30021 30311
rect 30055 30308 30067 30311
rect 30098 30308 30104 30320
rect 30055 30280 30104 30308
rect 30055 30277 30067 30280
rect 30009 30271 30067 30277
rect 30098 30268 30104 30280
rect 30156 30268 30162 30320
rect 31297 30311 31355 30317
rect 31297 30277 31309 30311
rect 31343 30308 31355 30311
rect 31938 30308 31944 30320
rect 31343 30280 31944 30308
rect 31343 30277 31355 30280
rect 31297 30271 31355 30277
rect 31938 30268 31944 30280
rect 31996 30308 32002 30320
rect 31996 30280 32352 30308
rect 31996 30268 32002 30280
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30240 25927 30243
rect 25958 30240 25964 30252
rect 25915 30212 25964 30240
rect 25915 30209 25927 30212
rect 25869 30203 25927 30209
rect 25958 30200 25964 30212
rect 26016 30200 26022 30252
rect 28629 30243 28687 30249
rect 28629 30209 28641 30243
rect 28675 30240 28687 30243
rect 28994 30240 29000 30252
rect 28675 30212 29000 30240
rect 28675 30209 28687 30212
rect 28629 30203 28687 30209
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 30285 30243 30343 30249
rect 30285 30240 30297 30243
rect 29104 30212 30297 30240
rect 24210 30132 24216 30184
rect 24268 30172 24274 30184
rect 25225 30175 25283 30181
rect 25225 30172 25237 30175
rect 24268 30144 25237 30172
rect 24268 30132 24274 30144
rect 25225 30141 25237 30144
rect 25271 30141 25283 30175
rect 25225 30135 25283 30141
rect 28445 30175 28503 30181
rect 28445 30141 28457 30175
rect 28491 30172 28503 30175
rect 29104 30172 29132 30212
rect 30285 30209 30297 30212
rect 30331 30209 30343 30243
rect 31110 30240 31116 30252
rect 31071 30212 31116 30240
rect 30285 30203 30343 30209
rect 31110 30200 31116 30212
rect 31168 30240 31174 30252
rect 32324 30249 32352 30280
rect 34238 30268 34244 30320
rect 34296 30268 34302 30320
rect 32125 30243 32183 30249
rect 32125 30240 32137 30243
rect 31168 30212 32137 30240
rect 31168 30200 31174 30212
rect 32125 30209 32137 30212
rect 32171 30209 32183 30243
rect 32125 30203 32183 30209
rect 32309 30243 32367 30249
rect 32309 30209 32321 30243
rect 32355 30209 32367 30243
rect 32309 30203 32367 30209
rect 37461 30243 37519 30249
rect 37461 30209 37473 30243
rect 37507 30240 37519 30243
rect 37642 30240 37648 30252
rect 37507 30212 37648 30240
rect 37507 30209 37519 30212
rect 37461 30203 37519 30209
rect 37642 30200 37648 30212
rect 37700 30200 37706 30252
rect 38470 30240 38476 30252
rect 38431 30212 38476 30240
rect 38470 30200 38476 30212
rect 38528 30200 38534 30252
rect 28491 30144 29132 30172
rect 30193 30175 30251 30181
rect 28491 30141 28503 30144
rect 28445 30135 28503 30141
rect 29012 30116 29040 30144
rect 30193 30141 30205 30175
rect 30239 30172 30251 30175
rect 31018 30172 31024 30184
rect 30239 30144 31024 30172
rect 30239 30141 30251 30144
rect 30193 30135 30251 30141
rect 31018 30132 31024 30144
rect 31076 30132 31082 30184
rect 32214 30132 32220 30184
rect 32272 30172 32278 30184
rect 32674 30172 32680 30184
rect 32272 30144 32680 30172
rect 32272 30132 32278 30144
rect 32674 30132 32680 30144
rect 32732 30172 32738 30184
rect 33502 30172 33508 30184
rect 32732 30144 33508 30172
rect 32732 30132 32738 30144
rect 33502 30132 33508 30144
rect 33560 30132 33566 30184
rect 33781 30175 33839 30181
rect 33781 30141 33793 30175
rect 33827 30172 33839 30175
rect 35342 30172 35348 30184
rect 33827 30144 35348 30172
rect 33827 30141 33839 30144
rect 33781 30135 33839 30141
rect 35342 30132 35348 30144
rect 35400 30132 35406 30184
rect 35986 30132 35992 30184
rect 36044 30172 36050 30184
rect 37090 30172 37096 30184
rect 36044 30144 37096 30172
rect 36044 30132 36050 30144
rect 37090 30132 37096 30144
rect 37148 30172 37154 30184
rect 37369 30175 37427 30181
rect 37369 30172 37381 30175
rect 37148 30144 37381 30172
rect 37148 30132 37154 30144
rect 37369 30141 37381 30144
rect 37415 30141 37427 30175
rect 38286 30172 38292 30184
rect 38247 30144 38292 30172
rect 37369 30135 37427 30141
rect 38286 30132 38292 30144
rect 38344 30132 38350 30184
rect 24946 30104 24952 30116
rect 23952 30076 24952 30104
rect 24946 30064 24952 30076
rect 25004 30064 25010 30116
rect 25130 30104 25136 30116
rect 25091 30076 25136 30104
rect 25130 30064 25136 30076
rect 25188 30064 25194 30116
rect 27798 30104 27804 30116
rect 25332 30076 27804 30104
rect 9950 30036 9956 30048
rect 9911 30008 9956 30036
rect 9950 29996 9956 30008
rect 10008 29996 10014 30048
rect 22094 29996 22100 30048
rect 22152 30036 22158 30048
rect 22152 30008 22197 30036
rect 22152 29996 22158 30008
rect 23290 29996 23296 30048
rect 23348 30036 23354 30048
rect 23385 30039 23443 30045
rect 23385 30036 23397 30039
rect 23348 30008 23397 30036
rect 23348 29996 23354 30008
rect 23385 30005 23397 30008
rect 23431 30005 23443 30039
rect 23385 29999 23443 30005
rect 24121 30039 24179 30045
rect 24121 30005 24133 30039
rect 24167 30036 24179 30039
rect 24210 30036 24216 30048
rect 24167 30008 24216 30036
rect 24167 30005 24179 30008
rect 24121 29999 24179 30005
rect 24210 29996 24216 30008
rect 24268 29996 24274 30048
rect 24305 30039 24363 30045
rect 24305 30005 24317 30039
rect 24351 30036 24363 30039
rect 24394 30036 24400 30048
rect 24351 30008 24400 30036
rect 24351 30005 24363 30008
rect 24305 29999 24363 30005
rect 24394 29996 24400 30008
rect 24452 29996 24458 30048
rect 24670 29996 24676 30048
rect 24728 30036 24734 30048
rect 25332 30036 25360 30076
rect 27798 30064 27804 30076
rect 27856 30104 27862 30116
rect 28626 30104 28632 30116
rect 27856 30076 28632 30104
rect 27856 30064 27862 30076
rect 28626 30064 28632 30076
rect 28684 30064 28690 30116
rect 28994 30064 29000 30116
rect 29052 30064 29058 30116
rect 35434 30064 35440 30116
rect 35492 30104 35498 30116
rect 37826 30104 37832 30116
rect 35492 30076 37832 30104
rect 35492 30064 35498 30076
rect 37826 30064 37832 30076
rect 37884 30064 37890 30116
rect 24728 30008 25360 30036
rect 24728 29996 24734 30008
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 25869 30039 25927 30045
rect 25869 30036 25881 30039
rect 25464 30008 25881 30036
rect 25464 29996 25470 30008
rect 25869 30005 25881 30008
rect 25915 30036 25927 30039
rect 26142 30036 26148 30048
rect 25915 30008 26148 30036
rect 25915 30005 25927 30008
rect 25869 29999 25927 30005
rect 26142 29996 26148 30008
rect 26200 29996 26206 30048
rect 28258 29996 28264 30048
rect 28316 30036 28322 30048
rect 28813 30039 28871 30045
rect 28813 30036 28825 30039
rect 28316 30008 28825 30036
rect 28316 29996 28322 30008
rect 28813 30005 28825 30008
rect 28859 30005 28871 30039
rect 30006 30036 30012 30048
rect 29967 30008 30012 30036
rect 28813 29999 28871 30005
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 30469 30039 30527 30045
rect 30469 30005 30481 30039
rect 30515 30036 30527 30039
rect 30558 30036 30564 30048
rect 30515 30008 30564 30036
rect 30515 30005 30527 30008
rect 30469 29999 30527 30005
rect 30558 29996 30564 30008
rect 30616 29996 30622 30048
rect 31478 30036 31484 30048
rect 31439 30008 31484 30036
rect 31478 29996 31484 30008
rect 31536 29996 31542 30048
rect 32217 30039 32275 30045
rect 32217 30005 32229 30039
rect 32263 30036 32275 30039
rect 32858 30036 32864 30048
rect 32263 30008 32864 30036
rect 32263 30005 32275 30008
rect 32217 29999 32275 30005
rect 32858 29996 32864 30008
rect 32916 29996 32922 30048
rect 34514 29996 34520 30048
rect 34572 30036 34578 30048
rect 35253 30039 35311 30045
rect 35253 30036 35265 30039
rect 34572 30008 35265 30036
rect 34572 29996 34578 30008
rect 35253 30005 35265 30008
rect 35299 30005 35311 30039
rect 35253 29999 35311 30005
rect 37458 29996 37464 30048
rect 37516 30036 37522 30048
rect 37737 30039 37795 30045
rect 37737 30036 37749 30039
rect 37516 30008 37749 30036
rect 37516 29996 37522 30008
rect 37737 30005 37749 30008
rect 37783 30005 37795 30039
rect 37737 29999 37795 30005
rect 38010 29996 38016 30048
rect 38068 30036 38074 30048
rect 38657 30039 38715 30045
rect 38657 30036 38669 30039
rect 38068 30008 38669 30036
rect 38068 29996 38074 30008
rect 38657 30005 38669 30008
rect 38703 30005 38715 30039
rect 38657 29999 38715 30005
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 12529 29835 12587 29841
rect 12529 29801 12541 29835
rect 12575 29832 12587 29835
rect 13170 29832 13176 29844
rect 12575 29804 13176 29832
rect 12575 29801 12587 29804
rect 12529 29795 12587 29801
rect 13170 29792 13176 29804
rect 13228 29792 13234 29844
rect 13262 29792 13268 29844
rect 13320 29832 13326 29844
rect 23385 29835 23443 29841
rect 13320 29804 13365 29832
rect 13320 29792 13326 29804
rect 23385 29801 23397 29835
rect 23431 29801 23443 29835
rect 23385 29795 23443 29801
rect 24581 29835 24639 29841
rect 24581 29801 24593 29835
rect 24627 29832 24639 29835
rect 24670 29832 24676 29844
rect 24627 29804 24676 29832
rect 24627 29801 24639 29804
rect 24581 29795 24639 29801
rect 11514 29696 11520 29708
rect 11427 29668 11520 29696
rect 8386 29628 8392 29640
rect 8347 29600 8392 29628
rect 8386 29588 8392 29600
rect 8444 29588 8450 29640
rect 8938 29628 8944 29640
rect 8899 29600 8944 29628
rect 8938 29588 8944 29600
rect 8996 29588 9002 29640
rect 11440 29637 11468 29668
rect 11514 29656 11520 29668
rect 11572 29696 11578 29708
rect 13280 29696 13308 29792
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 20530 29764 20536 29776
rect 13504 29736 20536 29764
rect 13504 29724 13510 29736
rect 20530 29724 20536 29736
rect 20588 29724 20594 29776
rect 23106 29724 23112 29776
rect 23164 29764 23170 29776
rect 23400 29764 23428 29795
rect 24670 29792 24676 29804
rect 24728 29792 24734 29844
rect 25222 29792 25228 29844
rect 25280 29832 25286 29844
rect 25409 29835 25467 29841
rect 25409 29832 25421 29835
rect 25280 29804 25421 29832
rect 25280 29792 25286 29804
rect 25409 29801 25421 29804
rect 25455 29801 25467 29835
rect 25409 29795 25467 29801
rect 27512 29835 27570 29841
rect 27512 29801 27524 29835
rect 27558 29832 27570 29835
rect 28718 29832 28724 29844
rect 27558 29804 28724 29832
rect 27558 29801 27570 29804
rect 27512 29795 27570 29801
rect 28718 29792 28724 29804
rect 28776 29792 28782 29844
rect 28994 29832 29000 29844
rect 28955 29804 29000 29832
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 31110 29792 31116 29844
rect 31168 29832 31174 29844
rect 31297 29835 31355 29841
rect 31297 29832 31309 29835
rect 31168 29804 31309 29832
rect 31168 29792 31174 29804
rect 31297 29801 31309 29804
rect 31343 29801 31355 29835
rect 31662 29832 31668 29844
rect 31623 29804 31668 29832
rect 31297 29795 31355 29801
rect 31312 29764 31340 29795
rect 31662 29792 31668 29804
rect 31720 29792 31726 29844
rect 33965 29835 34023 29841
rect 33965 29801 33977 29835
rect 34011 29832 34023 29835
rect 34238 29832 34244 29844
rect 34011 29804 34244 29832
rect 34011 29801 34023 29804
rect 33965 29795 34023 29801
rect 34238 29792 34244 29804
rect 34296 29792 34302 29844
rect 35342 29832 35348 29844
rect 35303 29804 35348 29832
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 35986 29832 35992 29844
rect 35947 29804 35992 29832
rect 35986 29792 35992 29804
rect 36044 29792 36050 29844
rect 36078 29792 36084 29844
rect 36136 29832 36142 29844
rect 36909 29835 36967 29841
rect 36909 29832 36921 29835
rect 36136 29804 36921 29832
rect 36136 29792 36142 29804
rect 36909 29801 36921 29804
rect 36955 29832 36967 29835
rect 37642 29832 37648 29844
rect 36955 29804 37648 29832
rect 36955 29801 36967 29804
rect 36909 29795 36967 29801
rect 37642 29792 37648 29804
rect 37700 29792 37706 29844
rect 23164 29736 27384 29764
rect 31312 29736 33456 29764
rect 23164 29724 23170 29736
rect 17218 29696 17224 29708
rect 11572 29668 13308 29696
rect 17179 29668 17224 29696
rect 11572 29656 11578 29668
rect 17218 29656 17224 29668
rect 17276 29656 17282 29708
rect 17681 29699 17739 29705
rect 17681 29665 17693 29699
rect 17727 29696 17739 29699
rect 18230 29696 18236 29708
rect 17727 29668 18236 29696
rect 17727 29665 17739 29668
rect 17681 29659 17739 29665
rect 18230 29656 18236 29668
rect 18288 29656 18294 29708
rect 23477 29699 23535 29705
rect 22480 29668 23336 29696
rect 11425 29631 11483 29637
rect 11425 29597 11437 29631
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 12437 29631 12495 29637
rect 12437 29597 12449 29631
rect 12483 29628 12495 29631
rect 12618 29628 12624 29640
rect 12483 29600 12624 29628
rect 12483 29597 12495 29600
rect 12437 29591 12495 29597
rect 12618 29588 12624 29600
rect 12676 29588 12682 29640
rect 12894 29588 12900 29640
rect 12952 29628 12958 29640
rect 13081 29631 13139 29637
rect 13081 29628 13093 29631
rect 12952 29600 13093 29628
rect 12952 29588 12958 29600
rect 13081 29597 13093 29600
rect 13127 29597 13139 29631
rect 13081 29591 13139 29597
rect 13354 29588 13360 29640
rect 13412 29628 13418 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 13412 29600 14289 29628
rect 13412 29588 13418 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 15841 29631 15899 29637
rect 15841 29597 15853 29631
rect 15887 29628 15899 29631
rect 16298 29628 16304 29640
rect 15887 29600 16304 29628
rect 15887 29597 15899 29600
rect 15841 29591 15899 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 17310 29628 17316 29640
rect 17271 29600 17316 29628
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 18138 29628 18144 29640
rect 18099 29600 18144 29628
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 19242 29628 19248 29640
rect 19155 29600 19248 29628
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 22480 29637 22508 29668
rect 23308 29640 23336 29668
rect 23477 29665 23489 29699
rect 23523 29696 23535 29699
rect 23523 29668 24440 29696
rect 23523 29665 23535 29668
rect 23477 29659 23535 29665
rect 24412 29640 24440 29668
rect 25332 29668 26188 29696
rect 22465 29631 22523 29637
rect 22465 29597 22477 29631
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 22554 29588 22560 29640
rect 22612 29628 22618 29640
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 22612 29600 22661 29628
rect 22612 29588 22618 29600
rect 22649 29597 22661 29600
rect 22695 29597 22707 29631
rect 23290 29628 23296 29640
rect 23251 29600 23296 29628
rect 22649 29591 22707 29597
rect 9217 29563 9275 29569
rect 9217 29529 9229 29563
rect 9263 29529 9275 29563
rect 9217 29523 9275 29529
rect 8205 29495 8263 29501
rect 8205 29461 8217 29495
rect 8251 29492 8263 29495
rect 9232 29492 9260 29523
rect 9950 29520 9956 29572
rect 10008 29520 10014 29572
rect 14550 29560 14556 29572
rect 14511 29532 14556 29560
rect 14550 29520 14556 29532
rect 14608 29520 14614 29572
rect 16316 29560 16344 29588
rect 19260 29560 19288 29588
rect 16316 29532 19288 29560
rect 22664 29560 22692 29591
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23566 29628 23572 29640
rect 23527 29600 23572 29628
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 24394 29628 24400 29640
rect 24355 29600 24400 29628
rect 24394 29588 24400 29600
rect 24452 29588 24458 29640
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 25332 29637 25360 29668
rect 25317 29631 25375 29637
rect 24544 29600 24589 29628
rect 24544 29588 24550 29600
rect 25317 29597 25329 29631
rect 25363 29597 25375 29631
rect 25317 29591 25375 29597
rect 25501 29631 25559 29637
rect 25501 29597 25513 29631
rect 25547 29597 25559 29631
rect 25501 29591 25559 29597
rect 25516 29560 25544 29591
rect 22664 29532 25544 29560
rect 26160 29560 26188 29668
rect 26234 29656 26240 29708
rect 26292 29696 26298 29708
rect 27246 29696 27252 29708
rect 26292 29668 27252 29696
rect 26292 29656 26298 29668
rect 27246 29656 27252 29668
rect 27304 29656 27310 29708
rect 27356 29696 27384 29736
rect 31018 29696 31024 29708
rect 27356 29668 31024 29696
rect 31018 29656 31024 29668
rect 31076 29656 31082 29708
rect 31389 29699 31447 29705
rect 31389 29665 31401 29699
rect 31435 29696 31447 29699
rect 31938 29696 31944 29708
rect 31435 29668 31944 29696
rect 31435 29665 31447 29668
rect 31389 29659 31447 29665
rect 31938 29656 31944 29668
rect 31996 29656 32002 29708
rect 32401 29699 32459 29705
rect 32401 29665 32413 29699
rect 32447 29696 32459 29699
rect 33428 29696 33456 29736
rect 33502 29724 33508 29776
rect 33560 29764 33566 29776
rect 33560 29736 37596 29764
rect 33560 29724 33566 29736
rect 32447 29668 33180 29696
rect 33428 29668 34468 29696
rect 32447 29665 32459 29668
rect 32401 29659 32459 29665
rect 26326 29588 26332 29640
rect 26384 29628 26390 29640
rect 26513 29631 26571 29637
rect 26513 29628 26525 29631
rect 26384 29600 26525 29628
rect 26384 29588 26390 29600
rect 26513 29597 26525 29600
rect 26559 29597 26571 29631
rect 26513 29591 26571 29597
rect 29822 29588 29828 29640
rect 29880 29628 29886 29640
rect 29880 29600 30512 29628
rect 29880 29588 29886 29600
rect 27522 29560 27528 29572
rect 26160 29532 27528 29560
rect 10686 29492 10692 29504
rect 8251 29464 9260 29492
rect 10647 29464 10692 29492
rect 8251 29461 8263 29464
rect 8205 29455 8263 29461
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 11422 29452 11428 29504
rect 11480 29492 11486 29504
rect 11517 29495 11575 29501
rect 11517 29492 11529 29495
rect 11480 29464 11529 29492
rect 11480 29452 11486 29464
rect 11517 29461 11529 29464
rect 11563 29461 11575 29495
rect 15930 29492 15936 29504
rect 15891 29464 15936 29492
rect 11517 29455 11575 29461
rect 15930 29452 15936 29464
rect 15988 29452 15994 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 18325 29495 18383 29501
rect 18325 29492 18337 29495
rect 18012 29464 18337 29492
rect 18012 29452 18018 29464
rect 18325 29461 18337 29464
rect 18371 29461 18383 29495
rect 19334 29492 19340 29504
rect 19295 29464 19340 29492
rect 18325 29455 18383 29461
rect 19334 29452 19340 29464
rect 19392 29452 19398 29504
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 22557 29495 22615 29501
rect 22557 29492 22569 29495
rect 22520 29464 22569 29492
rect 22520 29452 22526 29464
rect 22557 29461 22569 29464
rect 22603 29461 22615 29495
rect 22557 29455 22615 29461
rect 23753 29495 23811 29501
rect 23753 29461 23765 29495
rect 23799 29492 23811 29495
rect 23934 29492 23940 29504
rect 23799 29464 23940 29492
rect 23799 29461 23811 29464
rect 23753 29455 23811 29461
rect 23934 29452 23940 29464
rect 23992 29452 23998 29504
rect 24780 29501 24808 29532
rect 27522 29520 27528 29532
rect 27580 29520 27586 29572
rect 28534 29520 28540 29572
rect 28592 29520 28598 29572
rect 30009 29563 30067 29569
rect 30009 29560 30021 29563
rect 28828 29532 30021 29560
rect 24765 29495 24823 29501
rect 24765 29461 24777 29495
rect 24811 29461 24823 29495
rect 26602 29492 26608 29504
rect 26563 29464 26608 29492
rect 24765 29455 24823 29461
rect 26602 29452 26608 29464
rect 26660 29452 26666 29504
rect 27798 29452 27804 29504
rect 27856 29492 27862 29504
rect 28828 29492 28856 29532
rect 30009 29529 30021 29532
rect 30055 29529 30067 29563
rect 30484 29560 30512 29600
rect 30742 29588 30748 29640
rect 30800 29628 30806 29640
rect 31297 29631 31355 29637
rect 31297 29628 31309 29631
rect 30800 29600 31309 29628
rect 30800 29588 30806 29600
rect 31297 29597 31309 29600
rect 31343 29597 31355 29631
rect 31297 29591 31355 29597
rect 31478 29588 31484 29640
rect 31536 29628 31542 29640
rect 32217 29631 32275 29637
rect 32217 29628 32229 29631
rect 31536 29600 32229 29628
rect 31536 29588 31542 29600
rect 32217 29597 32229 29600
rect 32263 29597 32275 29631
rect 32217 29591 32275 29597
rect 32416 29560 32444 29659
rect 32858 29628 32864 29640
rect 32819 29600 32864 29628
rect 32858 29588 32864 29600
rect 32916 29588 32922 29640
rect 33152 29637 33180 29668
rect 33137 29631 33195 29637
rect 33137 29597 33149 29631
rect 33183 29597 33195 29631
rect 33137 29591 33195 29597
rect 33226 29588 33232 29640
rect 33284 29628 33290 29640
rect 33873 29631 33931 29637
rect 33873 29628 33885 29631
rect 33284 29600 33885 29628
rect 33284 29588 33290 29600
rect 33873 29597 33885 29600
rect 33919 29628 33931 29631
rect 33962 29628 33968 29640
rect 33919 29600 33968 29628
rect 33919 29597 33931 29600
rect 33873 29591 33931 29597
rect 33962 29588 33968 29600
rect 34020 29588 34026 29640
rect 34440 29628 34468 29668
rect 34514 29656 34520 29708
rect 34572 29696 34578 29708
rect 35434 29696 35440 29708
rect 34572 29668 35020 29696
rect 34572 29656 34578 29668
rect 34606 29628 34612 29640
rect 34440 29600 34612 29628
rect 34606 29588 34612 29600
rect 34664 29588 34670 29640
rect 34701 29631 34759 29637
rect 34701 29597 34713 29631
rect 34747 29597 34759 29631
rect 34701 29591 34759 29597
rect 33045 29563 33103 29569
rect 33045 29560 33057 29563
rect 30484 29532 32444 29560
rect 32784 29532 33057 29560
rect 30009 29523 30067 29529
rect 32784 29504 32812 29532
rect 33045 29529 33057 29532
rect 33091 29529 33103 29563
rect 33045 29523 33103 29529
rect 27856 29464 28856 29492
rect 27856 29452 27862 29464
rect 29730 29452 29736 29504
rect 29788 29492 29794 29504
rect 30101 29495 30159 29501
rect 30101 29492 30113 29495
rect 29788 29464 30113 29492
rect 29788 29452 29794 29464
rect 30101 29461 30113 29464
rect 30147 29492 30159 29495
rect 32766 29492 32772 29504
rect 30147 29464 32772 29492
rect 30147 29461 30159 29464
rect 30101 29455 30159 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 32950 29492 32956 29504
rect 32911 29464 32956 29492
rect 32950 29452 32956 29464
rect 33008 29452 33014 29504
rect 34716 29492 34744 29591
rect 34790 29588 34796 29640
rect 34848 29628 34854 29640
rect 34992 29628 35020 29668
rect 35268 29668 35440 29696
rect 35069 29631 35127 29637
rect 35069 29628 35081 29631
rect 34848 29600 34893 29628
rect 34992 29600 35081 29628
rect 34848 29588 34854 29600
rect 35069 29597 35081 29600
rect 35115 29597 35127 29631
rect 35069 29591 35127 29597
rect 35166 29631 35224 29637
rect 35166 29597 35178 29631
rect 35212 29628 35224 29631
rect 35268 29628 35296 29668
rect 35434 29656 35440 29668
rect 35492 29656 35498 29708
rect 36173 29699 36231 29705
rect 36173 29665 36185 29699
rect 36219 29696 36231 29699
rect 36814 29696 36820 29708
rect 36219 29668 36492 29696
rect 36775 29668 36820 29696
rect 36219 29665 36231 29668
rect 36173 29659 36231 29665
rect 36464 29640 36492 29668
rect 36814 29656 36820 29668
rect 36872 29656 36878 29708
rect 37568 29705 37596 29736
rect 37553 29699 37611 29705
rect 37553 29665 37565 29699
rect 37599 29665 37611 29699
rect 37553 29659 37611 29665
rect 46934 29656 46940 29708
rect 46992 29696 46998 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 46992 29668 47593 29696
rect 46992 29656 46998 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 35802 29628 35808 29640
rect 35212 29600 35296 29628
rect 35360 29600 35808 29628
rect 35212 29597 35224 29600
rect 35166 29591 35224 29597
rect 34977 29563 35035 29569
rect 34977 29529 34989 29563
rect 35023 29560 35035 29563
rect 35360 29560 35388 29600
rect 35802 29588 35808 29600
rect 35860 29588 35866 29640
rect 35897 29631 35955 29637
rect 35897 29597 35909 29631
rect 35943 29628 35955 29631
rect 36078 29628 36084 29640
rect 35943 29600 36084 29628
rect 35943 29597 35955 29600
rect 35897 29591 35955 29597
rect 36078 29588 36084 29600
rect 36136 29588 36142 29640
rect 36446 29588 36452 29640
rect 36504 29628 36510 29640
rect 36909 29631 36967 29637
rect 36909 29628 36921 29631
rect 36504 29600 36921 29628
rect 36504 29588 36510 29600
rect 36909 29597 36921 29600
rect 36955 29597 36967 29631
rect 36909 29591 36967 29597
rect 47305 29631 47363 29637
rect 47305 29597 47317 29631
rect 47351 29628 47363 29631
rect 47394 29628 47400 29640
rect 47351 29600 47400 29628
rect 47351 29597 47363 29600
rect 47305 29591 47363 29597
rect 47394 29588 47400 29600
rect 47452 29588 47458 29640
rect 35023 29532 35388 29560
rect 35023 29529 35035 29532
rect 34977 29523 35035 29529
rect 35710 29520 35716 29572
rect 35768 29560 35774 29572
rect 36633 29563 36691 29569
rect 35768 29532 36308 29560
rect 35768 29520 35774 29532
rect 35986 29492 35992 29504
rect 34716 29464 35992 29492
rect 35986 29452 35992 29464
rect 36044 29452 36050 29504
rect 36170 29492 36176 29504
rect 36131 29464 36176 29492
rect 36170 29452 36176 29464
rect 36228 29452 36234 29504
rect 36280 29492 36308 29532
rect 36633 29529 36645 29563
rect 36679 29560 36691 29563
rect 36998 29560 37004 29572
rect 36679 29532 37004 29560
rect 36679 29529 36691 29532
rect 36633 29523 36691 29529
rect 36998 29520 37004 29532
rect 37056 29520 37062 29572
rect 37829 29563 37887 29569
rect 37829 29529 37841 29563
rect 37875 29560 37887 29563
rect 37918 29560 37924 29572
rect 37875 29532 37924 29560
rect 37875 29529 37887 29532
rect 37829 29523 37887 29529
rect 37918 29520 37924 29532
rect 37976 29520 37982 29572
rect 38470 29520 38476 29572
rect 38528 29520 38534 29572
rect 37093 29495 37151 29501
rect 37093 29492 37105 29495
rect 36280 29464 37105 29492
rect 37093 29461 37105 29464
rect 37139 29461 37151 29495
rect 37093 29455 37151 29461
rect 37642 29452 37648 29504
rect 37700 29492 37706 29504
rect 39301 29495 39359 29501
rect 39301 29492 39313 29495
rect 37700 29464 39313 29492
rect 37700 29452 37706 29464
rect 39301 29461 39313 29464
rect 39347 29461 39359 29495
rect 39301 29455 39359 29461
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 8386 29248 8392 29300
rect 8444 29288 8450 29300
rect 9217 29291 9275 29297
rect 9217 29288 9229 29291
rect 8444 29260 9229 29288
rect 8444 29248 8450 29260
rect 9217 29257 9229 29260
rect 9263 29257 9275 29291
rect 9217 29251 9275 29257
rect 11977 29291 12035 29297
rect 11977 29257 11989 29291
rect 12023 29288 12035 29291
rect 13354 29288 13360 29300
rect 12023 29260 13360 29288
rect 12023 29257 12035 29260
rect 11977 29251 12035 29257
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 17310 29248 17316 29300
rect 17368 29288 17374 29300
rect 19705 29291 19763 29297
rect 19705 29288 19717 29291
rect 17368 29260 19717 29288
rect 17368 29248 17374 29260
rect 19705 29257 19717 29260
rect 19751 29257 19763 29291
rect 19705 29251 19763 29257
rect 20717 29291 20775 29297
rect 20717 29257 20729 29291
rect 20763 29288 20775 29291
rect 20990 29288 20996 29300
rect 20763 29260 20996 29288
rect 20763 29257 20775 29260
rect 20717 29251 20775 29257
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 22925 29291 22983 29297
rect 22925 29257 22937 29291
rect 22971 29288 22983 29291
rect 23658 29288 23664 29300
rect 22971 29260 23664 29288
rect 22971 29257 22983 29260
rect 22925 29251 22983 29257
rect 23658 29248 23664 29260
rect 23716 29248 23722 29300
rect 25130 29248 25136 29300
rect 25188 29288 25194 29300
rect 25225 29291 25283 29297
rect 25225 29288 25237 29291
rect 25188 29260 25237 29288
rect 25188 29248 25194 29260
rect 25225 29257 25237 29260
rect 25271 29257 25283 29291
rect 25225 29251 25283 29257
rect 27338 29248 27344 29300
rect 27396 29288 27402 29300
rect 28718 29288 28724 29300
rect 27396 29260 27660 29288
rect 28679 29260 28724 29288
rect 27396 29248 27402 29260
rect 8205 29223 8263 29229
rect 8205 29189 8217 29223
rect 8251 29220 8263 29223
rect 8938 29220 8944 29232
rect 8251 29192 8944 29220
rect 8251 29189 8263 29192
rect 8205 29183 8263 29189
rect 8938 29180 8944 29192
rect 8996 29180 9002 29232
rect 14829 29223 14887 29229
rect 14829 29189 14841 29223
rect 14875 29220 14887 29223
rect 18230 29220 18236 29232
rect 14875 29192 17816 29220
rect 18191 29192 18236 29220
rect 14875 29189 14887 29192
rect 14829 29183 14887 29189
rect 7098 29112 7104 29164
rect 7156 29152 7162 29164
rect 7929 29155 7987 29161
rect 7929 29152 7941 29155
rect 7156 29124 7941 29152
rect 7156 29112 7162 29124
rect 7929 29121 7941 29124
rect 7975 29121 7987 29155
rect 8754 29152 8760 29164
rect 8715 29124 8760 29152
rect 7929 29115 7987 29121
rect 7944 29084 7972 29115
rect 8754 29112 8760 29124
rect 8812 29112 8818 29164
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10413 29115 10471 29121
rect 10428 29084 10456 29115
rect 11514 29112 11520 29164
rect 11572 29152 11578 29164
rect 11793 29155 11851 29161
rect 11793 29152 11805 29155
rect 11572 29124 11805 29152
rect 11572 29112 11578 29124
rect 11793 29121 11805 29124
rect 11839 29121 11851 29155
rect 15470 29152 15476 29164
rect 15431 29124 15476 29152
rect 11793 29115 11851 29121
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 17034 29112 17040 29164
rect 17092 29152 17098 29164
rect 17221 29155 17279 29161
rect 17221 29152 17233 29155
rect 17092 29124 17233 29152
rect 17092 29112 17098 29124
rect 17221 29121 17233 29124
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 11146 29084 11152 29096
rect 7944 29056 11152 29084
rect 11146 29044 11152 29056
rect 11204 29044 11210 29096
rect 12158 29044 12164 29096
rect 12216 29084 12222 29096
rect 12989 29087 13047 29093
rect 12989 29084 13001 29087
rect 12216 29056 13001 29084
rect 12216 29044 12222 29056
rect 12989 29053 13001 29056
rect 13035 29053 13047 29087
rect 13170 29084 13176 29096
rect 13131 29056 13176 29084
rect 12989 29047 13047 29053
rect 13170 29044 13176 29056
rect 13228 29044 13234 29096
rect 15565 29087 15623 29093
rect 15565 29053 15577 29087
rect 15611 29084 15623 29087
rect 16206 29084 16212 29096
rect 15611 29056 16212 29084
rect 15611 29053 15623 29056
rect 15565 29047 15623 29053
rect 16206 29044 16212 29056
rect 16264 29044 16270 29096
rect 16850 29044 16856 29096
rect 16908 29084 16914 29096
rect 17129 29087 17187 29093
rect 17129 29084 17141 29087
rect 16908 29056 17141 29084
rect 16908 29044 16914 29056
rect 17129 29053 17141 29056
rect 17175 29053 17187 29087
rect 17310 29084 17316 29096
rect 17271 29056 17316 29084
rect 17129 29047 17187 29053
rect 17310 29044 17316 29056
rect 17368 29044 17374 29096
rect 17405 29087 17463 29093
rect 17405 29053 17417 29087
rect 17451 29053 17463 29087
rect 17788 29084 17816 29192
rect 18230 29180 18236 29192
rect 18288 29180 18294 29232
rect 26237 29223 26295 29229
rect 22296 29192 25176 29220
rect 17954 29152 17960 29164
rect 17915 29124 17960 29152
rect 17954 29112 17960 29124
rect 18012 29112 18018 29164
rect 19334 29112 19340 29164
rect 19392 29112 19398 29164
rect 20530 29152 20536 29164
rect 20491 29124 20536 29152
rect 20530 29112 20536 29124
rect 20588 29152 20594 29164
rect 22296 29161 22324 29192
rect 22281 29155 22339 29161
rect 20588 29124 22232 29152
rect 20588 29112 20594 29124
rect 22204 29084 22232 29124
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 23106 29152 23112 29164
rect 23067 29124 23112 29152
rect 22281 29115 22339 29121
rect 23106 29112 23112 29124
rect 23164 29112 23170 29164
rect 23216 29124 24624 29152
rect 23216 29084 23244 29124
rect 23566 29084 23572 29096
rect 17788 29056 22094 29084
rect 22204 29056 23244 29084
rect 23527 29056 23572 29084
rect 17405 29047 17463 29053
rect 9030 29016 9036 29028
rect 8991 28988 9036 29016
rect 9030 28976 9036 28988
rect 9088 28976 9094 29028
rect 17420 29016 17448 29047
rect 17954 29016 17960 29028
rect 17420 28988 17960 29016
rect 17954 28976 17960 28988
rect 18012 28976 18018 29028
rect 22066 29016 22094 29056
rect 23566 29044 23572 29056
rect 23624 29044 23630 29096
rect 23845 29087 23903 29093
rect 23845 29053 23857 29087
rect 23891 29084 23903 29087
rect 24394 29084 24400 29096
rect 23891 29056 24400 29084
rect 23891 29053 23903 29056
rect 23845 29047 23903 29053
rect 24394 29044 24400 29056
rect 24452 29044 24458 29096
rect 24596 29084 24624 29124
rect 24670 29112 24676 29164
rect 24728 29152 24734 29164
rect 24857 29155 24915 29161
rect 24857 29152 24869 29155
rect 24728 29124 24869 29152
rect 24728 29112 24734 29124
rect 24857 29121 24869 29124
rect 24903 29121 24915 29155
rect 24857 29115 24915 29121
rect 24946 29112 24952 29164
rect 25004 29152 25010 29164
rect 25148 29152 25176 29192
rect 26237 29189 26249 29223
rect 26283 29220 26295 29223
rect 27430 29220 27436 29232
rect 26283 29192 27436 29220
rect 26283 29189 26295 29192
rect 26237 29183 26295 29189
rect 27430 29180 27436 29192
rect 27488 29180 27494 29232
rect 27632 29220 27660 29260
rect 28718 29248 28724 29260
rect 28776 29248 28782 29300
rect 28810 29248 28816 29300
rect 28868 29288 28874 29300
rect 46842 29288 46848 29300
rect 28868 29260 46848 29288
rect 28868 29248 28874 29260
rect 46842 29248 46848 29260
rect 46900 29248 46906 29300
rect 29917 29223 29975 29229
rect 27632 29192 29868 29220
rect 26326 29152 26332 29164
rect 25004 29124 25049 29152
rect 25148 29124 26332 29152
rect 25004 29112 25010 29124
rect 26326 29112 26332 29124
rect 26384 29112 26390 29164
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27338 29152 27344 29164
rect 27120 29124 27344 29152
rect 27120 29112 27126 29124
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 27522 29112 27528 29164
rect 27580 29150 27586 29164
rect 27982 29152 27988 29164
rect 27580 29122 27623 29150
rect 27943 29124 27988 29152
rect 27580 29112 27586 29122
rect 27982 29112 27988 29124
rect 28040 29112 28046 29164
rect 28169 29155 28227 29161
rect 28169 29121 28181 29155
rect 28215 29121 28227 29155
rect 28169 29115 28227 29121
rect 24762 29084 24768 29096
rect 24596 29056 24768 29084
rect 24762 29044 24768 29056
rect 24820 29044 24826 29096
rect 27433 29087 27491 29093
rect 24872 29056 26924 29084
rect 24872 29016 24900 29056
rect 22066 28988 24900 29016
rect 26234 28976 26240 29028
rect 26292 29016 26298 29028
rect 26421 29019 26479 29025
rect 26421 29016 26433 29019
rect 26292 28988 26433 29016
rect 26292 28976 26298 28988
rect 26421 28985 26433 28988
rect 26467 28985 26479 29019
rect 26896 29016 26924 29056
rect 27433 29053 27445 29087
rect 27479 29084 27491 29087
rect 28184 29084 28212 29115
rect 28258 29112 28264 29164
rect 28316 29152 28322 29164
rect 28537 29155 28595 29161
rect 28316 29124 28361 29152
rect 28316 29112 28322 29124
rect 28537 29121 28549 29155
rect 28583 29152 28595 29155
rect 28994 29152 29000 29164
rect 28583 29124 29000 29152
rect 28583 29121 28595 29124
rect 28537 29115 28595 29121
rect 28994 29112 29000 29124
rect 29052 29112 29058 29164
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29840 29152 29868 29192
rect 29917 29189 29929 29223
rect 29963 29220 29975 29223
rect 30558 29220 30564 29232
rect 29963 29192 30564 29220
rect 29963 29189 29975 29192
rect 29917 29183 29975 29189
rect 30558 29180 30564 29192
rect 30616 29180 30622 29232
rect 34977 29223 35035 29229
rect 34977 29220 34989 29223
rect 34178 29192 34989 29220
rect 34977 29189 34989 29192
rect 35023 29189 35035 29223
rect 38010 29220 38016 29232
rect 34977 29183 35035 29189
rect 37292 29192 38016 29220
rect 30837 29155 30895 29161
rect 29840 29124 30604 29152
rect 29733 29115 29791 29121
rect 28350 29084 28356 29096
rect 27479 29056 28212 29084
rect 28311 29056 28356 29084
rect 27479 29053 27491 29056
rect 27433 29047 27491 29053
rect 28350 29044 28356 29056
rect 28408 29044 28414 29096
rect 28810 29044 28816 29096
rect 28868 29044 28874 29096
rect 28828 29016 28856 29044
rect 29748 29016 29776 29115
rect 26896 28988 28856 29016
rect 29196 28988 29776 29016
rect 30101 29019 30159 29025
rect 26421 28979 26479 28985
rect 10410 28948 10416 28960
rect 10371 28920 10416 28948
rect 10410 28908 10416 28920
rect 10468 28908 10474 28960
rect 15286 28908 15292 28960
rect 15344 28948 15350 28960
rect 15749 28951 15807 28957
rect 15749 28948 15761 28951
rect 15344 28920 15761 28948
rect 15344 28908 15350 28920
rect 15749 28917 15761 28920
rect 15795 28917 15807 28951
rect 15749 28911 15807 28917
rect 16945 28951 17003 28957
rect 16945 28917 16957 28951
rect 16991 28948 17003 28951
rect 17402 28948 17408 28960
rect 16991 28920 17408 28948
rect 16991 28917 17003 28920
rect 16945 28911 17003 28917
rect 17402 28908 17408 28920
rect 17460 28908 17466 28960
rect 22370 28948 22376 28960
rect 22331 28920 22376 28948
rect 22370 28908 22376 28920
rect 22428 28908 22434 28960
rect 24394 28908 24400 28960
rect 24452 28948 24458 28960
rect 24857 28951 24915 28957
rect 24857 28948 24869 28951
rect 24452 28920 24869 28948
rect 24452 28908 24458 28920
rect 24857 28917 24869 28920
rect 24903 28917 24915 28951
rect 24857 28911 24915 28917
rect 25682 28908 25688 28960
rect 25740 28948 25746 28960
rect 28810 28948 28816 28960
rect 25740 28920 28816 28948
rect 25740 28908 25746 28920
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 28902 28908 28908 28960
rect 28960 28948 28966 28960
rect 29196 28948 29224 28988
rect 30101 28985 30113 29019
rect 30147 29016 30159 29019
rect 30466 29016 30472 29028
rect 30147 28988 30472 29016
rect 30147 28985 30159 28988
rect 30101 28979 30159 28985
rect 30466 28976 30472 28988
rect 30524 28976 30530 29028
rect 30576 29016 30604 29124
rect 30837 29121 30849 29155
rect 30883 29152 30895 29155
rect 30926 29152 30932 29164
rect 30883 29124 30932 29152
rect 30883 29121 30895 29124
rect 30837 29115 30895 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 32674 29152 32680 29164
rect 32635 29124 32680 29152
rect 32674 29112 32680 29124
rect 32732 29112 32738 29164
rect 34790 29112 34796 29164
rect 34848 29152 34854 29164
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34848 29124 34897 29152
rect 34848 29112 34854 29124
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 35342 29152 35348 29164
rect 34885 29115 34943 29121
rect 34992 29124 35348 29152
rect 30742 29084 30748 29096
rect 30703 29056 30748 29084
rect 30742 29044 30748 29056
rect 30800 29044 30806 29096
rect 33042 29044 33048 29096
rect 33100 29084 33106 29096
rect 34425 29087 34483 29093
rect 34425 29084 34437 29087
rect 33100 29056 34437 29084
rect 33100 29044 33106 29056
rect 34425 29053 34437 29056
rect 34471 29053 34483 29087
rect 34425 29047 34483 29053
rect 34606 29044 34612 29096
rect 34664 29084 34670 29096
rect 34992 29084 35020 29124
rect 35342 29112 35348 29124
rect 35400 29152 35406 29164
rect 37292 29161 37320 29192
rect 38010 29180 38016 29192
rect 38068 29180 38074 29232
rect 38470 29220 38476 29232
rect 38431 29192 38476 29220
rect 38470 29180 38476 29192
rect 38528 29180 38534 29232
rect 37458 29161 37464 29164
rect 35989 29155 36047 29161
rect 35989 29152 36001 29155
rect 35400 29124 36001 29152
rect 35400 29112 35406 29124
rect 35989 29121 36001 29124
rect 36035 29121 36047 29155
rect 35989 29115 36047 29121
rect 37277 29155 37335 29161
rect 37277 29121 37289 29155
rect 37323 29121 37335 29155
rect 37277 29115 37335 29121
rect 37425 29155 37464 29161
rect 37425 29121 37437 29155
rect 37425 29115 37464 29121
rect 37458 29112 37464 29115
rect 37516 29112 37522 29164
rect 37553 29155 37611 29161
rect 37553 29121 37565 29155
rect 37599 29121 37611 29155
rect 37553 29115 37611 29121
rect 35710 29084 35716 29096
rect 34664 29056 35020 29084
rect 35671 29056 35716 29084
rect 34664 29044 34670 29056
rect 35710 29044 35716 29056
rect 35768 29044 35774 29096
rect 35802 29044 35808 29096
rect 35860 29084 35866 29096
rect 37568 29084 37596 29115
rect 37642 29112 37648 29164
rect 37700 29152 37706 29164
rect 37826 29161 37832 29164
rect 37783 29155 37832 29161
rect 37700 29124 37745 29152
rect 37700 29112 37706 29124
rect 37783 29121 37795 29155
rect 37829 29121 37832 29155
rect 37783 29115 37832 29121
rect 37826 29112 37832 29115
rect 37884 29112 37890 29164
rect 38381 29155 38439 29161
rect 38381 29121 38393 29155
rect 38427 29121 38439 29155
rect 38381 29115 38439 29121
rect 38396 29084 38424 29115
rect 35860 29056 37596 29084
rect 37752 29056 38424 29084
rect 35860 29044 35866 29056
rect 37752 29028 37780 29056
rect 31021 29019 31079 29025
rect 31021 29016 31033 29019
rect 30576 28988 31033 29016
rect 31021 28985 31033 28988
rect 31067 28985 31079 29019
rect 31021 28979 31079 28985
rect 34790 28976 34796 29028
rect 34848 29016 34854 29028
rect 37274 29016 37280 29028
rect 34848 28988 37280 29016
rect 34848 28976 34854 28988
rect 37274 28976 37280 28988
rect 37332 29016 37338 29028
rect 37734 29016 37740 29028
rect 37332 28988 37740 29016
rect 37332 28976 37338 28988
rect 37734 28976 37740 28988
rect 37792 28976 37798 29028
rect 37918 29016 37924 29028
rect 37879 28988 37924 29016
rect 37918 28976 37924 28988
rect 37976 28976 37982 29028
rect 30834 28948 30840 28960
rect 28960 28920 29224 28948
rect 30795 28920 30840 28948
rect 28960 28908 28966 28920
rect 30834 28908 30840 28920
rect 30892 28908 30898 28960
rect 32398 28908 32404 28960
rect 32456 28948 32462 28960
rect 32934 28951 32992 28957
rect 32934 28948 32946 28951
rect 32456 28920 32946 28948
rect 32456 28908 32462 28920
rect 32934 28917 32946 28920
rect 32980 28917 32992 28951
rect 32934 28911 32992 28917
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 12158 28744 12164 28756
rect 9600 28716 12164 28744
rect 9490 28608 9496 28620
rect 9451 28580 9496 28608
rect 9490 28568 9496 28580
rect 9548 28568 9554 28620
rect 9600 28552 9628 28716
rect 12158 28704 12164 28716
rect 12216 28704 12222 28756
rect 12713 28747 12771 28753
rect 12713 28713 12725 28747
rect 12759 28744 12771 28747
rect 13170 28744 13176 28756
rect 12759 28716 13176 28744
rect 12759 28713 12771 28716
rect 12713 28707 12771 28713
rect 13170 28704 13176 28716
rect 13228 28704 13234 28756
rect 15470 28704 15476 28756
rect 15528 28744 15534 28756
rect 16393 28747 16451 28753
rect 16393 28744 16405 28747
rect 15528 28716 16405 28744
rect 15528 28704 15534 28716
rect 16393 28713 16405 28716
rect 16439 28744 16451 28747
rect 17310 28744 17316 28756
rect 16439 28716 17316 28744
rect 16439 28713 16451 28716
rect 16393 28707 16451 28713
rect 17310 28704 17316 28716
rect 17368 28704 17374 28756
rect 23658 28704 23664 28756
rect 23716 28744 23722 28756
rect 24489 28747 24547 28753
rect 24489 28744 24501 28747
rect 23716 28716 24501 28744
rect 23716 28704 23722 28716
rect 24489 28713 24501 28716
rect 24535 28744 24547 28747
rect 24670 28744 24676 28756
rect 24535 28716 24676 28744
rect 24535 28713 24547 28716
rect 24489 28707 24547 28713
rect 24670 28704 24676 28716
rect 24728 28704 24734 28756
rect 24946 28704 24952 28756
rect 25004 28744 25010 28756
rect 26973 28747 27031 28753
rect 26973 28744 26985 28747
rect 25004 28716 26985 28744
rect 25004 28704 25010 28716
rect 26973 28713 26985 28716
rect 27019 28713 27031 28747
rect 26973 28707 27031 28713
rect 28445 28747 28503 28753
rect 28445 28713 28457 28747
rect 28491 28744 28503 28747
rect 28534 28744 28540 28756
rect 28491 28716 28540 28744
rect 28491 28713 28503 28716
rect 28445 28707 28503 28713
rect 28534 28704 28540 28716
rect 28592 28704 28598 28756
rect 30834 28744 30840 28756
rect 30747 28716 30840 28744
rect 30834 28704 30840 28716
rect 30892 28704 30898 28756
rect 31018 28744 31024 28756
rect 30979 28716 31024 28744
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 32398 28744 32404 28756
rect 32359 28716 32404 28744
rect 32398 28704 32404 28716
rect 32456 28704 32462 28756
rect 33502 28704 33508 28756
rect 33560 28744 33566 28756
rect 33778 28744 33784 28756
rect 33560 28716 33784 28744
rect 33560 28704 33566 28716
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 35986 28704 35992 28756
rect 36044 28744 36050 28756
rect 38841 28747 38899 28753
rect 38841 28744 38853 28747
rect 36044 28716 38853 28744
rect 36044 28704 36050 28716
rect 38841 28713 38853 28716
rect 38887 28713 38899 28747
rect 38841 28707 38899 28713
rect 17402 28676 17408 28688
rect 17363 28648 17408 28676
rect 17402 28636 17408 28648
rect 17460 28636 17466 28688
rect 17770 28636 17776 28688
rect 17828 28676 17834 28688
rect 23474 28676 23480 28688
rect 17828 28648 22508 28676
rect 17828 28636 17834 28648
rect 10410 28608 10416 28620
rect 10371 28580 10416 28608
rect 10410 28568 10416 28580
rect 10468 28568 10474 28620
rect 14550 28568 14556 28620
rect 14608 28608 14614 28620
rect 14645 28611 14703 28617
rect 14645 28608 14657 28611
rect 14608 28580 14657 28608
rect 14608 28568 14614 28580
rect 14645 28577 14657 28580
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 14921 28611 14979 28617
rect 14921 28577 14933 28611
rect 14967 28608 14979 28611
rect 15286 28608 15292 28620
rect 14967 28580 15292 28608
rect 14967 28577 14979 28580
rect 14921 28571 14979 28577
rect 15286 28568 15292 28580
rect 15344 28568 15350 28620
rect 17129 28611 17187 28617
rect 17129 28577 17141 28611
rect 17175 28608 17187 28611
rect 17218 28608 17224 28620
rect 17175 28580 17224 28608
rect 17175 28577 17187 28580
rect 17129 28571 17187 28577
rect 17218 28568 17224 28580
rect 17276 28568 17282 28620
rect 17310 28568 17316 28620
rect 17368 28608 17374 28620
rect 17368 28580 18276 28608
rect 17368 28568 17374 28580
rect 9582 28540 9588 28552
rect 9495 28512 9588 28540
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 12618 28540 12624 28552
rect 12579 28512 12624 28540
rect 12618 28500 12624 28512
rect 12676 28500 12682 28552
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28540 13415 28543
rect 13446 28540 13452 28552
rect 13403 28512 13452 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 13446 28500 13452 28512
rect 13504 28500 13510 28552
rect 17954 28500 17960 28552
rect 18012 28540 18018 28552
rect 18248 28549 18276 28580
rect 18049 28543 18107 28549
rect 18049 28540 18061 28543
rect 18012 28512 18061 28540
rect 18012 28500 18018 28512
rect 18049 28509 18061 28512
rect 18095 28509 18107 28543
rect 18049 28503 18107 28509
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28540 18291 28543
rect 20165 28543 20223 28549
rect 20165 28540 20177 28543
rect 18279 28512 20177 28540
rect 18279 28509 18291 28512
rect 18233 28503 18291 28509
rect 20165 28509 20177 28512
rect 20211 28509 20223 28543
rect 20165 28503 20223 28509
rect 10689 28475 10747 28481
rect 10689 28441 10701 28475
rect 10735 28441 10747 28475
rect 10689 28435 10747 28441
rect 9953 28407 10011 28413
rect 9953 28373 9965 28407
rect 9999 28404 10011 28407
rect 10704 28404 10732 28435
rect 11422 28432 11428 28484
rect 11480 28432 11486 28484
rect 15930 28432 15936 28484
rect 15988 28432 15994 28484
rect 16942 28432 16948 28484
rect 17000 28472 17006 28484
rect 18417 28475 18475 28481
rect 18417 28472 18429 28475
rect 17000 28444 18429 28472
rect 17000 28432 17006 28444
rect 18417 28441 18429 28444
rect 18463 28441 18475 28475
rect 20346 28472 20352 28484
rect 20307 28444 20352 28472
rect 18417 28435 18475 28441
rect 20346 28432 20352 28444
rect 20404 28432 20410 28484
rect 22002 28472 22008 28484
rect 21963 28444 22008 28472
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 22480 28472 22508 28648
rect 22848 28648 23480 28676
rect 22848 28608 22876 28648
rect 23474 28636 23480 28648
rect 23532 28676 23538 28688
rect 24210 28676 24216 28688
rect 23532 28648 24216 28676
rect 23532 28636 23538 28648
rect 24210 28636 24216 28648
rect 24268 28636 24274 28688
rect 25130 28676 25136 28688
rect 24320 28648 25136 28676
rect 23750 28608 23756 28620
rect 22756 28580 22876 28608
rect 23124 28580 23756 28608
rect 22756 28549 22784 28580
rect 23124 28549 23152 28580
rect 23750 28568 23756 28580
rect 23808 28568 23814 28620
rect 22741 28543 22799 28549
rect 22741 28509 22753 28543
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 23109 28543 23167 28549
rect 23109 28509 23121 28543
rect 23155 28509 23167 28543
rect 23109 28503 23167 28509
rect 23661 28543 23719 28549
rect 23661 28509 23673 28543
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28540 23903 28543
rect 24320 28540 24348 28648
rect 25130 28636 25136 28648
rect 25188 28636 25194 28688
rect 30852 28676 30880 28704
rect 35710 28676 35716 28688
rect 30852 28648 35716 28676
rect 35710 28636 35716 28648
rect 35768 28636 35774 28688
rect 46106 28636 46112 28688
rect 46164 28676 46170 28688
rect 46164 28648 47072 28676
rect 46164 28636 46170 28648
rect 24673 28611 24731 28617
rect 24673 28577 24685 28611
rect 24719 28608 24731 28611
rect 24946 28608 24952 28620
rect 24719 28580 24952 28608
rect 24719 28577 24731 28580
rect 24673 28571 24731 28577
rect 24946 28568 24952 28580
rect 25004 28568 25010 28620
rect 26234 28608 26240 28620
rect 25240 28580 26240 28608
rect 25240 28552 25268 28580
rect 26234 28568 26240 28580
rect 26292 28568 26298 28620
rect 27798 28608 27804 28620
rect 27632 28580 27804 28608
rect 23891 28512 24348 28540
rect 23891 28509 23903 28512
rect 23845 28503 23903 28509
rect 22848 28472 22876 28503
rect 22480 28444 22876 28472
rect 22940 28472 22968 28503
rect 23474 28472 23480 28484
rect 22940 28444 23480 28472
rect 23474 28432 23480 28444
rect 23532 28432 23538 28484
rect 23676 28472 23704 28503
rect 24394 28500 24400 28552
rect 24452 28540 24458 28552
rect 25222 28540 25228 28552
rect 24452 28512 24497 28540
rect 25183 28512 25228 28540
rect 24452 28500 24458 28512
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 26602 28500 26608 28552
rect 26660 28500 26666 28552
rect 27632 28549 27660 28580
rect 27798 28568 27804 28580
rect 27856 28568 27862 28620
rect 28810 28568 28816 28620
rect 28868 28608 28874 28620
rect 30742 28608 30748 28620
rect 28868 28580 29776 28608
rect 30655 28580 30748 28608
rect 28868 28568 28874 28580
rect 27617 28543 27675 28549
rect 27617 28509 27629 28543
rect 27663 28509 27675 28543
rect 27617 28503 27675 28509
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 28353 28543 28411 28549
rect 28353 28540 28365 28543
rect 27764 28512 28365 28540
rect 27764 28500 27770 28512
rect 28353 28509 28365 28512
rect 28399 28509 28411 28543
rect 29638 28540 29644 28552
rect 29599 28512 29644 28540
rect 28353 28503 28411 28509
rect 29638 28500 29644 28512
rect 29696 28500 29702 28552
rect 29748 28549 29776 28580
rect 30742 28568 30748 28580
rect 30800 28608 30806 28620
rect 31478 28608 31484 28620
rect 30800 28580 31484 28608
rect 30800 28568 30806 28580
rect 31478 28568 31484 28580
rect 31536 28568 31542 28620
rect 32950 28608 32956 28620
rect 31680 28580 32956 28608
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28509 29791 28543
rect 29733 28503 29791 28509
rect 30466 28500 30472 28552
rect 30524 28540 30530 28552
rect 31680 28549 31708 28580
rect 32950 28568 32956 28580
rect 33008 28568 33014 28620
rect 36170 28608 36176 28620
rect 35176 28580 36176 28608
rect 30561 28543 30619 28549
rect 30561 28540 30573 28543
rect 30524 28512 30573 28540
rect 30524 28500 30530 28512
rect 30561 28509 30573 28512
rect 30607 28509 30619 28543
rect 30561 28503 30619 28509
rect 30837 28543 30895 28549
rect 30837 28509 30849 28543
rect 30883 28509 30895 28543
rect 30837 28503 30895 28509
rect 31665 28543 31723 28549
rect 31665 28509 31677 28543
rect 31711 28509 31723 28543
rect 31846 28540 31852 28552
rect 31807 28512 31852 28540
rect 31665 28503 31723 28509
rect 24673 28475 24731 28481
rect 24673 28472 24685 28475
rect 23676 28444 24685 28472
rect 24673 28441 24685 28444
rect 24719 28441 24731 28475
rect 25498 28472 25504 28484
rect 25459 28444 25504 28472
rect 24673 28435 24731 28441
rect 25498 28432 25504 28444
rect 25556 28432 25562 28484
rect 27522 28432 27528 28484
rect 27580 28472 27586 28484
rect 27801 28475 27859 28481
rect 27801 28472 27813 28475
rect 27580 28444 27813 28472
rect 27580 28432 27586 28444
rect 27801 28441 27813 28444
rect 27847 28472 27859 28475
rect 29178 28472 29184 28484
rect 27847 28444 29184 28472
rect 27847 28441 27859 28444
rect 27801 28435 27859 28441
rect 29178 28432 29184 28444
rect 29236 28432 29242 28484
rect 29917 28475 29975 28481
rect 29917 28441 29929 28475
rect 29963 28472 29975 28475
rect 30190 28472 30196 28484
rect 29963 28444 30196 28472
rect 29963 28441 29975 28444
rect 29917 28435 29975 28441
rect 30190 28432 30196 28444
rect 30248 28432 30254 28484
rect 30852 28472 30880 28503
rect 31846 28500 31852 28512
rect 31904 28500 31910 28552
rect 31938 28500 31944 28552
rect 31996 28540 32002 28552
rect 32122 28549 32128 28552
rect 32079 28543 32128 28549
rect 31996 28512 32041 28540
rect 31996 28500 32002 28512
rect 32079 28509 32091 28543
rect 32125 28509 32128 28543
rect 32079 28503 32128 28509
rect 32122 28500 32128 28503
rect 32180 28500 32186 28552
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28540 32275 28543
rect 32674 28540 32680 28552
rect 32263 28512 32680 28540
rect 32263 28509 32275 28512
rect 32217 28503 32275 28509
rect 32674 28500 32680 28512
rect 32732 28500 32738 28552
rect 33042 28540 33048 28552
rect 33003 28512 33048 28540
rect 33042 28500 33048 28512
rect 33100 28500 33106 28552
rect 35176 28549 35204 28580
rect 36170 28568 36176 28580
rect 36228 28568 36234 28620
rect 36449 28611 36507 28617
rect 36449 28577 36461 28611
rect 36495 28608 36507 28611
rect 36538 28608 36544 28620
rect 36495 28580 36544 28608
rect 36495 28577 36507 28580
rect 36449 28571 36507 28577
rect 36538 28568 36544 28580
rect 36596 28568 36602 28620
rect 38286 28568 38292 28620
rect 38344 28608 38350 28620
rect 38473 28611 38531 28617
rect 38473 28608 38485 28611
rect 38344 28580 38485 28608
rect 38344 28568 38350 28580
rect 38473 28577 38485 28580
rect 38519 28577 38531 28611
rect 38473 28571 38531 28577
rect 46477 28611 46535 28617
rect 46477 28577 46489 28611
rect 46523 28608 46535 28611
rect 46934 28608 46940 28620
rect 46523 28580 46940 28608
rect 46523 28577 46535 28580
rect 46477 28571 46535 28577
rect 46934 28568 46940 28580
rect 46992 28568 46998 28620
rect 47044 28617 47072 28648
rect 47029 28611 47087 28617
rect 47029 28577 47041 28611
rect 47075 28577 47087 28611
rect 47029 28571 47087 28577
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28509 35219 28543
rect 35342 28540 35348 28552
rect 35303 28512 35348 28540
rect 35161 28503 35219 28509
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 38657 28543 38715 28549
rect 38657 28509 38669 28543
rect 38703 28540 38715 28543
rect 39022 28540 39028 28552
rect 38703 28512 39028 28540
rect 38703 28509 38715 28512
rect 38657 28503 38715 28509
rect 39022 28500 39028 28512
rect 39080 28500 39086 28552
rect 46290 28540 46296 28552
rect 46251 28512 46296 28540
rect 46290 28500 46296 28512
rect 46348 28500 46354 28552
rect 30926 28472 30932 28484
rect 30839 28444 30932 28472
rect 30926 28432 30932 28444
rect 30984 28472 30990 28484
rect 33060 28472 33088 28500
rect 30984 28444 33088 28472
rect 30984 28432 30990 28444
rect 33502 28432 33508 28484
rect 33560 28472 33566 28484
rect 33689 28475 33747 28481
rect 33689 28472 33701 28475
rect 33560 28444 33701 28472
rect 33560 28432 33566 28444
rect 33689 28441 33701 28444
rect 33735 28441 33747 28475
rect 33689 28435 33747 28441
rect 36173 28475 36231 28481
rect 36173 28441 36185 28475
rect 36219 28472 36231 28475
rect 36446 28472 36452 28484
rect 36219 28444 36452 28472
rect 36219 28441 36231 28444
rect 36173 28435 36231 28441
rect 36446 28432 36452 28444
rect 36504 28432 36510 28484
rect 13446 28404 13452 28416
rect 9999 28376 10732 28404
rect 13407 28376 13452 28404
rect 9999 28373 10011 28376
rect 9953 28367 10011 28373
rect 13446 28364 13452 28376
rect 13504 28364 13510 28416
rect 17402 28364 17408 28416
rect 17460 28404 17466 28416
rect 17589 28407 17647 28413
rect 17589 28404 17601 28407
rect 17460 28376 17601 28404
rect 17460 28364 17466 28376
rect 17589 28373 17601 28376
rect 17635 28373 17647 28407
rect 17589 28367 17647 28373
rect 22094 28364 22100 28416
rect 22152 28404 22158 28416
rect 22465 28407 22523 28413
rect 22465 28404 22477 28407
rect 22152 28376 22477 28404
rect 22152 28364 22158 28376
rect 22465 28373 22477 28376
rect 22511 28373 22523 28407
rect 23842 28404 23848 28416
rect 23803 28376 23848 28404
rect 22465 28367 22523 28373
rect 23842 28364 23848 28376
rect 23900 28364 23906 28416
rect 28350 28364 28356 28416
rect 28408 28404 28414 28416
rect 31846 28404 31852 28416
rect 28408 28376 31852 28404
rect 28408 28364 28414 28376
rect 31846 28364 31852 28376
rect 31904 28364 31910 28416
rect 31938 28364 31944 28416
rect 31996 28404 32002 28416
rect 32861 28407 32919 28413
rect 32861 28404 32873 28407
rect 31996 28376 32873 28404
rect 31996 28364 32002 28376
rect 32861 28373 32873 28376
rect 32907 28373 32919 28407
rect 35342 28404 35348 28416
rect 35303 28376 35348 28404
rect 32861 28367 32919 28373
rect 35342 28364 35348 28376
rect 35400 28364 35406 28416
rect 35805 28407 35863 28413
rect 35805 28373 35817 28407
rect 35851 28404 35863 28407
rect 36078 28404 36084 28416
rect 35851 28376 36084 28404
rect 35851 28373 35863 28376
rect 35805 28367 35863 28373
rect 36078 28364 36084 28376
rect 36136 28364 36142 28416
rect 36262 28364 36268 28416
rect 36320 28404 36326 28416
rect 36320 28376 36365 28404
rect 36320 28364 36326 28376
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 15933 28203 15991 28209
rect 15933 28169 15945 28203
rect 15979 28200 15991 28203
rect 16298 28200 16304 28212
rect 15979 28172 16304 28200
rect 15979 28169 15991 28172
rect 15933 28163 15991 28169
rect 16298 28160 16304 28172
rect 16356 28160 16362 28212
rect 16850 28160 16856 28212
rect 16908 28200 16914 28212
rect 17145 28203 17203 28209
rect 17145 28200 17157 28203
rect 16908 28172 17157 28200
rect 16908 28160 16914 28172
rect 17145 28169 17157 28172
rect 17191 28169 17203 28203
rect 17310 28200 17316 28212
rect 17271 28172 17316 28200
rect 17145 28163 17203 28169
rect 17310 28160 17316 28172
rect 17368 28160 17374 28212
rect 20257 28203 20315 28209
rect 20257 28169 20269 28203
rect 20303 28200 20315 28203
rect 20346 28200 20352 28212
rect 20303 28172 20352 28200
rect 20303 28169 20315 28172
rect 20257 28163 20315 28169
rect 20346 28160 20352 28172
rect 20404 28160 20410 28212
rect 25222 28200 25228 28212
rect 21836 28172 25228 28200
rect 9674 28132 9680 28144
rect 7944 28104 9680 28132
rect 7944 28073 7972 28104
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 12894 28092 12900 28144
rect 12952 28132 12958 28144
rect 13446 28132 13452 28144
rect 12952 28104 13452 28132
rect 12952 28092 12958 28104
rect 13446 28092 13452 28104
rect 13504 28132 13510 28144
rect 16942 28132 16948 28144
rect 13504 28104 15792 28132
rect 16903 28104 16948 28132
rect 13504 28092 13510 28104
rect 7929 28067 7987 28073
rect 7929 28033 7941 28067
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 11422 28024 11428 28076
rect 11480 28064 11486 28076
rect 15764 28073 15792 28104
rect 16942 28092 16948 28104
rect 17000 28092 17006 28144
rect 17954 28092 17960 28144
rect 18012 28132 18018 28144
rect 18049 28135 18107 28141
rect 18049 28132 18061 28135
rect 18012 28104 18061 28132
rect 18012 28092 18018 28104
rect 18049 28101 18061 28104
rect 18095 28101 18107 28135
rect 19334 28132 19340 28144
rect 19274 28104 19340 28132
rect 18049 28095 18107 28101
rect 19334 28092 19340 28104
rect 19392 28092 19398 28144
rect 11517 28067 11575 28073
rect 11517 28064 11529 28067
rect 11480 28036 11529 28064
rect 11480 28024 11486 28036
rect 11517 28033 11529 28036
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 20162 28064 20168 28076
rect 19484 28036 20168 28064
rect 19484 28024 19490 28036
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 21836 28073 21864 28172
rect 25222 28160 25228 28172
rect 25280 28160 25286 28212
rect 25498 28160 25504 28212
rect 25556 28200 25562 28212
rect 25869 28203 25927 28209
rect 25869 28200 25881 28203
rect 25556 28172 25881 28200
rect 25556 28160 25562 28172
rect 25869 28169 25881 28172
rect 25915 28169 25927 28203
rect 30374 28200 30380 28212
rect 25869 28163 25927 28169
rect 27356 28172 30380 28200
rect 22094 28092 22100 28144
rect 22152 28132 22158 28144
rect 22152 28104 22197 28132
rect 22152 28092 22158 28104
rect 22370 28092 22376 28144
rect 22428 28132 22434 28144
rect 22428 28104 22586 28132
rect 22428 28092 22434 28104
rect 23842 28092 23848 28144
rect 23900 28132 23906 28144
rect 23900 28104 25360 28132
rect 23900 28092 23906 28104
rect 21821 28067 21879 28073
rect 21821 28033 21833 28067
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 23474 28024 23480 28076
rect 23532 28064 23538 28076
rect 24029 28067 24087 28073
rect 24029 28064 24041 28067
rect 23532 28036 24041 28064
rect 23532 28024 23538 28036
rect 24029 28033 24041 28036
rect 24075 28033 24087 28067
rect 24029 28027 24087 28033
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 8110 27996 8116 28008
rect 8071 27968 8116 27996
rect 8110 27956 8116 27968
rect 8168 27956 8174 28008
rect 8389 27999 8447 28005
rect 8389 27965 8401 27999
rect 8435 27965 8447 27999
rect 12710 27996 12716 28008
rect 12671 27968 12716 27996
rect 8389 27959 8447 27965
rect 3970 27888 3976 27940
rect 4028 27928 4034 27940
rect 8404 27928 8432 27959
rect 12710 27956 12716 27968
rect 12768 27956 12774 28008
rect 12894 27996 12900 28008
rect 12855 27968 12900 27996
rect 12894 27956 12900 27968
rect 12952 27956 12958 28008
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27965 13231 27999
rect 13173 27959 13231 27965
rect 17773 27999 17831 28005
rect 17773 27965 17785 27999
rect 17819 27965 17831 27999
rect 17773 27959 17831 27965
rect 4028 27900 8432 27928
rect 8496 27900 12434 27928
rect 4028 27888 4034 27900
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8496 27860 8524 27900
rect 8352 27832 8524 27860
rect 8352 27820 8358 27832
rect 11146 27820 11152 27872
rect 11204 27860 11210 27872
rect 11701 27863 11759 27869
rect 11701 27860 11713 27863
rect 11204 27832 11713 27860
rect 11204 27820 11210 27832
rect 11701 27829 11713 27832
rect 11747 27829 11759 27863
rect 12406 27860 12434 27900
rect 13188 27860 13216 27959
rect 12406 27832 13216 27860
rect 11701 27823 11759 27829
rect 17034 27820 17040 27872
rect 17092 27860 17098 27872
rect 17129 27863 17187 27869
rect 17129 27860 17141 27863
rect 17092 27832 17141 27860
rect 17092 27820 17098 27832
rect 17129 27829 17141 27832
rect 17175 27829 17187 27863
rect 17788 27860 17816 27959
rect 18046 27956 18052 28008
rect 18104 27996 18110 28008
rect 19242 27996 19248 28008
rect 18104 27968 19248 27996
rect 18104 27956 18110 27968
rect 19242 27956 19248 27968
rect 19300 27996 19306 28008
rect 19521 27999 19579 28005
rect 19521 27996 19533 27999
rect 19300 27968 19533 27996
rect 19300 27956 19306 27968
rect 19521 27965 19533 27968
rect 19567 27965 19579 27999
rect 23566 27996 23572 28008
rect 23527 27968 23572 27996
rect 19521 27959 19579 27965
rect 23566 27956 23572 27968
rect 23624 27956 23630 28008
rect 24228 27928 24256 28027
rect 24302 28024 24308 28076
rect 24360 28064 24366 28076
rect 24486 28064 24492 28076
rect 24360 28036 24405 28064
rect 24447 28036 24492 28064
rect 24360 28024 24366 28036
rect 24486 28024 24492 28036
rect 24544 28024 24550 28076
rect 24578 28024 24584 28076
rect 24636 28064 24642 28076
rect 25222 28064 25228 28076
rect 24636 28036 24681 28064
rect 25183 28036 25228 28064
rect 24636 28024 24642 28036
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25332 28073 25360 28104
rect 25318 28067 25376 28073
rect 25318 28033 25330 28067
rect 25364 28033 25376 28067
rect 25498 28064 25504 28076
rect 25459 28036 25504 28064
rect 25318 28027 25376 28033
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 25731 28067 25789 28073
rect 25731 28033 25743 28067
rect 25777 28064 25789 28067
rect 27356 28064 27384 28172
rect 30374 28160 30380 28172
rect 30432 28160 30438 28212
rect 31202 28160 31208 28212
rect 31260 28200 31266 28212
rect 31938 28200 31944 28212
rect 31260 28172 31944 28200
rect 31260 28160 31266 28172
rect 31938 28160 31944 28172
rect 31996 28160 32002 28212
rect 35342 28160 35348 28212
rect 35400 28200 35406 28212
rect 36081 28203 36139 28209
rect 36081 28200 36093 28203
rect 35400 28172 36093 28200
rect 35400 28160 35406 28172
rect 36081 28169 36093 28172
rect 36127 28169 36139 28203
rect 36081 28163 36139 28169
rect 27433 28135 27491 28141
rect 27433 28101 27445 28135
rect 27479 28132 27491 28135
rect 31386 28132 31392 28144
rect 27479 28104 31392 28132
rect 27479 28101 27491 28104
rect 27433 28095 27491 28101
rect 31386 28092 31392 28104
rect 31444 28132 31450 28144
rect 32769 28135 32827 28141
rect 32769 28132 32781 28135
rect 31444 28104 32781 28132
rect 31444 28092 31450 28104
rect 32769 28101 32781 28104
rect 32815 28101 32827 28135
rect 32769 28095 32827 28101
rect 27614 28064 27620 28076
rect 25777 28036 27384 28064
rect 27575 28036 27620 28064
rect 25777 28033 25789 28036
rect 25731 28027 25789 28033
rect 24946 27956 24952 28008
rect 25004 27996 25010 28008
rect 25608 27996 25636 28027
rect 27614 28024 27620 28036
rect 27672 28024 27678 28076
rect 29733 28067 29791 28073
rect 29733 28033 29745 28067
rect 29779 28064 29791 28067
rect 29822 28064 29828 28076
rect 29779 28036 29828 28064
rect 29779 28033 29791 28036
rect 29733 28027 29791 28033
rect 29822 28024 29828 28036
rect 29880 28024 29886 28076
rect 29914 28024 29920 28076
rect 29972 28064 29978 28076
rect 30929 28067 30987 28073
rect 30929 28064 30941 28067
rect 29972 28036 30941 28064
rect 29972 28024 29978 28036
rect 30929 28033 30941 28036
rect 30975 28033 30987 28067
rect 31110 28064 31116 28076
rect 31071 28036 31116 28064
rect 30929 28027 30987 28033
rect 25004 27968 25636 27996
rect 30009 27999 30067 28005
rect 25004 27956 25010 27968
rect 30009 27965 30021 27999
rect 30055 27965 30067 27999
rect 30009 27959 30067 27965
rect 26234 27928 26240 27940
rect 24228 27900 26240 27928
rect 26234 27888 26240 27900
rect 26292 27888 26298 27940
rect 29638 27888 29644 27940
rect 29696 27928 29702 27940
rect 29917 27931 29975 27937
rect 29917 27928 29929 27931
rect 29696 27900 29929 27928
rect 29696 27888 29702 27900
rect 29917 27897 29929 27900
rect 29963 27897 29975 27931
rect 29917 27891 29975 27897
rect 18046 27860 18052 27872
rect 17788 27832 18052 27860
rect 17129 27823 17187 27829
rect 18046 27820 18052 27832
rect 18104 27820 18110 27872
rect 29822 27860 29828 27872
rect 29783 27832 29828 27860
rect 29822 27820 29828 27832
rect 29880 27820 29886 27872
rect 30024 27860 30052 27959
rect 30944 27928 30972 28027
rect 31110 28024 31116 28036
rect 31168 28024 31174 28076
rect 31205 28067 31263 28073
rect 31205 28033 31217 28067
rect 31251 28033 31263 28067
rect 32214 28064 32220 28076
rect 31205 28027 31263 28033
rect 31312 28036 32220 28064
rect 31018 27956 31024 28008
rect 31076 27996 31082 28008
rect 31220 27996 31248 28027
rect 31076 27968 31248 27996
rect 31076 27956 31082 27968
rect 31312 27928 31340 28036
rect 32214 28024 32220 28036
rect 32272 28024 32278 28076
rect 32306 28024 32312 28076
rect 32364 28064 32370 28076
rect 33597 28067 33655 28073
rect 33597 28064 33609 28067
rect 32364 28036 33609 28064
rect 32364 28024 32370 28036
rect 33597 28033 33609 28036
rect 33643 28033 33655 28067
rect 35986 28064 35992 28076
rect 35947 28036 35992 28064
rect 33597 28027 33655 28033
rect 35986 28024 35992 28036
rect 36044 28024 36050 28076
rect 36078 28024 36084 28076
rect 36136 28064 36142 28076
rect 37461 28067 37519 28073
rect 37461 28064 37473 28067
rect 36136 28036 37473 28064
rect 36136 28024 36142 28036
rect 37461 28033 37473 28036
rect 37507 28033 37519 28067
rect 37461 28027 37519 28033
rect 37734 28024 37740 28076
rect 37792 28064 37798 28076
rect 37921 28067 37979 28073
rect 37921 28064 37933 28067
rect 37792 28036 37933 28064
rect 37792 28024 37798 28036
rect 37921 28033 37933 28036
rect 37967 28033 37979 28067
rect 37921 28027 37979 28033
rect 46566 28024 46572 28076
rect 46624 28064 46630 28076
rect 47578 28064 47584 28076
rect 46624 28036 47584 28064
rect 46624 28024 46630 28036
rect 47578 28024 47584 28036
rect 47636 28024 47642 28076
rect 31570 27956 31576 28008
rect 31628 27996 31634 28008
rect 35802 27996 35808 28008
rect 31628 27968 35808 27996
rect 31628 27956 31634 27968
rect 35802 27956 35808 27968
rect 35860 27956 35866 28008
rect 36170 27996 36176 28008
rect 36083 27968 36176 27996
rect 36170 27956 36176 27968
rect 36228 27996 36234 28008
rect 36354 27996 36360 28008
rect 36228 27968 36360 27996
rect 36228 27956 36234 27968
rect 36354 27956 36360 27968
rect 36412 27956 36418 28008
rect 30944 27900 31340 27928
rect 32953 27931 33011 27937
rect 32953 27897 32965 27931
rect 32999 27928 33011 27931
rect 33502 27928 33508 27940
rect 32999 27900 33508 27928
rect 32999 27897 33011 27900
rect 32953 27891 33011 27897
rect 33502 27888 33508 27900
rect 33560 27888 33566 27940
rect 35621 27931 35679 27937
rect 35621 27897 35633 27931
rect 35667 27928 35679 27931
rect 36262 27928 36268 27940
rect 35667 27900 36268 27928
rect 35667 27897 35679 27900
rect 35621 27891 35679 27897
rect 36262 27888 36268 27900
rect 36320 27888 36326 27940
rect 31018 27860 31024 27872
rect 30024 27832 31024 27860
rect 31018 27820 31024 27832
rect 31076 27820 31082 27872
rect 31202 27860 31208 27872
rect 31163 27832 31208 27860
rect 31202 27820 31208 27832
rect 31260 27820 31266 27872
rect 31294 27820 31300 27872
rect 31352 27860 31358 27872
rect 31389 27863 31447 27869
rect 31389 27860 31401 27863
rect 31352 27832 31401 27860
rect 31352 27820 31358 27832
rect 31389 27829 31401 27832
rect 31435 27829 31447 27863
rect 33410 27860 33416 27872
rect 33371 27832 33416 27860
rect 31389 27823 31447 27829
rect 33410 27820 33416 27832
rect 33468 27820 33474 27872
rect 36354 27820 36360 27872
rect 36412 27860 36418 27872
rect 37277 27863 37335 27869
rect 37277 27860 37289 27863
rect 36412 27832 37289 27860
rect 36412 27820 36418 27832
rect 37277 27829 37289 27832
rect 37323 27829 37335 27863
rect 38010 27860 38016 27872
rect 37971 27832 38016 27860
rect 37277 27823 37335 27829
rect 38010 27820 38016 27832
rect 38068 27820 38074 27872
rect 47026 27860 47032 27872
rect 46987 27832 47032 27860
rect 47026 27820 47032 27832
rect 47084 27820 47090 27872
rect 47670 27860 47676 27872
rect 47631 27832 47676 27860
rect 47670 27820 47676 27832
rect 47728 27820 47734 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 7653 27659 7711 27665
rect 7653 27625 7665 27659
rect 7699 27656 7711 27659
rect 8110 27656 8116 27668
rect 7699 27628 8116 27656
rect 7699 27625 7711 27628
rect 7653 27619 7711 27625
rect 8110 27616 8116 27628
rect 8168 27616 8174 27668
rect 12894 27616 12900 27668
rect 12952 27656 12958 27668
rect 13173 27659 13231 27665
rect 13173 27656 13185 27659
rect 12952 27628 13185 27656
rect 12952 27616 12958 27628
rect 13173 27625 13185 27628
rect 13219 27625 13231 27659
rect 17954 27656 17960 27668
rect 13173 27619 13231 27625
rect 17880 27628 17960 27656
rect 9030 27588 9036 27600
rect 8991 27560 9036 27588
rect 9030 27548 9036 27560
rect 9088 27548 9094 27600
rect 9674 27588 9680 27600
rect 9232 27560 9680 27588
rect 9232 27529 9260 27560
rect 9674 27548 9680 27560
rect 9732 27588 9738 27600
rect 10137 27591 10195 27597
rect 10137 27588 10149 27591
rect 9732 27560 10149 27588
rect 9732 27548 9738 27560
rect 10137 27557 10149 27560
rect 10183 27588 10195 27591
rect 10686 27588 10692 27600
rect 10183 27560 10692 27588
rect 10183 27557 10195 27560
rect 10137 27551 10195 27557
rect 10686 27548 10692 27560
rect 10744 27548 10750 27600
rect 17221 27591 17279 27597
rect 17221 27557 17233 27591
rect 17267 27588 17279 27591
rect 17880 27588 17908 27628
rect 17954 27616 17960 27628
rect 18012 27616 18018 27668
rect 23569 27659 23627 27665
rect 23569 27625 23581 27659
rect 23615 27656 23627 27659
rect 25406 27656 25412 27668
rect 23615 27628 25412 27656
rect 23615 27625 23627 27628
rect 23569 27619 23627 27625
rect 25406 27616 25412 27628
rect 25464 27616 25470 27668
rect 25498 27616 25504 27668
rect 25556 27656 25562 27668
rect 27890 27656 27896 27668
rect 25556 27628 27896 27656
rect 25556 27616 25562 27628
rect 27890 27616 27896 27628
rect 27948 27656 27954 27668
rect 27948 27628 30972 27656
rect 27948 27616 27954 27628
rect 18046 27588 18052 27600
rect 17267 27560 17908 27588
rect 18007 27560 18052 27588
rect 17267 27557 17279 27560
rect 17221 27551 17279 27557
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 19334 27588 19340 27600
rect 19295 27560 19340 27588
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 23658 27588 23664 27600
rect 23492 27560 23664 27588
rect 9217 27523 9275 27529
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9217 27483 9275 27489
rect 9309 27523 9367 27529
rect 9309 27489 9321 27523
rect 9355 27520 9367 27523
rect 9582 27520 9588 27532
rect 9355 27492 9588 27520
rect 9355 27489 9367 27492
rect 9309 27483 9367 27489
rect 9582 27480 9588 27492
rect 9640 27520 9646 27532
rect 23492 27529 23520 27560
rect 23658 27548 23664 27560
rect 23716 27548 23722 27600
rect 23750 27548 23756 27600
rect 23808 27588 23814 27600
rect 23845 27591 23903 27597
rect 23845 27588 23857 27591
rect 23808 27560 23857 27588
rect 23808 27548 23814 27560
rect 23845 27557 23857 27560
rect 23891 27557 23903 27591
rect 23845 27551 23903 27557
rect 24670 27548 24676 27600
rect 24728 27588 24734 27600
rect 24949 27591 25007 27597
rect 24949 27588 24961 27591
rect 24728 27560 24961 27588
rect 24728 27548 24734 27560
rect 24949 27557 24961 27560
rect 24995 27588 25007 27591
rect 24995 27560 27108 27588
rect 24995 27557 25007 27560
rect 24949 27551 25007 27557
rect 23477 27523 23535 27529
rect 23477 27520 23489 27523
rect 9640 27492 10364 27520
rect 9640 27480 9646 27492
rect 7558 27452 7564 27464
rect 7519 27424 7564 27452
rect 7558 27412 7564 27424
rect 7616 27412 7622 27464
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8846 27452 8852 27464
rect 8435 27424 8852 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8846 27412 8852 27424
rect 8904 27452 8910 27464
rect 9677 27455 9735 27461
rect 8904 27446 9536 27452
rect 8904 27424 9628 27446
rect 8904 27412 8910 27424
rect 9508 27418 9628 27424
rect 9600 27384 9628 27418
rect 9677 27421 9689 27455
rect 9723 27452 9735 27455
rect 10042 27452 10048 27464
rect 9723 27424 10048 27452
rect 9723 27421 9735 27424
rect 9677 27415 9735 27421
rect 10042 27412 10048 27424
rect 10100 27412 10106 27464
rect 10336 27461 10364 27492
rect 22756 27492 23489 27520
rect 10321 27455 10379 27461
rect 10321 27421 10333 27455
rect 10367 27421 10379 27455
rect 11146 27452 11152 27464
rect 11107 27424 11152 27452
rect 10321 27415 10379 27421
rect 11146 27412 11152 27424
rect 11204 27412 11210 27464
rect 12618 27412 12624 27464
rect 12676 27452 12682 27464
rect 13078 27452 13084 27464
rect 12676 27424 13084 27452
rect 12676 27412 12682 27424
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 17402 27452 17408 27464
rect 17363 27424 17408 27452
rect 17402 27412 17408 27424
rect 17460 27412 17466 27464
rect 18046 27452 18052 27464
rect 18007 27424 18052 27452
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 19150 27412 19156 27464
rect 19208 27452 19214 27464
rect 22756 27461 22784 27492
rect 23477 27489 23489 27492
rect 23523 27489 23535 27523
rect 24486 27520 24492 27532
rect 23477 27483 23535 27489
rect 23584 27492 24492 27520
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 19208 27424 19257 27452
rect 19208 27412 19214 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 22741 27455 22799 27461
rect 22741 27421 22753 27455
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23584 27452 23612 27492
rect 24486 27480 24492 27492
rect 24544 27480 24550 27532
rect 22971 27424 23612 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23658 27412 23664 27464
rect 23716 27452 23722 27464
rect 24762 27452 24768 27464
rect 23716 27424 23761 27452
rect 24723 27424 24768 27452
rect 23716 27412 23722 27424
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 26237 27455 26295 27461
rect 26237 27421 26249 27455
rect 26283 27452 26295 27455
rect 26326 27452 26332 27464
rect 26283 27424 26332 27452
rect 26283 27421 26295 27424
rect 26237 27415 26295 27421
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 27080 27452 27108 27560
rect 30944 27520 30972 27628
rect 31018 27616 31024 27668
rect 31076 27656 31082 27668
rect 36354 27665 36360 27668
rect 32125 27659 32183 27665
rect 32125 27656 32137 27659
rect 31076 27628 32137 27656
rect 31076 27616 31082 27628
rect 32125 27625 32137 27628
rect 32171 27625 32183 27659
rect 32125 27619 32183 27625
rect 36344 27659 36360 27665
rect 36344 27625 36356 27659
rect 36344 27619 36360 27625
rect 36354 27616 36360 27619
rect 36412 27616 36418 27668
rect 31386 27588 31392 27600
rect 31347 27560 31392 27588
rect 31386 27548 31392 27560
rect 31444 27548 31450 27600
rect 31478 27548 31484 27600
rect 31536 27588 31542 27600
rect 32585 27591 32643 27597
rect 32585 27588 32597 27591
rect 31536 27560 32597 27588
rect 31536 27548 31542 27560
rect 32585 27557 32597 27560
rect 32631 27557 32643 27591
rect 32585 27551 32643 27557
rect 34790 27548 34796 27600
rect 34848 27588 34854 27600
rect 34885 27591 34943 27597
rect 34885 27588 34897 27591
rect 34848 27560 34897 27588
rect 34848 27548 34854 27560
rect 34885 27557 34897 27560
rect 34931 27557 34943 27591
rect 34885 27551 34943 27557
rect 41414 27548 41420 27600
rect 41472 27588 41478 27600
rect 42058 27588 42064 27600
rect 41472 27560 42064 27588
rect 41472 27548 41478 27560
rect 42058 27548 42064 27560
rect 42116 27548 42122 27600
rect 31570 27520 31576 27532
rect 30944 27492 31576 27520
rect 31570 27480 31576 27492
rect 31628 27480 31634 27532
rect 32214 27520 32220 27532
rect 32175 27492 32220 27520
rect 32214 27480 32220 27492
rect 32272 27480 32278 27532
rect 32324 27492 33640 27520
rect 32324 27452 32352 27492
rect 27080 27424 32352 27452
rect 32401 27455 32459 27461
rect 32401 27421 32413 27455
rect 32447 27452 32459 27455
rect 32582 27452 32588 27464
rect 32447 27424 32588 27452
rect 32447 27421 32459 27424
rect 32401 27415 32459 27421
rect 32582 27412 32588 27424
rect 32640 27412 32646 27464
rect 33612 27461 33640 27492
rect 33778 27480 33784 27532
rect 33836 27520 33842 27532
rect 36081 27523 36139 27529
rect 36081 27520 36093 27523
rect 33836 27492 36093 27520
rect 33836 27480 33842 27492
rect 36081 27489 36093 27492
rect 36127 27489 36139 27523
rect 36081 27483 36139 27489
rect 36446 27480 36452 27532
rect 36504 27520 36510 27532
rect 37829 27523 37887 27529
rect 37829 27520 37841 27523
rect 36504 27492 37841 27520
rect 36504 27480 36510 27492
rect 37829 27489 37841 27492
rect 37875 27489 37887 27523
rect 37829 27483 37887 27489
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27520 46351 27523
rect 47026 27520 47032 27532
rect 46339 27492 47032 27520
rect 46339 27489 46351 27492
rect 46293 27483 46351 27489
rect 47026 27480 47032 27492
rect 47084 27480 47090 27532
rect 48130 27520 48136 27532
rect 48091 27492 48136 27520
rect 48130 27480 48136 27492
rect 48188 27480 48194 27532
rect 33597 27455 33655 27461
rect 33060 27424 33364 27452
rect 10505 27387 10563 27393
rect 10505 27384 10517 27387
rect 8220 27356 9536 27384
rect 9600 27356 10517 27384
rect 8220 27328 8248 27356
rect 8202 27316 8208 27328
rect 8163 27288 8208 27316
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 9214 27276 9220 27328
rect 9272 27316 9278 27328
rect 9401 27319 9459 27325
rect 9401 27316 9413 27319
rect 9272 27288 9413 27316
rect 9272 27276 9278 27288
rect 9401 27285 9413 27288
rect 9447 27285 9459 27319
rect 9508 27316 9536 27356
rect 10505 27353 10517 27356
rect 10551 27353 10563 27387
rect 10505 27347 10563 27353
rect 22833 27387 22891 27393
rect 22833 27353 22845 27387
rect 22879 27384 22891 27387
rect 23385 27387 23443 27393
rect 23385 27384 23397 27387
rect 22879 27356 23397 27384
rect 22879 27353 22891 27356
rect 22833 27347 22891 27353
rect 23385 27353 23397 27356
rect 23431 27384 23443 27387
rect 24302 27384 24308 27396
rect 23431 27356 24308 27384
rect 23431 27353 23443 27356
rect 23385 27347 23443 27353
rect 24302 27344 24308 27356
rect 24360 27344 24366 27396
rect 29914 27384 29920 27396
rect 29875 27356 29920 27384
rect 29914 27344 29920 27356
rect 29972 27344 29978 27396
rect 32030 27344 32036 27396
rect 32088 27384 32094 27396
rect 32125 27387 32183 27393
rect 32125 27384 32137 27387
rect 32088 27356 32137 27384
rect 32088 27344 32094 27356
rect 32125 27353 32137 27356
rect 32171 27353 32183 27387
rect 32125 27347 32183 27353
rect 9585 27319 9643 27325
rect 9585 27316 9597 27319
rect 9508 27288 9597 27316
rect 9401 27279 9459 27285
rect 9585 27285 9597 27288
rect 9631 27285 9643 27319
rect 9585 27279 9643 27285
rect 10226 27276 10232 27328
rect 10284 27316 10290 27328
rect 10413 27319 10471 27325
rect 10413 27316 10425 27319
rect 10284 27288 10425 27316
rect 10284 27276 10290 27288
rect 10413 27285 10425 27288
rect 10459 27285 10471 27319
rect 10413 27279 10471 27285
rect 10689 27319 10747 27325
rect 10689 27285 10701 27319
rect 10735 27316 10747 27319
rect 11238 27316 11244 27328
rect 10735 27288 11244 27316
rect 10735 27285 10747 27288
rect 10689 27279 10747 27285
rect 11238 27276 11244 27288
rect 11296 27276 11302 27328
rect 11333 27319 11391 27325
rect 11333 27285 11345 27319
rect 11379 27316 11391 27319
rect 11514 27316 11520 27328
rect 11379 27288 11520 27316
rect 11379 27285 11391 27288
rect 11333 27279 11391 27285
rect 11514 27276 11520 27288
rect 11572 27276 11578 27328
rect 26329 27319 26387 27325
rect 26329 27285 26341 27319
rect 26375 27316 26387 27319
rect 26418 27316 26424 27328
rect 26375 27288 26424 27316
rect 26375 27285 26387 27288
rect 26329 27279 26387 27285
rect 26418 27276 26424 27288
rect 26476 27276 26482 27328
rect 30190 27276 30196 27328
rect 30248 27316 30254 27328
rect 33060 27316 33088 27424
rect 33336 27384 33364 27424
rect 33597 27421 33609 27455
rect 33643 27452 33655 27455
rect 33962 27452 33968 27464
rect 33643 27424 33968 27452
rect 33643 27421 33655 27424
rect 33597 27415 33655 27421
rect 33962 27412 33968 27424
rect 34020 27452 34026 27464
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 34020 27424 34713 27452
rect 34020 27412 34026 27424
rect 34701 27421 34713 27424
rect 34747 27421 34759 27455
rect 34701 27415 34759 27421
rect 37734 27412 37740 27464
rect 37792 27452 37798 27464
rect 38289 27455 38347 27461
rect 38289 27452 38301 27455
rect 37792 27424 38301 27452
rect 37792 27412 37798 27424
rect 38289 27421 38301 27424
rect 38335 27421 38347 27455
rect 38289 27415 38347 27421
rect 35434 27384 35440 27396
rect 33336 27356 35440 27384
rect 35434 27344 35440 27356
rect 35492 27344 35498 27396
rect 38010 27384 38016 27396
rect 37582 27356 38016 27384
rect 38010 27344 38016 27356
rect 38068 27344 38074 27396
rect 46477 27387 46535 27393
rect 46477 27353 46489 27387
rect 46523 27384 46535 27387
rect 47670 27384 47676 27396
rect 46523 27356 47676 27384
rect 46523 27353 46535 27356
rect 46477 27347 46535 27353
rect 47670 27344 47676 27356
rect 47728 27344 47734 27396
rect 30248 27288 33088 27316
rect 30248 27276 30254 27288
rect 33318 27276 33324 27328
rect 33376 27316 33382 27328
rect 33686 27316 33692 27328
rect 33376 27288 33692 27316
rect 33376 27276 33382 27288
rect 33686 27276 33692 27288
rect 33744 27316 33750 27328
rect 33781 27319 33839 27325
rect 33781 27316 33793 27319
rect 33744 27288 33793 27316
rect 33744 27276 33750 27288
rect 33781 27285 33793 27288
rect 33827 27285 33839 27319
rect 38378 27316 38384 27328
rect 38339 27288 38384 27316
rect 33781 27279 33839 27285
rect 38378 27276 38384 27288
rect 38436 27276 38442 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 7558 27072 7564 27124
rect 7616 27112 7622 27124
rect 8018 27112 8024 27124
rect 7616 27084 8024 27112
rect 7616 27072 7622 27084
rect 8018 27072 8024 27084
rect 8076 27112 8082 27124
rect 12526 27112 12532 27124
rect 8076 27084 12532 27112
rect 8076 27072 8082 27084
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 13265 27115 13323 27121
rect 13265 27112 13277 27115
rect 12768 27084 13277 27112
rect 12768 27072 12774 27084
rect 13265 27081 13277 27084
rect 13311 27081 13323 27115
rect 27890 27112 27896 27124
rect 27851 27084 27896 27112
rect 13265 27075 13323 27081
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 29549 27115 29607 27121
rect 29549 27081 29561 27115
rect 29595 27112 29607 27115
rect 31294 27112 31300 27124
rect 29595 27084 31300 27112
rect 29595 27081 29607 27084
rect 29549 27075 29607 27081
rect 31294 27072 31300 27084
rect 31352 27072 31358 27124
rect 33410 27112 33416 27124
rect 32508 27084 33416 27112
rect 8389 27047 8447 27053
rect 8389 27013 8401 27047
rect 8435 27044 8447 27047
rect 9030 27044 9036 27056
rect 8435 27016 9036 27044
rect 8435 27013 8447 27016
rect 8389 27007 8447 27013
rect 9030 27004 9036 27016
rect 9088 27044 9094 27056
rect 9217 27047 9275 27053
rect 9217 27044 9229 27047
rect 9088 27016 9229 27044
rect 9088 27004 9094 27016
rect 9217 27013 9229 27016
rect 9263 27044 9275 27047
rect 9263 27016 10364 27044
rect 9263 27013 9275 27016
rect 9217 27007 9275 27013
rect 8202 26936 8208 26988
rect 8260 26976 8266 26988
rect 9122 26976 9128 26988
rect 8260 26948 9128 26976
rect 8260 26936 8266 26948
rect 9122 26936 9128 26948
rect 9180 26976 9186 26988
rect 9401 26979 9459 26985
rect 9401 26976 9413 26979
rect 9180 26948 9413 26976
rect 9180 26936 9186 26948
rect 9401 26945 9413 26948
rect 9447 26945 9459 26979
rect 9401 26939 9459 26945
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26976 9551 26979
rect 10226 26976 10232 26988
rect 9539 26948 10232 26976
rect 9539 26945 9551 26948
rect 9493 26939 9551 26945
rect 8021 26843 8079 26849
rect 8021 26809 8033 26843
rect 8067 26840 8079 26843
rect 8294 26840 8300 26852
rect 8067 26812 8300 26840
rect 8067 26809 8079 26812
rect 8021 26803 8079 26809
rect 8294 26800 8300 26812
rect 8352 26800 8358 26852
rect 9214 26800 9220 26852
rect 9272 26840 9278 26852
rect 9508 26840 9536 26939
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 10336 26985 10364 27016
rect 12250 27004 12256 27056
rect 12308 27004 12314 27056
rect 13078 27004 13084 27056
rect 13136 27044 13142 27056
rect 17221 27047 17279 27053
rect 13136 27016 17172 27044
rect 13136 27004 13142 27016
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26945 10379 26979
rect 11514 26976 11520 26988
rect 11475 26948 11520 26976
rect 10321 26939 10379 26945
rect 11514 26936 11520 26948
rect 11572 26936 11578 26988
rect 17144 26985 17172 27016
rect 17221 27013 17233 27047
rect 17267 27044 17279 27047
rect 17957 27047 18015 27053
rect 17957 27044 17969 27047
rect 17267 27016 17969 27044
rect 17267 27013 17279 27016
rect 17221 27007 17279 27013
rect 17957 27013 17969 27016
rect 18003 27013 18015 27047
rect 17957 27007 18015 27013
rect 18138 27004 18144 27056
rect 18196 27044 18202 27056
rect 23566 27044 23572 27056
rect 18196 27016 23572 27044
rect 18196 27004 18202 27016
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 30190 27044 30196 27056
rect 24872 27016 29316 27044
rect 30151 27016 30196 27044
rect 24872 26988 24900 27016
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26976 17187 26979
rect 17586 26976 17592 26988
rect 17175 26948 17592 26976
rect 17175 26945 17187 26948
rect 17129 26939 17187 26945
rect 10042 26908 10048 26920
rect 9955 26880 10048 26908
rect 10042 26868 10048 26880
rect 10100 26868 10106 26920
rect 11790 26908 11796 26920
rect 11751 26880 11796 26908
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 12526 26868 12532 26920
rect 12584 26908 12590 26920
rect 14936 26908 14964 26939
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 17678 26936 17684 26988
rect 17736 26976 17742 26988
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 17736 26948 17785 26976
rect 17736 26936 17742 26948
rect 17773 26945 17785 26948
rect 17819 26945 17831 26979
rect 20073 26979 20131 26985
rect 20073 26976 20085 26979
rect 17773 26939 17831 26945
rect 19168 26948 20085 26976
rect 17034 26908 17040 26920
rect 12584 26880 17040 26908
rect 12584 26868 12590 26880
rect 17034 26868 17040 26880
rect 17092 26868 17098 26920
rect 17604 26908 17632 26936
rect 19168 26908 19196 26948
rect 20073 26945 20085 26948
rect 20119 26945 20131 26979
rect 22554 26976 22560 26988
rect 22515 26948 22560 26976
rect 20073 26939 20131 26945
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 23474 26976 23480 26988
rect 23435 26948 23480 26976
rect 23474 26936 23480 26948
rect 23532 26936 23538 26988
rect 24118 26976 24124 26988
rect 24079 26948 24124 26976
rect 24118 26936 24124 26948
rect 24176 26936 24182 26988
rect 24854 26976 24860 26988
rect 24767 26948 24860 26976
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 27154 26976 27160 26988
rect 27115 26948 27160 26976
rect 27154 26936 27160 26948
rect 27212 26936 27218 26988
rect 27709 26979 27767 26985
rect 27709 26945 27721 26979
rect 27755 26976 27767 26979
rect 27798 26976 27804 26988
rect 27755 26948 27804 26976
rect 27755 26945 27767 26948
rect 27709 26939 27767 26945
rect 27798 26936 27804 26948
rect 27856 26936 27862 26988
rect 17604 26880 19196 26908
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26908 19671 26911
rect 20254 26908 20260 26920
rect 19659 26880 20260 26908
rect 19659 26877 19671 26880
rect 19613 26871 19671 26877
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 21082 26868 21088 26920
rect 21140 26908 21146 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 21140 26880 22845 26908
rect 21140 26868 21146 26880
rect 22833 26877 22845 26880
rect 22879 26908 22891 26911
rect 23106 26908 23112 26920
rect 22879 26880 23112 26908
rect 22879 26877 22891 26880
rect 22833 26871 22891 26877
rect 23106 26868 23112 26880
rect 23164 26908 23170 26920
rect 23658 26908 23664 26920
rect 23164 26880 23664 26908
rect 23164 26868 23170 26880
rect 23658 26868 23664 26880
rect 23716 26908 23722 26920
rect 24949 26911 25007 26917
rect 24949 26908 24961 26911
rect 23716 26880 24961 26908
rect 23716 26868 23722 26880
rect 24949 26877 24961 26880
rect 24995 26877 25007 26911
rect 29178 26908 29184 26920
rect 29139 26880 29184 26908
rect 24949 26871 25007 26877
rect 29178 26868 29184 26880
rect 29236 26868 29242 26920
rect 29288 26908 29316 27016
rect 30190 27004 30196 27016
rect 30248 27004 30254 27056
rect 30374 27044 30380 27056
rect 30335 27016 30380 27044
rect 30374 27004 30380 27016
rect 30432 27004 30438 27056
rect 32508 27053 32536 27084
rect 33410 27072 33416 27084
rect 33468 27072 33474 27124
rect 32493 27047 32551 27053
rect 32493 27013 32505 27047
rect 32539 27013 32551 27047
rect 33778 27044 33784 27056
rect 33718 27016 33784 27044
rect 32493 27007 32551 27013
rect 33778 27004 33784 27016
rect 33836 27004 33842 27056
rect 29638 26936 29644 26988
rect 29696 26976 29702 26988
rect 29696 26948 29741 26976
rect 29696 26936 29702 26948
rect 33870 26936 33876 26988
rect 33928 26976 33934 26988
rect 34701 26979 34759 26985
rect 34701 26976 34713 26979
rect 33928 26948 34713 26976
rect 33928 26936 33934 26948
rect 34701 26945 34713 26948
rect 34747 26945 34759 26979
rect 34701 26939 34759 26945
rect 38286 26936 38292 26988
rect 38344 26976 38350 26988
rect 38381 26979 38439 26985
rect 38381 26976 38393 26979
rect 38344 26948 38393 26976
rect 38344 26936 38350 26948
rect 38381 26945 38393 26948
rect 38427 26945 38439 26979
rect 38381 26939 38439 26945
rect 38565 26979 38623 26985
rect 38565 26945 38577 26979
rect 38611 26976 38623 26979
rect 44266 26976 44272 26988
rect 38611 26948 44272 26976
rect 38611 26945 38623 26948
rect 38565 26939 38623 26945
rect 44266 26936 44272 26948
rect 44324 26936 44330 26988
rect 31938 26908 31944 26920
rect 29288 26880 31944 26908
rect 31938 26868 31944 26880
rect 31996 26868 32002 26920
rect 32217 26911 32275 26917
rect 32217 26877 32229 26911
rect 32263 26877 32275 26911
rect 32217 26871 32275 26877
rect 9272 26812 9536 26840
rect 9272 26800 9278 26812
rect 7374 26732 7380 26784
rect 7432 26772 7438 26784
rect 8202 26772 8208 26784
rect 7432 26744 8208 26772
rect 7432 26732 7438 26744
rect 8202 26732 8208 26744
rect 8260 26772 8266 26784
rect 8389 26775 8447 26781
rect 8389 26772 8401 26775
rect 8260 26744 8401 26772
rect 8260 26732 8266 26744
rect 8389 26741 8401 26744
rect 8435 26741 8447 26775
rect 8570 26772 8576 26784
rect 8531 26744 8576 26772
rect 8389 26735 8447 26741
rect 8570 26732 8576 26744
rect 8628 26732 8634 26784
rect 9490 26772 9496 26784
rect 9451 26744 9496 26772
rect 9490 26732 9496 26744
rect 9548 26732 9554 26784
rect 10060 26772 10088 26868
rect 17862 26800 17868 26852
rect 17920 26840 17926 26852
rect 32122 26840 32128 26852
rect 17920 26812 32128 26840
rect 17920 26800 17926 26812
rect 32122 26800 32128 26812
rect 32180 26800 32186 26852
rect 12342 26772 12348 26784
rect 10060 26744 12348 26772
rect 12342 26732 12348 26744
rect 12400 26732 12406 26784
rect 15010 26772 15016 26784
rect 14971 26744 15016 26772
rect 15010 26732 15016 26744
rect 15068 26732 15074 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 20165 26775 20223 26781
rect 20165 26772 20177 26775
rect 19484 26744 20177 26772
rect 19484 26732 19490 26744
rect 20165 26741 20177 26744
rect 20211 26741 20223 26775
rect 20165 26735 20223 26741
rect 22373 26775 22431 26781
rect 22373 26741 22385 26775
rect 22419 26772 22431 26775
rect 22646 26772 22652 26784
rect 22419 26744 22652 26772
rect 22419 26741 22431 26744
rect 22373 26735 22431 26741
rect 22646 26732 22652 26744
rect 22704 26732 22710 26784
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23566 26772 23572 26784
rect 22796 26744 22841 26772
rect 23527 26744 23572 26772
rect 22796 26732 22802 26744
rect 23566 26732 23572 26744
rect 23624 26732 23630 26784
rect 24302 26772 24308 26784
rect 24263 26744 24308 26772
rect 24302 26732 24308 26744
rect 24360 26732 24366 26784
rect 25958 26732 25964 26784
rect 26016 26772 26022 26784
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26016 26744 26985 26772
rect 26016 26732 26022 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 26973 26735 27031 26741
rect 28994 26732 29000 26784
rect 29052 26772 29058 26784
rect 29365 26775 29423 26781
rect 29365 26772 29377 26775
rect 29052 26744 29377 26772
rect 29052 26732 29058 26744
rect 29365 26741 29377 26744
rect 29411 26741 29423 26775
rect 32232 26772 32260 26871
rect 32582 26868 32588 26920
rect 32640 26908 32646 26920
rect 33965 26911 34023 26917
rect 33965 26908 33977 26911
rect 32640 26880 33977 26908
rect 32640 26868 32646 26880
rect 33965 26877 33977 26880
rect 34011 26877 34023 26911
rect 33965 26871 34023 26877
rect 33594 26800 33600 26852
rect 33652 26840 33658 26852
rect 37734 26840 37740 26852
rect 33652 26812 37740 26840
rect 33652 26800 33658 26812
rect 37734 26800 37740 26812
rect 37792 26800 37798 26852
rect 33042 26772 33048 26784
rect 32232 26744 33048 26772
rect 29365 26735 29423 26741
rect 33042 26732 33048 26744
rect 33100 26732 33106 26784
rect 34790 26772 34796 26784
rect 34751 26744 34796 26772
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 38654 26732 38660 26784
rect 38712 26772 38718 26784
rect 38749 26775 38807 26781
rect 38749 26772 38761 26775
rect 38712 26744 38761 26772
rect 38712 26732 38718 26744
rect 38749 26741 38761 26744
rect 38795 26741 38807 26775
rect 38749 26735 38807 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 8386 26528 8392 26580
rect 8444 26568 8450 26580
rect 9490 26568 9496 26580
rect 8444 26540 9496 26568
rect 8444 26528 8450 26540
rect 9490 26528 9496 26540
rect 9548 26528 9554 26580
rect 12250 26568 12256 26580
rect 12211 26540 12256 26568
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 12400 26540 17141 26568
rect 12400 26528 12406 26540
rect 17129 26537 17141 26540
rect 17175 26537 17187 26571
rect 17129 26531 17187 26537
rect 17586 26528 17592 26580
rect 17644 26568 17650 26580
rect 18417 26571 18475 26577
rect 18417 26568 18429 26571
rect 17644 26540 18429 26568
rect 17644 26528 17650 26540
rect 18417 26537 18429 26540
rect 18463 26537 18475 26571
rect 18417 26531 18475 26537
rect 22554 26528 22560 26580
rect 22612 26568 22618 26580
rect 22830 26568 22836 26580
rect 22612 26540 22836 26568
rect 22612 26528 22618 26540
rect 22830 26528 22836 26540
rect 22888 26568 22894 26580
rect 23293 26571 23351 26577
rect 23293 26568 23305 26571
rect 22888 26540 23305 26568
rect 22888 26528 22894 26540
rect 23293 26537 23305 26540
rect 23339 26537 23351 26571
rect 23293 26531 23351 26537
rect 24302 26528 24308 26580
rect 24360 26568 24366 26580
rect 24360 26540 31432 26568
rect 24360 26528 24366 26540
rect 9030 26500 9036 26512
rect 7208 26472 9036 26500
rect 7208 26373 7236 26472
rect 9030 26460 9036 26472
rect 9088 26500 9094 26512
rect 11241 26503 11299 26509
rect 9088 26472 10916 26500
rect 9088 26460 9094 26472
rect 8570 26432 8576 26444
rect 8036 26404 8576 26432
rect 7193 26367 7251 26373
rect 7193 26333 7205 26367
rect 7239 26333 7251 26367
rect 7374 26364 7380 26376
rect 7335 26336 7380 26364
rect 7193 26327 7251 26333
rect 7374 26324 7380 26336
rect 7432 26324 7438 26376
rect 8036 26373 8064 26404
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 10888 26441 10916 26472
rect 11241 26469 11253 26503
rect 11287 26500 11299 26503
rect 12805 26503 12863 26509
rect 12805 26500 12817 26503
rect 11287 26472 12817 26500
rect 11287 26469 11299 26472
rect 11241 26463 11299 26469
rect 12805 26469 12817 26472
rect 12851 26469 12863 26503
rect 12805 26463 12863 26469
rect 15838 26460 15844 26512
rect 15896 26500 15902 26512
rect 15896 26472 17816 26500
rect 15896 26460 15902 26472
rect 9309 26435 9367 26441
rect 9309 26401 9321 26435
rect 9355 26432 9367 26435
rect 10873 26435 10931 26441
rect 9355 26404 9996 26432
rect 9355 26401 9367 26404
rect 9309 26395 9367 26401
rect 8021 26367 8079 26373
rect 8021 26333 8033 26367
rect 8067 26333 8079 26367
rect 8021 26327 8079 26333
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26364 8355 26367
rect 8386 26364 8392 26376
rect 8343 26336 8392 26364
rect 8343 26333 8355 26336
rect 8297 26327 8355 26333
rect 7285 26299 7343 26305
rect 7285 26265 7297 26299
rect 7331 26296 7343 26299
rect 8312 26296 8340 26327
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9490 26324 9496 26376
rect 9548 26364 9554 26376
rect 9968 26373 9996 26404
rect 10873 26401 10885 26435
rect 10919 26401 10931 26435
rect 10873 26395 10931 26401
rect 12710 26392 12716 26444
rect 12768 26432 12774 26444
rect 12989 26435 13047 26441
rect 12989 26432 13001 26435
rect 12768 26404 13001 26432
rect 12768 26392 12774 26404
rect 12989 26401 13001 26404
rect 13035 26401 13047 26435
rect 15010 26432 15016 26444
rect 14971 26404 15016 26432
rect 12989 26395 13047 26401
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 16482 26432 16488 26444
rect 16443 26404 16488 26432
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 17512 26404 17724 26432
rect 9769 26367 9827 26373
rect 9769 26364 9781 26367
rect 9548 26336 9781 26364
rect 9548 26324 9554 26336
rect 9769 26333 9781 26336
rect 9815 26333 9827 26367
rect 9769 26327 9827 26333
rect 9953 26367 10011 26373
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 12161 26367 12219 26373
rect 12161 26333 12173 26367
rect 12207 26364 12219 26367
rect 12526 26364 12532 26376
rect 12207 26336 12532 26364
rect 12207 26333 12219 26336
rect 12161 26327 12219 26333
rect 12526 26324 12532 26336
rect 12584 26364 12590 26376
rect 12894 26364 12900 26376
rect 12584 26336 12900 26364
rect 12584 26324 12590 26336
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 13081 26367 13139 26373
rect 13081 26333 13093 26367
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26364 13507 26367
rect 13906 26364 13912 26376
rect 13495 26336 13912 26364
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 7331 26268 8340 26296
rect 7331 26265 7343 26268
rect 7285 26259 7343 26265
rect 8938 26256 8944 26308
rect 8996 26305 9002 26308
rect 8996 26299 9017 26305
rect 9005 26265 9017 26299
rect 9122 26296 9128 26308
rect 9083 26268 9128 26296
rect 8996 26259 9017 26265
rect 8996 26256 9002 26259
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 12986 26256 12992 26308
rect 13044 26296 13050 26308
rect 13096 26296 13124 26327
rect 13906 26324 13912 26336
rect 13964 26324 13970 26376
rect 14458 26324 14464 26376
rect 14516 26364 14522 26376
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 14516 26336 14841 26364
rect 14516 26324 14522 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 17402 26364 17408 26376
rect 17363 26336 17408 26364
rect 14829 26327 14887 26333
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 17512 26373 17540 26404
rect 17497 26367 17555 26373
rect 17497 26333 17509 26367
rect 17543 26333 17555 26367
rect 17497 26327 17555 26333
rect 17589 26367 17647 26373
rect 17589 26333 17601 26367
rect 17635 26333 17647 26367
rect 17589 26327 17647 26333
rect 13044 26268 13124 26296
rect 13357 26299 13415 26305
rect 13044 26256 13050 26268
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 14476 26296 14504 26324
rect 13403 26268 14504 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 15746 26256 15752 26308
rect 15804 26296 15810 26308
rect 17604 26296 17632 26327
rect 15804 26268 17632 26296
rect 17696 26296 17724 26404
rect 17788 26373 17816 26472
rect 19242 26432 19248 26444
rect 19203 26404 19248 26432
rect 19242 26392 19248 26404
rect 19300 26392 19306 26444
rect 19426 26432 19432 26444
rect 19387 26404 19432 26432
rect 19426 26392 19432 26404
rect 19484 26392 19490 26444
rect 21545 26435 21603 26441
rect 21545 26401 21557 26435
rect 21591 26432 21603 26435
rect 22370 26432 22376 26444
rect 21591 26404 22376 26432
rect 21591 26401 21603 26404
rect 21545 26395 21603 26401
rect 22370 26392 22376 26404
rect 22428 26432 22434 26444
rect 25685 26435 25743 26441
rect 25685 26432 25697 26435
rect 22428 26404 25697 26432
rect 22428 26392 22434 26404
rect 25685 26401 25697 26404
rect 25731 26432 25743 26435
rect 27246 26432 27252 26444
rect 25731 26404 27252 26432
rect 25731 26401 25743 26404
rect 25685 26395 25743 26401
rect 27246 26392 27252 26404
rect 27304 26432 27310 26444
rect 29549 26435 29607 26441
rect 29549 26432 29561 26435
rect 27304 26404 29561 26432
rect 27304 26392 27310 26404
rect 29549 26401 29561 26404
rect 29595 26401 29607 26435
rect 29549 26395 29607 26401
rect 31018 26392 31024 26444
rect 31076 26432 31082 26444
rect 31297 26435 31355 26441
rect 31297 26432 31309 26435
rect 31076 26404 31309 26432
rect 31076 26392 31082 26404
rect 31297 26401 31309 26404
rect 31343 26401 31355 26435
rect 31297 26395 31355 26401
rect 17773 26367 17831 26373
rect 17773 26333 17785 26367
rect 17819 26333 17831 26367
rect 17773 26327 17831 26333
rect 17862 26324 17868 26376
rect 17920 26364 17926 26376
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 17920 26336 18245 26364
rect 17920 26324 17926 26336
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 25406 26364 25412 26376
rect 24903 26336 25412 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 25406 26324 25412 26336
rect 25464 26324 25470 26376
rect 18138 26296 18144 26308
rect 17696 26268 18144 26296
rect 15804 26256 15810 26268
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 21085 26299 21143 26305
rect 21085 26265 21097 26299
rect 21131 26296 21143 26299
rect 21174 26296 21180 26308
rect 21131 26268 21180 26296
rect 21131 26265 21143 26268
rect 21085 26259 21143 26265
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 21818 26296 21824 26308
rect 21779 26268 21824 26296
rect 21818 26256 21824 26268
rect 21876 26256 21882 26308
rect 22094 26256 22100 26308
rect 22152 26296 22158 26308
rect 22152 26268 22310 26296
rect 22152 26256 22158 26268
rect 24946 26256 24952 26308
rect 25004 26296 25010 26308
rect 25041 26299 25099 26305
rect 25041 26296 25053 26299
rect 25004 26268 25053 26296
rect 25004 26256 25010 26268
rect 25041 26265 25053 26268
rect 25087 26265 25099 26299
rect 25958 26296 25964 26308
rect 25919 26268 25964 26296
rect 25041 26259 25099 26265
rect 25958 26256 25964 26268
rect 26016 26256 26022 26308
rect 26418 26256 26424 26308
rect 26476 26256 26482 26308
rect 29822 26296 29828 26308
rect 29783 26268 29828 26296
rect 29822 26256 29828 26268
rect 29880 26256 29886 26308
rect 30374 26256 30380 26308
rect 30432 26256 30438 26308
rect 31404 26296 31432 26540
rect 31754 26528 31760 26580
rect 31812 26568 31818 26580
rect 33594 26568 33600 26580
rect 31812 26540 33600 26568
rect 31812 26528 31818 26540
rect 33594 26528 33600 26540
rect 33652 26528 33658 26580
rect 33778 26568 33784 26580
rect 33739 26540 33784 26568
rect 33778 26528 33784 26540
rect 33836 26528 33842 26580
rect 47854 26568 47860 26580
rect 33888 26540 47860 26568
rect 31938 26460 31944 26512
rect 31996 26500 32002 26512
rect 33888 26500 33916 26540
rect 47854 26528 47860 26540
rect 47912 26528 47918 26580
rect 31996 26472 33916 26500
rect 35069 26503 35127 26509
rect 31996 26460 32002 26472
rect 35069 26469 35081 26503
rect 35115 26500 35127 26503
rect 36170 26500 36176 26512
rect 35115 26472 36176 26500
rect 35115 26469 35127 26472
rect 35069 26463 35127 26469
rect 36170 26460 36176 26472
rect 36228 26460 36234 26512
rect 32401 26435 32459 26441
rect 32401 26401 32413 26435
rect 32447 26432 32459 26435
rect 32582 26432 32588 26444
rect 32447 26404 32588 26432
rect 32447 26401 32459 26404
rect 32401 26395 32459 26401
rect 32582 26392 32588 26404
rect 32640 26392 32646 26444
rect 33042 26392 33048 26444
rect 33100 26432 33106 26444
rect 37553 26435 37611 26441
rect 37553 26432 37565 26435
rect 33100 26404 37565 26432
rect 33100 26392 33106 26404
rect 37553 26401 37565 26404
rect 37599 26401 37611 26435
rect 37553 26395 37611 26401
rect 37826 26392 37832 26444
rect 37884 26432 37890 26444
rect 40218 26432 40224 26444
rect 37884 26404 40224 26432
rect 37884 26392 37890 26404
rect 40218 26392 40224 26404
rect 40276 26432 40282 26444
rect 41141 26435 41199 26441
rect 41141 26432 41153 26435
rect 40276 26404 41153 26432
rect 40276 26392 40282 26404
rect 41141 26401 41153 26404
rect 41187 26401 41199 26435
rect 41141 26395 41199 26401
rect 31938 26324 31944 26376
rect 31996 26364 32002 26376
rect 32677 26367 32735 26373
rect 32677 26364 32689 26367
rect 31996 26336 32689 26364
rect 31996 26324 32002 26336
rect 32677 26333 32689 26336
rect 32723 26333 32735 26367
rect 33686 26364 33692 26376
rect 33647 26336 33692 26364
rect 32677 26327 32735 26333
rect 33686 26324 33692 26336
rect 33744 26324 33750 26376
rect 34882 26364 34888 26376
rect 34843 26336 34888 26364
rect 34882 26324 34888 26336
rect 34940 26324 34946 26376
rect 40865 26367 40923 26373
rect 40865 26333 40877 26367
rect 40911 26364 40923 26367
rect 41414 26364 41420 26376
rect 40911 26336 41420 26364
rect 40911 26333 40923 26336
rect 40865 26327 40923 26333
rect 41414 26324 41420 26336
rect 41472 26324 41478 26376
rect 45186 26324 45192 26376
rect 45244 26364 45250 26376
rect 47673 26367 47731 26373
rect 47673 26364 47685 26367
rect 45244 26336 47685 26364
rect 45244 26324 45250 26336
rect 47673 26333 47685 26336
rect 47719 26333 47731 26367
rect 47673 26327 47731 26333
rect 31754 26296 31760 26308
rect 31404 26268 31760 26296
rect 31754 26256 31760 26268
rect 31812 26256 31818 26308
rect 37826 26296 37832 26308
rect 37787 26268 37832 26296
rect 37826 26256 37832 26268
rect 37884 26256 37890 26308
rect 38378 26256 38384 26308
rect 38436 26256 38442 26308
rect 43990 26256 43996 26308
rect 44048 26296 44054 26308
rect 46842 26296 46848 26308
rect 44048 26268 46848 26296
rect 44048 26256 44054 26268
rect 46842 26256 46848 26268
rect 46900 26256 46906 26308
rect 7834 26228 7840 26240
rect 7795 26200 7840 26228
rect 7834 26188 7840 26200
rect 7892 26188 7898 26240
rect 8205 26231 8263 26237
rect 8205 26197 8217 26231
rect 8251 26228 8263 26231
rect 8294 26228 8300 26240
rect 8251 26200 8300 26228
rect 8251 26197 8263 26200
rect 8205 26191 8263 26197
rect 8294 26188 8300 26200
rect 8352 26228 8358 26240
rect 9214 26228 9220 26240
rect 8352 26200 9220 26228
rect 8352 26188 8358 26200
rect 9214 26188 9220 26200
rect 9272 26188 9278 26240
rect 9766 26188 9772 26240
rect 9824 26228 9830 26240
rect 10137 26231 10195 26237
rect 10137 26228 10149 26231
rect 9824 26200 10149 26228
rect 9824 26188 9830 26200
rect 10137 26197 10149 26200
rect 10183 26197 10195 26231
rect 10137 26191 10195 26197
rect 11333 26231 11391 26237
rect 11333 26197 11345 26231
rect 11379 26228 11391 26231
rect 11698 26228 11704 26240
rect 11379 26200 11704 26228
rect 11379 26197 11391 26200
rect 11333 26191 11391 26197
rect 11698 26188 11704 26200
rect 11756 26188 11762 26240
rect 13262 26228 13268 26240
rect 13223 26200 13268 26228
rect 13262 26188 13268 26200
rect 13320 26188 13326 26240
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 27433 26231 27491 26237
rect 27433 26228 27445 26231
rect 26844 26200 27445 26228
rect 26844 26188 26850 26200
rect 27433 26197 27445 26200
rect 27479 26197 27491 26231
rect 27433 26191 27491 26197
rect 38746 26188 38752 26240
rect 38804 26228 38810 26240
rect 39301 26231 39359 26237
rect 39301 26228 39313 26231
rect 38804 26200 39313 26228
rect 38804 26188 38810 26200
rect 39301 26197 39313 26200
rect 39347 26197 39359 26231
rect 39301 26191 39359 26197
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 11517 26027 11575 26033
rect 11517 25993 11529 26027
rect 11563 26024 11575 26027
rect 11790 26024 11796 26036
rect 11563 25996 11796 26024
rect 11563 25993 11575 25996
rect 11517 25987 11575 25993
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 12894 25984 12900 26036
rect 12952 26024 12958 26036
rect 13081 26027 13139 26033
rect 13081 26024 13093 26027
rect 12952 25996 13093 26024
rect 12952 25984 12958 25996
rect 13081 25993 13093 25996
rect 13127 25993 13139 26027
rect 13081 25987 13139 25993
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 14001 26027 14059 26033
rect 14001 26024 14013 26027
rect 13320 25996 14013 26024
rect 13320 25984 13326 25996
rect 14001 25993 14013 25996
rect 14047 25993 14059 26027
rect 14001 25987 14059 25993
rect 14277 26027 14335 26033
rect 14277 25993 14289 26027
rect 14323 26024 14335 26027
rect 15746 26024 15752 26036
rect 14323 25996 15752 26024
rect 14323 25993 14335 25996
rect 14277 25987 14335 25993
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 17862 26024 17868 26036
rect 16960 25996 17868 26024
rect 7561 25959 7619 25965
rect 7561 25925 7573 25959
rect 7607 25956 7619 25959
rect 7834 25956 7840 25968
rect 7607 25928 7840 25956
rect 7607 25925 7619 25928
rect 7561 25919 7619 25925
rect 7834 25916 7840 25928
rect 7892 25916 7898 25968
rect 9030 25956 9036 25968
rect 8786 25928 9036 25956
rect 9030 25916 9036 25928
rect 9088 25916 9094 25968
rect 12710 25916 12716 25968
rect 12768 25956 12774 25968
rect 13725 25959 13783 25965
rect 13725 25956 13737 25959
rect 12768 25928 13737 25956
rect 12768 25916 12774 25928
rect 13725 25925 13737 25928
rect 13771 25925 13783 25959
rect 13725 25919 13783 25925
rect 15381 25959 15439 25965
rect 15381 25925 15393 25959
rect 15427 25956 15439 25959
rect 16850 25956 16856 25968
rect 15427 25928 16856 25956
rect 15427 25925 15439 25928
rect 15381 25919 15439 25925
rect 16850 25916 16856 25928
rect 16908 25916 16914 25968
rect 16960 25965 16988 25996
rect 17862 25984 17868 25996
rect 17920 25984 17926 26036
rect 21821 26027 21879 26033
rect 21821 26024 21833 26027
rect 20640 25996 21833 26024
rect 16945 25959 17003 25965
rect 16945 25925 16957 25959
rect 16991 25925 17003 25959
rect 19610 25956 19616 25968
rect 19571 25928 19616 25956
rect 16945 25919 17003 25925
rect 19610 25916 19616 25928
rect 19668 25916 19674 25968
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25888 6791 25891
rect 7098 25888 7104 25900
rect 6779 25860 7104 25888
rect 6779 25857 6791 25860
rect 6733 25851 6791 25857
rect 7098 25848 7104 25860
rect 7156 25848 7162 25900
rect 11698 25888 11704 25900
rect 11659 25860 11704 25888
rect 11698 25848 11704 25860
rect 11756 25848 11762 25900
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 12492 25860 12537 25888
rect 12492 25848 12498 25860
rect 12802 25848 12808 25900
rect 12860 25888 12866 25900
rect 12897 25891 12955 25897
rect 12897 25888 12909 25891
rect 12860 25860 12909 25888
rect 12860 25848 12866 25860
rect 12897 25857 12909 25860
rect 12943 25857 12955 25891
rect 12897 25851 12955 25857
rect 12986 25848 12992 25900
rect 13044 25888 13050 25900
rect 13909 25891 13967 25897
rect 13909 25888 13921 25891
rect 13044 25860 13921 25888
rect 13044 25848 13050 25860
rect 13909 25857 13921 25860
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 14093 25891 14151 25897
rect 14093 25857 14105 25891
rect 14139 25888 14151 25891
rect 14458 25888 14464 25900
rect 14139 25860 14464 25888
rect 14139 25857 14151 25860
rect 14093 25851 14151 25857
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25888 14795 25891
rect 15010 25888 15016 25900
rect 14783 25860 15016 25888
rect 14783 25857 14795 25860
rect 14737 25851 14795 25857
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25888 15715 25891
rect 15746 25888 15752 25900
rect 15703 25860 15752 25888
rect 15703 25857 15715 25860
rect 15657 25851 15715 25857
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 20640 25897 20668 25996
rect 21821 25993 21833 25996
rect 21867 25993 21879 26027
rect 21821 25987 21879 25993
rect 21910 25984 21916 26036
rect 21968 26024 21974 26036
rect 23934 26024 23940 26036
rect 21968 25996 23940 26024
rect 21968 25984 21974 25996
rect 23934 25984 23940 25996
rect 23992 25984 23998 26036
rect 26973 26027 27031 26033
rect 26973 25993 26985 26027
rect 27019 26024 27031 26027
rect 27154 26024 27160 26036
rect 27019 25996 27160 26024
rect 27019 25993 27031 25996
rect 26973 25987 27031 25993
rect 27154 25984 27160 25996
rect 27212 25984 27218 26036
rect 27982 25984 27988 26036
rect 28040 26024 28046 26036
rect 28537 26027 28595 26033
rect 28537 26024 28549 26027
rect 28040 25996 28549 26024
rect 28040 25984 28046 25996
rect 28537 25993 28549 25996
rect 28583 25993 28595 26027
rect 28537 25987 28595 25993
rect 29546 25984 29552 26036
rect 29604 25984 29610 26036
rect 29733 26027 29791 26033
rect 29733 25993 29745 26027
rect 29779 26024 29791 26027
rect 29822 26024 29828 26036
rect 29779 25996 29828 26024
rect 29779 25993 29791 25996
rect 29733 25987 29791 25993
rect 29822 25984 29828 25996
rect 29880 25984 29886 26036
rect 30190 26024 30196 26036
rect 29932 25996 30196 26024
rect 22189 25959 22247 25965
rect 22189 25925 22201 25959
rect 22235 25925 22247 25959
rect 22189 25919 22247 25925
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25857 15899 25891
rect 15841 25851 15899 25857
rect 20625 25891 20683 25897
rect 20625 25857 20637 25891
rect 20671 25857 20683 25891
rect 21082 25888 21088 25900
rect 21043 25860 21088 25888
rect 20625 25851 20683 25857
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25820 6883 25823
rect 7285 25823 7343 25829
rect 7285 25820 7297 25823
rect 6871 25792 7297 25820
rect 6871 25789 6883 25792
rect 6825 25783 6883 25789
rect 7285 25789 7297 25792
rect 7331 25789 7343 25823
rect 7285 25783 7343 25789
rect 11238 25780 11244 25832
rect 11296 25820 11302 25832
rect 15856 25820 15884 25851
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 21266 25888 21272 25900
rect 21227 25860 21272 25888
rect 21266 25848 21272 25860
rect 21324 25848 21330 25900
rect 22204 25888 22232 25919
rect 22278 25916 22284 25968
rect 22336 25956 22342 25968
rect 22336 25928 22381 25956
rect 22336 25916 22342 25928
rect 23566 25916 23572 25968
rect 23624 25956 23630 25968
rect 25317 25959 25375 25965
rect 23624 25928 24992 25956
rect 23624 25916 23630 25928
rect 22554 25888 22560 25900
rect 22204 25860 22560 25888
rect 22554 25848 22560 25860
rect 22612 25888 22618 25900
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22612 25860 22845 25888
rect 22612 25848 22618 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23385 25891 23443 25897
rect 23385 25857 23397 25891
rect 23431 25888 23443 25891
rect 24026 25888 24032 25900
rect 23431 25860 24032 25888
rect 23431 25857 23443 25860
rect 23385 25851 23443 25857
rect 24026 25848 24032 25860
rect 24084 25848 24090 25900
rect 24670 25888 24676 25900
rect 24631 25860 24676 25888
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 24854 25888 24860 25900
rect 24815 25860 24860 25888
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 24964 25897 24992 25928
rect 25317 25925 25329 25959
rect 25363 25956 25375 25959
rect 27798 25956 27804 25968
rect 25363 25928 27804 25956
rect 25363 25925 25375 25928
rect 25317 25919 25375 25925
rect 27798 25916 27804 25928
rect 27856 25916 27862 25968
rect 28169 25959 28227 25965
rect 28169 25925 28181 25959
rect 28215 25956 28227 25959
rect 28718 25956 28724 25968
rect 28215 25928 28724 25956
rect 28215 25925 28227 25928
rect 28169 25919 28227 25925
rect 28718 25916 28724 25928
rect 28776 25916 28782 25968
rect 29365 25959 29423 25965
rect 29365 25925 29377 25959
rect 29411 25956 29423 25959
rect 29564 25956 29592 25984
rect 29932 25956 29960 25996
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 30285 26027 30343 26033
rect 30285 25993 30297 26027
rect 30331 26024 30343 26027
rect 30374 26024 30380 26036
rect 30331 25996 30380 26024
rect 30331 25993 30343 25996
rect 30285 25987 30343 25993
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 31573 26027 31631 26033
rect 31573 25993 31585 26027
rect 31619 26024 31631 26027
rect 36170 26024 36176 26036
rect 31619 25996 32168 26024
rect 31619 25993 31631 25996
rect 31573 25987 31631 25993
rect 29411 25928 29960 25956
rect 30208 25928 32076 25956
rect 29411 25925 29423 25928
rect 29365 25919 29423 25925
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25857 25007 25891
rect 24949 25851 25007 25857
rect 25042 25891 25100 25897
rect 25042 25857 25054 25891
rect 25088 25888 25100 25891
rect 25130 25888 25136 25900
rect 25088 25860 25136 25888
rect 25088 25857 25100 25860
rect 25042 25851 25100 25857
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 25774 25888 25780 25900
rect 25735 25860 25780 25888
rect 25774 25848 25780 25860
rect 25832 25848 25838 25900
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 27338 25888 27344 25900
rect 27299 25860 27344 25888
rect 25961 25851 26019 25857
rect 11296 25792 15884 25820
rect 16117 25823 16175 25829
rect 11296 25780 11302 25792
rect 16117 25789 16129 25823
rect 16163 25820 16175 25823
rect 17126 25820 17132 25832
rect 16163 25792 17132 25820
rect 16163 25789 16175 25792
rect 16117 25783 16175 25789
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17770 25820 17776 25832
rect 17731 25792 17776 25820
rect 17770 25780 17776 25792
rect 17828 25780 17834 25832
rect 17954 25820 17960 25832
rect 17915 25792 17960 25820
rect 17954 25780 17960 25792
rect 18012 25780 18018 25832
rect 22465 25823 22523 25829
rect 22465 25789 22477 25823
rect 22511 25820 22523 25823
rect 23661 25823 23719 25829
rect 23661 25820 23673 25823
rect 22511 25792 23673 25820
rect 22511 25789 22523 25792
rect 22465 25783 22523 25789
rect 23661 25789 23673 25792
rect 23707 25820 23719 25823
rect 24118 25820 24124 25832
rect 23707 25792 24124 25820
rect 23707 25789 23719 25792
rect 23661 25783 23719 25789
rect 24118 25780 24124 25792
rect 24176 25820 24182 25832
rect 25976 25820 26004 25851
rect 27338 25848 27344 25860
rect 27396 25848 27402 25900
rect 28353 25891 28411 25897
rect 28353 25857 28365 25891
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 24176 25792 26004 25820
rect 24176 25780 24182 25792
rect 16025 25755 16083 25761
rect 16025 25721 16037 25755
rect 16071 25752 16083 25755
rect 18138 25752 18144 25764
rect 16071 25724 18144 25752
rect 16071 25721 16083 25724
rect 16025 25715 16083 25721
rect 18138 25712 18144 25724
rect 18196 25712 18202 25764
rect 21085 25755 21143 25761
rect 21085 25721 21097 25755
rect 21131 25752 21143 25755
rect 25976 25752 26004 25792
rect 27154 25780 27160 25832
rect 27212 25820 27218 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 27212 25792 27445 25820
rect 27212 25780 27218 25792
rect 27433 25789 27445 25792
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 27617 25823 27675 25829
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 28368 25820 28396 25851
rect 28994 25848 29000 25900
rect 29052 25888 29058 25900
rect 29089 25891 29147 25897
rect 29089 25888 29101 25891
rect 29052 25860 29101 25888
rect 29052 25848 29058 25860
rect 29089 25857 29101 25860
rect 29135 25857 29147 25891
rect 29089 25851 29147 25857
rect 29237 25891 29295 25897
rect 29237 25857 29249 25891
rect 29283 25888 29295 25891
rect 29283 25860 29408 25888
rect 29283 25857 29295 25860
rect 29237 25851 29295 25857
rect 27663 25792 28396 25820
rect 29380 25820 29408 25860
rect 29454 25848 29460 25900
rect 29512 25888 29518 25900
rect 29638 25897 29644 25900
rect 29595 25891 29644 25897
rect 29512 25860 29557 25888
rect 29512 25848 29518 25860
rect 29595 25857 29607 25891
rect 29641 25857 29644 25891
rect 29595 25851 29644 25857
rect 29638 25848 29644 25851
rect 29696 25848 29702 25900
rect 30208 25897 30236 25928
rect 30193 25891 30251 25897
rect 30193 25857 30205 25891
rect 30239 25857 30251 25891
rect 30193 25851 30251 25857
rect 31205 25891 31263 25897
rect 31205 25857 31217 25891
rect 31251 25888 31263 25891
rect 31938 25888 31944 25900
rect 31251 25860 31944 25888
rect 31251 25857 31263 25860
rect 31205 25851 31263 25857
rect 31938 25848 31944 25860
rect 31996 25848 32002 25900
rect 31018 25820 31024 25832
rect 29380 25792 31024 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 27632 25752 27660 25783
rect 31018 25780 31024 25792
rect 31076 25780 31082 25832
rect 31294 25820 31300 25832
rect 31255 25792 31300 25820
rect 31294 25780 31300 25792
rect 31352 25780 31358 25832
rect 21131 25724 21956 25752
rect 25976 25724 27660 25752
rect 32048 25752 32076 25928
rect 32140 25820 32168 25996
rect 33336 25996 36176 26024
rect 32493 25959 32551 25965
rect 32493 25925 32505 25959
rect 32539 25956 32551 25959
rect 32582 25956 32588 25968
rect 32539 25928 32588 25956
rect 32539 25925 32551 25928
rect 32493 25919 32551 25925
rect 32582 25916 32588 25928
rect 32640 25916 32646 25968
rect 32585 25823 32643 25829
rect 32585 25820 32597 25823
rect 32140 25792 32597 25820
rect 32585 25789 32597 25792
rect 32631 25789 32643 25823
rect 32585 25783 32643 25789
rect 32769 25823 32827 25829
rect 32769 25789 32781 25823
rect 32815 25820 32827 25823
rect 33336 25820 33364 25996
rect 36170 25984 36176 25996
rect 36228 25984 36234 26036
rect 37461 26027 37519 26033
rect 37461 25993 37473 26027
rect 37507 26024 37519 26027
rect 37826 26024 37832 26036
rect 37507 25996 37832 26024
rect 37507 25993 37519 25996
rect 37461 25987 37519 25993
rect 37826 25984 37832 25996
rect 37884 25984 37890 26036
rect 33502 25956 33508 25968
rect 33463 25928 33508 25956
rect 33502 25916 33508 25928
rect 33560 25916 33566 25968
rect 34790 25916 34796 25968
rect 34848 25956 34854 25968
rect 40402 25956 40408 25968
rect 34848 25928 35006 25956
rect 37844 25928 40408 25956
rect 34848 25916 34854 25928
rect 33686 25888 33692 25900
rect 32815 25792 33364 25820
rect 33428 25860 33692 25888
rect 32815 25789 32827 25792
rect 32769 25783 32827 25789
rect 33428 25752 33456 25860
rect 33686 25848 33692 25860
rect 33744 25848 33750 25900
rect 37734 25888 37740 25900
rect 37695 25860 37740 25888
rect 37734 25848 37740 25860
rect 37792 25848 37798 25900
rect 37844 25897 37872 25928
rect 40402 25916 40408 25928
rect 40460 25916 40466 25968
rect 41046 25956 41052 25968
rect 41007 25928 41052 25956
rect 41046 25916 41052 25928
rect 41104 25916 41110 25968
rect 41138 25916 41144 25968
rect 41196 25956 41202 25968
rect 45646 25956 45652 25968
rect 41196 25928 45652 25956
rect 41196 25916 41202 25928
rect 45646 25916 45652 25928
rect 45704 25916 45710 25968
rect 37829 25891 37887 25897
rect 37829 25857 37841 25891
rect 37875 25857 37887 25891
rect 37829 25851 37887 25857
rect 37918 25848 37924 25900
rect 37976 25888 37982 25900
rect 38105 25891 38163 25897
rect 37976 25860 38021 25888
rect 37976 25848 37982 25860
rect 38105 25857 38117 25891
rect 38151 25857 38163 25891
rect 38105 25851 38163 25857
rect 34241 25823 34299 25829
rect 34241 25820 34253 25823
rect 32048 25724 33456 25752
rect 33612 25792 34253 25820
rect 21131 25721 21143 25724
rect 21085 25715 21143 25721
rect 9033 25687 9091 25693
rect 9033 25653 9045 25687
rect 9079 25684 9091 25687
rect 9214 25684 9220 25696
rect 9079 25656 9220 25684
rect 9079 25653 9091 25656
rect 9033 25647 9091 25653
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 12066 25644 12072 25696
rect 12124 25684 12130 25696
rect 12253 25687 12311 25693
rect 12253 25684 12265 25687
rect 12124 25656 12265 25684
rect 12124 25644 12130 25656
rect 12253 25653 12265 25656
rect 12299 25653 12311 25687
rect 14826 25684 14832 25696
rect 14787 25656 14832 25684
rect 12253 25647 12311 25653
rect 14826 25644 14832 25656
rect 14884 25644 14890 25696
rect 17034 25684 17040 25696
rect 16995 25656 17040 25684
rect 17034 25644 17040 25656
rect 17092 25644 17098 25696
rect 20441 25687 20499 25693
rect 20441 25653 20453 25687
rect 20487 25684 20499 25687
rect 21818 25684 21824 25696
rect 20487 25656 21824 25684
rect 20487 25653 20499 25656
rect 20441 25647 20499 25653
rect 21818 25644 21824 25656
rect 21876 25644 21882 25696
rect 21928 25684 21956 25724
rect 22186 25684 22192 25696
rect 21928 25656 22192 25684
rect 22186 25644 22192 25656
rect 22244 25644 22250 25696
rect 25958 25644 25964 25696
rect 26016 25684 26022 25696
rect 26145 25687 26203 25693
rect 26145 25684 26157 25687
rect 26016 25656 26157 25684
rect 26016 25644 26022 25656
rect 26145 25653 26157 25656
rect 26191 25653 26203 25687
rect 26145 25647 26203 25653
rect 27338 25644 27344 25696
rect 27396 25684 27402 25696
rect 28074 25684 28080 25696
rect 27396 25656 28080 25684
rect 27396 25644 27402 25656
rect 28074 25644 28080 25656
rect 28132 25644 28138 25696
rect 32125 25687 32183 25693
rect 32125 25653 32137 25687
rect 32171 25684 32183 25687
rect 32398 25684 32404 25696
rect 32171 25656 32404 25684
rect 32171 25653 32183 25656
rect 32125 25647 32183 25653
rect 32398 25644 32404 25656
rect 32456 25644 32462 25696
rect 33042 25644 33048 25696
rect 33100 25684 33106 25696
rect 33612 25693 33640 25792
rect 34241 25789 34253 25792
rect 34287 25789 34299 25823
rect 34514 25820 34520 25832
rect 34475 25792 34520 25820
rect 34241 25783 34299 25789
rect 34514 25780 34520 25792
rect 34572 25780 34578 25832
rect 38120 25752 38148 25851
rect 38194 25848 38200 25900
rect 38252 25888 38258 25900
rect 38565 25891 38623 25897
rect 38565 25888 38577 25891
rect 38252 25860 38577 25888
rect 38252 25848 38258 25860
rect 38565 25857 38577 25860
rect 38611 25857 38623 25891
rect 38746 25888 38752 25900
rect 38707 25860 38752 25888
rect 38565 25851 38623 25857
rect 38746 25848 38752 25860
rect 38804 25848 38810 25900
rect 40218 25888 40224 25900
rect 40179 25860 40224 25888
rect 40218 25848 40224 25860
rect 40276 25848 40282 25900
rect 45554 25848 45560 25900
rect 45612 25888 45618 25900
rect 46477 25891 46535 25897
rect 46477 25888 46489 25891
rect 45612 25860 46489 25888
rect 45612 25848 45618 25860
rect 46477 25857 46489 25860
rect 46523 25857 46535 25891
rect 46477 25851 46535 25857
rect 38933 25755 38991 25761
rect 38933 25752 38945 25755
rect 38120 25724 38945 25752
rect 38933 25721 38945 25724
rect 38979 25721 38991 25755
rect 38933 25715 38991 25721
rect 33597 25687 33655 25693
rect 33597 25684 33609 25687
rect 33100 25656 33609 25684
rect 33100 25644 33106 25656
rect 33597 25653 33609 25656
rect 33643 25653 33655 25687
rect 33597 25647 33655 25653
rect 33686 25644 33692 25696
rect 33744 25684 33750 25696
rect 35526 25684 35532 25696
rect 33744 25656 35532 25684
rect 33744 25644 33750 25656
rect 35526 25644 35532 25656
rect 35584 25684 35590 25696
rect 35989 25687 36047 25693
rect 35989 25684 36001 25687
rect 35584 25656 36001 25684
rect 35584 25644 35590 25656
rect 35989 25653 36001 25656
rect 36035 25653 36047 25687
rect 35989 25647 36047 25653
rect 38286 25644 38292 25696
rect 38344 25684 38350 25696
rect 38565 25687 38623 25693
rect 38565 25684 38577 25687
rect 38344 25656 38577 25684
rect 38344 25644 38350 25656
rect 38565 25653 38577 25656
rect 38611 25653 38623 25687
rect 38565 25647 38623 25653
rect 46474 25644 46480 25696
rect 46532 25684 46538 25696
rect 46569 25687 46627 25693
rect 46569 25684 46581 25687
rect 46532 25656 46581 25684
rect 46532 25644 46538 25656
rect 46569 25653 46581 25656
rect 46615 25653 46627 25687
rect 47762 25684 47768 25696
rect 47723 25656 47768 25684
rect 46569 25647 46627 25653
rect 47762 25644 47768 25656
rect 47820 25644 47826 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 9030 25480 9036 25492
rect 8991 25452 9036 25480
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 13262 25440 13268 25492
rect 13320 25480 13326 25492
rect 13541 25483 13599 25489
rect 13541 25480 13553 25483
rect 13320 25452 13553 25480
rect 13320 25440 13326 25452
rect 13541 25449 13553 25452
rect 13587 25449 13599 25483
rect 13541 25443 13599 25449
rect 20993 25483 21051 25489
rect 20993 25449 21005 25483
rect 21039 25480 21051 25483
rect 22094 25480 22100 25492
rect 21039 25452 22100 25480
rect 21039 25449 21051 25452
rect 20993 25443 21051 25449
rect 12066 25344 12072 25356
rect 12027 25316 12072 25344
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7561 25279 7619 25285
rect 7561 25276 7573 25279
rect 7156 25248 7573 25276
rect 7156 25236 7162 25248
rect 7561 25245 7573 25248
rect 7607 25245 7619 25279
rect 7561 25239 7619 25245
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25276 8999 25279
rect 9030 25276 9036 25288
rect 8987 25248 9036 25276
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 9030 25236 9036 25248
rect 9088 25236 9094 25288
rect 9766 25276 9772 25288
rect 9727 25248 9772 25276
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 11790 25276 11796 25288
rect 11751 25248 11796 25276
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 13556 25276 13584 25443
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 22189 25483 22247 25489
rect 22189 25449 22201 25483
rect 22235 25480 22247 25483
rect 23474 25480 23480 25492
rect 22235 25452 23480 25480
rect 22235 25449 22247 25452
rect 22189 25443 22247 25449
rect 23474 25440 23480 25452
rect 23532 25440 23538 25492
rect 23934 25440 23940 25492
rect 23992 25480 23998 25492
rect 25501 25483 25559 25489
rect 23992 25452 24992 25480
rect 23992 25440 23998 25452
rect 19889 25415 19947 25421
rect 19889 25381 19901 25415
rect 19935 25412 19947 25415
rect 20070 25412 20076 25424
rect 19935 25384 20076 25412
rect 19935 25381 19947 25384
rect 19889 25375 19947 25381
rect 20070 25372 20076 25384
rect 20128 25412 20134 25424
rect 22738 25412 22744 25424
rect 20128 25384 22744 25412
rect 20128 25372 20134 25384
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 22925 25415 22983 25421
rect 22925 25381 22937 25415
rect 22971 25412 22983 25415
rect 23106 25412 23112 25424
rect 22971 25384 23112 25412
rect 22971 25381 22983 25384
rect 22925 25375 22983 25381
rect 23106 25372 23112 25384
rect 23164 25372 23170 25424
rect 23492 25412 23520 25440
rect 24765 25415 24823 25421
rect 24765 25412 24777 25415
rect 23492 25384 24777 25412
rect 24765 25381 24777 25384
rect 24811 25381 24823 25415
rect 24765 25375 24823 25381
rect 24854 25372 24860 25424
rect 24912 25372 24918 25424
rect 13906 25304 13912 25356
rect 13964 25344 13970 25356
rect 13964 25316 14596 25344
rect 13964 25304 13970 25316
rect 13814 25276 13820 25288
rect 13556 25248 13820 25276
rect 13814 25236 13820 25248
rect 13872 25276 13878 25288
rect 14568 25285 14596 25316
rect 14826 25304 14832 25356
rect 14884 25344 14890 25356
rect 15841 25347 15899 25353
rect 15841 25344 15853 25347
rect 14884 25316 15853 25344
rect 14884 25304 14890 25316
rect 15841 25313 15853 25316
rect 15887 25313 15899 25347
rect 17494 25344 17500 25356
rect 17455 25316 17500 25344
rect 15841 25307 15899 25313
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 21726 25344 21732 25356
rect 18524 25316 21732 25344
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 13872 25248 14289 25276
rect 13872 25236 13878 25248
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 14277 25239 14335 25245
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 15657 25279 15715 25285
rect 15657 25245 15669 25279
rect 15703 25245 15715 25279
rect 15657 25239 15715 25245
rect 1673 25211 1731 25217
rect 1673 25177 1685 25211
rect 1719 25208 1731 25211
rect 1762 25208 1768 25220
rect 1719 25180 1768 25208
rect 1719 25177 1731 25180
rect 1673 25171 1731 25177
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 13078 25168 13084 25220
rect 13136 25168 13142 25220
rect 14292 25208 14320 25239
rect 15672 25208 15700 25239
rect 17126 25236 17132 25288
rect 17184 25276 17190 25288
rect 18524 25285 18552 25316
rect 21726 25304 21732 25316
rect 21784 25304 21790 25356
rect 24872 25344 24900 25372
rect 24780 25316 24900 25344
rect 18509 25279 18567 25285
rect 18509 25276 18521 25279
rect 17184 25248 18521 25276
rect 17184 25236 17190 25248
rect 18509 25245 18521 25248
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 20990 25276 20996 25288
rect 20947 25248 20996 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 20990 25236 20996 25248
rect 21048 25236 21054 25288
rect 22830 25276 22836 25288
rect 22112 25248 22836 25276
rect 14292 25180 15700 25208
rect 18138 25168 18144 25220
rect 18196 25208 18202 25220
rect 18325 25211 18383 25217
rect 18325 25208 18337 25211
rect 18196 25180 18337 25208
rect 18196 25168 18202 25180
rect 18325 25177 18337 25180
rect 18371 25177 18383 25211
rect 18325 25171 18383 25177
rect 18693 25211 18751 25217
rect 18693 25177 18705 25211
rect 18739 25208 18751 25211
rect 19334 25208 19340 25220
rect 18739 25180 19340 25208
rect 18739 25177 18751 25180
rect 18693 25171 18751 25177
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19702 25208 19708 25220
rect 19484 25180 19708 25208
rect 19484 25168 19490 25180
rect 19702 25168 19708 25180
rect 19760 25168 19766 25220
rect 21266 25168 21272 25220
rect 21324 25208 21330 25220
rect 21821 25211 21879 25217
rect 21821 25208 21833 25211
rect 21324 25180 21833 25208
rect 21324 25168 21330 25180
rect 21821 25177 21833 25180
rect 21867 25177 21879 25211
rect 22002 25208 22008 25220
rect 21963 25180 22008 25208
rect 21821 25171 21879 25177
rect 7558 25100 7564 25152
rect 7616 25140 7622 25152
rect 7745 25143 7803 25149
rect 7745 25140 7757 25143
rect 7616 25112 7757 25140
rect 7616 25100 7622 25112
rect 7745 25109 7757 25112
rect 7791 25109 7803 25143
rect 9582 25140 9588 25152
rect 9543 25112 9588 25140
rect 7745 25103 7803 25109
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 14090 25140 14096 25152
rect 14051 25112 14096 25140
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14458 25140 14464 25152
rect 14371 25112 14464 25140
rect 14458 25100 14464 25112
rect 14516 25140 14522 25152
rect 15102 25140 15108 25152
rect 14516 25112 15108 25140
rect 14516 25100 14522 25112
rect 15102 25100 15108 25112
rect 15160 25100 15166 25152
rect 21836 25140 21864 25171
rect 22002 25168 22008 25180
rect 22060 25168 22066 25220
rect 22112 25140 22140 25248
rect 22830 25236 22836 25248
rect 22888 25236 22894 25288
rect 23017 25279 23075 25285
rect 23017 25254 23029 25279
rect 22940 25245 23029 25254
rect 23063 25245 23075 25279
rect 22940 25239 23075 25245
rect 23109 25279 23167 25285
rect 23109 25245 23121 25279
rect 23155 25254 23167 25279
rect 23155 25245 23244 25254
rect 23109 25239 23244 25245
rect 22940 25226 23060 25239
rect 23124 25226 23244 25239
rect 23290 25236 23296 25288
rect 23348 25276 23354 25288
rect 24611 25279 24669 25285
rect 24611 25276 24623 25279
rect 23348 25248 23393 25276
rect 23348 25236 23354 25248
rect 24596 25245 24623 25276
rect 24657 25270 24669 25279
rect 24780 25270 24808 25316
rect 24657 25245 24808 25270
rect 24596 25242 24808 25245
rect 24857 25279 24915 25285
rect 24857 25245 24869 25279
rect 24903 25276 24915 25279
rect 24964 25276 24992 25452
rect 25501 25449 25513 25483
rect 25547 25480 25559 25483
rect 26234 25480 26240 25492
rect 25547 25452 26240 25480
rect 25547 25449 25559 25452
rect 25501 25443 25559 25449
rect 26234 25440 26240 25452
rect 26292 25480 26298 25492
rect 26878 25480 26884 25492
rect 26292 25452 26884 25480
rect 26292 25440 26298 25452
rect 26878 25440 26884 25452
rect 26936 25440 26942 25492
rect 27154 25480 27160 25492
rect 27115 25452 27160 25480
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 28074 25440 28080 25492
rect 28132 25480 28138 25492
rect 28132 25452 33364 25480
rect 28132 25440 28138 25452
rect 29730 25372 29736 25424
rect 29788 25412 29794 25424
rect 30193 25415 30251 25421
rect 30193 25412 30205 25415
rect 29788 25384 30205 25412
rect 29788 25372 29794 25384
rect 30193 25381 30205 25384
rect 30239 25381 30251 25415
rect 30193 25375 30251 25381
rect 31941 25415 31999 25421
rect 31941 25381 31953 25415
rect 31987 25412 31999 25415
rect 32306 25412 32312 25424
rect 31987 25384 32312 25412
rect 31987 25381 31999 25384
rect 31941 25375 31999 25381
rect 32306 25372 32312 25384
rect 32364 25372 32370 25424
rect 33134 25372 33140 25424
rect 33192 25412 33198 25424
rect 33229 25415 33287 25421
rect 33229 25412 33241 25415
rect 33192 25384 33241 25412
rect 33192 25372 33198 25384
rect 33229 25381 33241 25384
rect 33275 25381 33287 25415
rect 33336 25412 33364 25452
rect 34514 25440 34520 25492
rect 34572 25480 34578 25492
rect 35345 25483 35403 25489
rect 35345 25480 35357 25483
rect 34572 25452 35357 25480
rect 34572 25440 34578 25452
rect 35345 25449 35357 25452
rect 35391 25449 35403 25483
rect 35345 25443 35403 25449
rect 37001 25483 37059 25489
rect 37001 25449 37013 25483
rect 37047 25480 37059 25483
rect 37918 25480 37924 25492
rect 37047 25452 37924 25480
rect 37047 25449 37059 25452
rect 37001 25443 37059 25449
rect 37918 25440 37924 25452
rect 37976 25440 37982 25492
rect 41138 25412 41144 25424
rect 33336 25384 41144 25412
rect 33229 25375 33287 25381
rect 41138 25372 41144 25384
rect 41196 25372 41202 25424
rect 26234 25304 26240 25356
rect 26292 25344 26298 25356
rect 26697 25347 26755 25353
rect 26697 25344 26709 25347
rect 26292 25316 26709 25344
rect 26292 25304 26298 25316
rect 26697 25313 26709 25316
rect 26743 25313 26755 25347
rect 32398 25344 32404 25356
rect 32359 25316 32404 25344
rect 26697 25307 26755 25313
rect 32398 25304 32404 25316
rect 32456 25304 32462 25356
rect 32490 25304 32496 25356
rect 32548 25344 32554 25356
rect 33413 25347 33471 25353
rect 32548 25316 32593 25344
rect 32548 25304 32554 25316
rect 33413 25313 33425 25347
rect 33459 25344 33471 25347
rect 33686 25344 33692 25356
rect 33459 25316 33692 25344
rect 33459 25313 33471 25316
rect 33413 25307 33471 25313
rect 33686 25304 33692 25316
rect 33744 25304 33750 25356
rect 33965 25347 34023 25353
rect 33965 25313 33977 25347
rect 34011 25344 34023 25347
rect 35526 25344 35532 25356
rect 34011 25316 34836 25344
rect 34011 25313 34023 25316
rect 33965 25307 34023 25313
rect 26786 25276 26792 25288
rect 24903 25248 24992 25276
rect 26747 25248 26792 25276
rect 24903 25245 24915 25248
rect 24611 25239 24669 25242
rect 24857 25239 24915 25245
rect 26786 25236 26792 25248
rect 26844 25236 26850 25288
rect 30009 25279 30067 25285
rect 30009 25245 30021 25279
rect 30055 25276 30067 25279
rect 30098 25276 30104 25288
rect 30055 25248 30104 25276
rect 30055 25245 30067 25248
rect 30009 25239 30067 25245
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 31938 25236 31944 25288
rect 31996 25276 32002 25288
rect 32309 25279 32367 25285
rect 32309 25276 32321 25279
rect 31996 25248 32321 25276
rect 31996 25236 32002 25248
rect 32309 25245 32321 25248
rect 32355 25276 32367 25279
rect 32950 25276 32956 25288
rect 32355 25248 32956 25276
rect 32355 25245 32367 25248
rect 32309 25239 32367 25245
rect 32950 25236 32956 25248
rect 33008 25276 33014 25288
rect 33137 25279 33195 25285
rect 33137 25276 33149 25279
rect 33008 25248 33149 25276
rect 33008 25236 33014 25248
rect 33137 25245 33149 25248
rect 33183 25245 33195 25279
rect 33137 25239 33195 25245
rect 33873 25279 33931 25285
rect 33873 25245 33885 25279
rect 33919 25245 33931 25279
rect 34054 25276 34060 25288
rect 34015 25248 34060 25276
rect 33873 25239 33931 25245
rect 22738 25168 22744 25220
rect 22796 25208 22802 25220
rect 22940 25208 22968 25226
rect 22796 25180 22968 25208
rect 23216 25208 23244 25226
rect 24302 25208 24308 25220
rect 23216 25180 24308 25208
rect 22796 25168 22802 25180
rect 24302 25168 24308 25180
rect 24360 25168 24366 25220
rect 24397 25211 24455 25217
rect 24397 25177 24409 25211
rect 24443 25208 24455 25211
rect 25409 25211 25467 25217
rect 25409 25208 25421 25211
rect 24443 25180 25421 25208
rect 24443 25177 24455 25180
rect 24397 25171 24455 25177
rect 25409 25177 25421 25180
rect 25455 25208 25467 25211
rect 28626 25208 28632 25220
rect 25455 25180 28632 25208
rect 25455 25177 25467 25180
rect 25409 25171 25467 25177
rect 28626 25168 28632 25180
rect 28684 25168 28690 25220
rect 33413 25211 33471 25217
rect 33413 25177 33425 25211
rect 33459 25208 33471 25211
rect 33888 25208 33916 25239
rect 34054 25236 34060 25248
rect 34112 25236 34118 25288
rect 34808 25285 34836 25316
rect 35084 25316 35532 25344
rect 35084 25285 35112 25316
rect 35526 25304 35532 25316
rect 35584 25304 35590 25356
rect 37458 25344 37464 25356
rect 36740 25316 37464 25344
rect 34701 25279 34759 25285
rect 34701 25245 34713 25279
rect 34747 25245 34759 25279
rect 34701 25239 34759 25245
rect 34794 25279 34852 25285
rect 34794 25245 34806 25279
rect 34840 25245 34852 25279
rect 34794 25239 34852 25245
rect 35069 25279 35127 25285
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 35207 25279 35265 25285
rect 35207 25245 35219 25279
rect 35253 25276 35265 25279
rect 35434 25276 35440 25288
rect 35253 25248 35440 25276
rect 35253 25245 35265 25248
rect 35207 25239 35265 25245
rect 33459 25180 33916 25208
rect 34716 25208 34744 25239
rect 35434 25236 35440 25248
rect 35492 25236 35498 25288
rect 36740 25285 36768 25316
rect 37458 25304 37464 25316
rect 37516 25304 37522 25356
rect 38286 25304 38292 25356
rect 38344 25344 38350 25356
rect 38381 25347 38439 25353
rect 38381 25344 38393 25347
rect 38344 25316 38393 25344
rect 38344 25304 38350 25316
rect 38381 25313 38393 25316
rect 38427 25313 38439 25347
rect 38381 25307 38439 25313
rect 40310 25304 40316 25356
rect 40368 25344 40374 25356
rect 40770 25344 40776 25356
rect 40368 25316 40776 25344
rect 40368 25304 40374 25316
rect 40770 25304 40776 25316
rect 40828 25344 40834 25356
rect 45738 25344 45744 25356
rect 40828 25316 45744 25344
rect 40828 25304 40834 25316
rect 45738 25304 45744 25316
rect 45796 25304 45802 25356
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 48130 25344 48136 25356
rect 48091 25316 48136 25344
rect 48130 25304 48136 25316
rect 48188 25304 48194 25356
rect 36725 25279 36783 25285
rect 36725 25245 36737 25279
rect 36771 25245 36783 25279
rect 36725 25239 36783 25245
rect 37001 25279 37059 25285
rect 37001 25245 37013 25279
rect 37047 25276 37059 25279
rect 37090 25276 37096 25288
rect 37047 25248 37096 25276
rect 37047 25245 37059 25248
rect 37001 25239 37059 25245
rect 37090 25236 37096 25248
rect 37148 25236 37154 25288
rect 38010 25236 38016 25288
rect 38068 25276 38074 25288
rect 38105 25279 38163 25285
rect 38105 25276 38117 25279
rect 38068 25248 38117 25276
rect 38068 25236 38074 25248
rect 38105 25245 38117 25248
rect 38151 25245 38163 25279
rect 40218 25276 40224 25288
rect 40179 25248 40224 25276
rect 38105 25239 38163 25245
rect 40218 25236 40224 25248
rect 40276 25236 40282 25288
rect 46290 25276 46296 25288
rect 46251 25248 46296 25276
rect 46290 25236 46296 25248
rect 46348 25236 46354 25288
rect 34977 25211 35035 25217
rect 34716 25180 34836 25208
rect 33459 25177 33471 25180
rect 33413 25171 33471 25177
rect 21836 25112 22140 25140
rect 22649 25143 22707 25149
rect 22649 25109 22661 25143
rect 22695 25140 22707 25143
rect 23474 25140 23480 25152
rect 22695 25112 23480 25140
rect 22695 25109 22707 25112
rect 22649 25103 22707 25109
rect 23474 25100 23480 25112
rect 23532 25100 23538 25152
rect 34808 25140 34836 25180
rect 34977 25177 34989 25211
rect 35023 25208 35035 25211
rect 35802 25208 35808 25220
rect 35023 25180 35808 25208
rect 35023 25177 35035 25180
rect 34977 25171 35035 25177
rect 35802 25168 35808 25180
rect 35860 25168 35866 25220
rect 36078 25168 36084 25220
rect 36136 25208 36142 25220
rect 36909 25211 36967 25217
rect 36909 25208 36921 25211
rect 36136 25180 36921 25208
rect 36136 25168 36142 25180
rect 36909 25177 36921 25180
rect 36955 25177 36967 25211
rect 36909 25171 36967 25177
rect 38654 25140 38660 25152
rect 34808 25112 38660 25140
rect 38654 25100 38660 25112
rect 38712 25100 38718 25152
rect 45646 25100 45652 25152
rect 45704 25140 45710 25152
rect 46106 25140 46112 25152
rect 45704 25112 46112 25140
rect 45704 25100 45710 25112
rect 46106 25100 46112 25112
rect 46164 25100 46170 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 12434 24896 12440 24948
rect 12492 24936 12498 24948
rect 13081 24939 13139 24945
rect 13081 24936 13093 24939
rect 12492 24908 13093 24936
rect 12492 24896 12498 24908
rect 13081 24905 13093 24908
rect 13127 24905 13139 24939
rect 13081 24899 13139 24905
rect 17221 24939 17279 24945
rect 17221 24905 17233 24939
rect 17267 24936 17279 24939
rect 17402 24936 17408 24948
rect 17267 24908 17408 24936
rect 17267 24905 17279 24908
rect 17221 24899 17279 24905
rect 14458 24868 14464 24880
rect 13740 24840 14464 24868
rect 7558 24800 7564 24812
rect 7519 24772 7564 24800
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 8938 24760 8944 24812
rect 8996 24760 9002 24812
rect 10318 24800 10324 24812
rect 10279 24772 10324 24800
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24800 11575 24803
rect 12897 24803 12955 24809
rect 11563 24772 12434 24800
rect 11563 24769 11575 24772
rect 11517 24763 11575 24769
rect 7837 24735 7895 24741
rect 7837 24701 7849 24735
rect 7883 24732 7895 24735
rect 9582 24732 9588 24744
rect 7883 24704 9588 24732
rect 7883 24701 7895 24704
rect 7837 24695 7895 24701
rect 9582 24692 9588 24704
rect 9640 24692 9646 24744
rect 9030 24624 9036 24676
rect 9088 24664 9094 24676
rect 11532 24664 11560 24763
rect 9088 24636 11560 24664
rect 12406 24664 12434 24772
rect 12897 24769 12909 24803
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 13541 24803 13599 24809
rect 13541 24769 13553 24803
rect 13587 24800 13599 24803
rect 13630 24800 13636 24812
rect 13587 24772 13636 24800
rect 13587 24769 13599 24772
rect 13541 24763 13599 24769
rect 12710 24732 12716 24744
rect 12671 24704 12716 24732
rect 12710 24692 12716 24704
rect 12768 24732 12774 24744
rect 12912 24732 12940 24763
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13740 24809 13768 24840
rect 14458 24828 14464 24840
rect 14516 24828 14522 24880
rect 17236 24868 17264 24899
rect 17402 24896 17408 24908
rect 17460 24936 17466 24948
rect 19426 24936 19432 24948
rect 17460 24908 19432 24936
rect 17460 24896 17466 24908
rect 19426 24896 19432 24908
rect 19484 24896 19490 24948
rect 23290 24936 23296 24948
rect 22572 24908 23296 24936
rect 16960 24840 17264 24868
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 15746 24800 15752 24812
rect 13872 24772 13917 24800
rect 15707 24772 15752 24800
rect 13872 24760 13878 24772
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16960 24800 16988 24840
rect 17126 24800 17132 24812
rect 16071 24772 16988 24800
rect 17087 24772 17132 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 17126 24760 17132 24772
rect 17184 24760 17190 24812
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24800 17831 24803
rect 17862 24800 17868 24812
rect 17819 24772 17868 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 20990 24800 20996 24812
rect 20951 24772 20996 24800
rect 20990 24760 20996 24772
rect 21048 24760 21054 24812
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22572 24809 22600 24908
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 24026 24896 24032 24948
rect 24084 24936 24090 24948
rect 24397 24939 24455 24945
rect 24397 24936 24409 24939
rect 24084 24908 24409 24936
rect 24084 24896 24090 24908
rect 24397 24905 24409 24908
rect 24443 24905 24455 24939
rect 24397 24899 24455 24905
rect 24854 24896 24860 24948
rect 24912 24936 24918 24948
rect 26053 24939 26111 24945
rect 26053 24936 26065 24939
rect 24912 24908 26065 24936
rect 24912 24896 24918 24908
rect 26053 24905 26065 24908
rect 26099 24905 26111 24939
rect 26053 24899 26111 24905
rect 29454 24896 29460 24948
rect 29512 24936 29518 24948
rect 30282 24936 30288 24948
rect 29512 24908 30288 24936
rect 29512 24896 29518 24908
rect 30282 24896 30288 24908
rect 30340 24896 30346 24948
rect 32490 24936 32496 24948
rect 31220 24908 32496 24936
rect 25130 24828 25136 24880
rect 25188 24868 25194 24880
rect 25188 24840 26464 24868
rect 25188 24828 25194 24840
rect 22557 24803 22615 24809
rect 22557 24800 22569 24803
rect 22060 24772 22569 24800
rect 22060 24760 22066 24772
rect 22557 24769 22569 24772
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 23474 24800 23480 24812
rect 22704 24772 22749 24800
rect 23435 24772 23480 24800
rect 22704 24760 22710 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 23661 24803 23719 24809
rect 23661 24769 23673 24803
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24800 23811 24803
rect 23934 24800 23940 24812
rect 23799 24772 23940 24800
rect 23799 24769 23811 24772
rect 23753 24763 23811 24769
rect 14090 24732 14096 24744
rect 12768 24704 12848 24732
rect 12912 24704 14096 24732
rect 12768 24692 12774 24704
rect 12526 24664 12532 24676
rect 12406 24636 12532 24664
rect 9088 24624 9094 24636
rect 12526 24624 12532 24636
rect 12584 24624 12590 24676
rect 12820 24664 12848 24704
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 22094 24732 22100 24744
rect 16132 24704 22100 24732
rect 13633 24667 13691 24673
rect 13633 24664 13645 24667
rect 12820 24636 13645 24664
rect 13633 24633 13645 24636
rect 13679 24633 13691 24667
rect 16132 24664 16160 24704
rect 22094 24692 22100 24704
rect 22152 24692 22158 24744
rect 22186 24692 22192 24744
rect 22244 24732 22250 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 22244 24704 22385 24732
rect 22244 24692 22250 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 22462 24692 22468 24744
rect 22520 24732 22526 24744
rect 23676 24732 23704 24763
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 22520 24704 22565 24732
rect 23676 24704 23796 24732
rect 22520 24692 22526 24704
rect 13633 24627 13691 24633
rect 13740 24636 16160 24664
rect 8846 24556 8852 24608
rect 8904 24596 8910 24608
rect 9309 24599 9367 24605
rect 9309 24596 9321 24599
rect 8904 24568 9321 24596
rect 8904 24556 8910 24568
rect 9309 24565 9321 24568
rect 9355 24565 9367 24599
rect 9309 24559 9367 24565
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10413 24599 10471 24605
rect 10413 24596 10425 24599
rect 10008 24568 10425 24596
rect 10008 24556 10014 24568
rect 10413 24565 10425 24568
rect 10459 24565 10471 24599
rect 11606 24596 11612 24608
rect 11567 24568 11612 24596
rect 10413 24559 10471 24565
rect 11606 24556 11612 24568
rect 11664 24556 11670 24608
rect 12894 24556 12900 24608
rect 12952 24596 12958 24608
rect 13740 24596 13768 24636
rect 20346 24624 20352 24676
rect 20404 24664 20410 24676
rect 23293 24667 23351 24673
rect 23293 24664 23305 24667
rect 20404 24636 23305 24664
rect 20404 24624 20410 24636
rect 23293 24633 23305 24636
rect 23339 24633 23351 24667
rect 23293 24627 23351 24633
rect 12952 24568 13768 24596
rect 12952 24556 12958 24568
rect 13814 24556 13820 24608
rect 13872 24596 13878 24608
rect 15565 24599 15623 24605
rect 15565 24596 15577 24599
rect 13872 24568 15577 24596
rect 13872 24556 13878 24568
rect 15565 24565 15577 24568
rect 15611 24565 15623 24599
rect 15565 24559 15623 24565
rect 15933 24599 15991 24605
rect 15933 24565 15945 24599
rect 15979 24596 15991 24599
rect 16850 24596 16856 24608
rect 15979 24568 16856 24596
rect 15979 24565 15991 24568
rect 15933 24559 15991 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17494 24556 17500 24608
rect 17552 24596 17558 24608
rect 17957 24599 18015 24605
rect 17957 24596 17969 24599
rect 17552 24568 17969 24596
rect 17552 24556 17558 24568
rect 17957 24565 17969 24568
rect 18003 24565 18015 24599
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 17957 24559 18015 24565
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 22189 24599 22247 24605
rect 22189 24565 22201 24599
rect 22235 24596 22247 24599
rect 22278 24596 22284 24608
rect 22235 24568 22284 24596
rect 22235 24565 22247 24568
rect 22189 24559 22247 24565
rect 22278 24556 22284 24568
rect 22336 24556 22342 24608
rect 23768 24596 23796 24704
rect 24320 24664 24348 24763
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 25961 24803 26019 24809
rect 25961 24800 25973 24803
rect 25924 24772 25973 24800
rect 25924 24760 25930 24772
rect 25961 24769 25973 24772
rect 26007 24769 26019 24803
rect 25961 24763 26019 24769
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26326 24800 26332 24812
rect 26191 24772 26332 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 26326 24760 26332 24772
rect 26384 24760 26390 24812
rect 26436 24809 26464 24840
rect 29472 24840 30696 24868
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24769 26479 24803
rect 26421 24763 26479 24769
rect 27065 24803 27123 24809
rect 27065 24769 27077 24803
rect 27111 24800 27123 24803
rect 27614 24800 27620 24812
rect 27111 24772 27620 24800
rect 27111 24769 27123 24772
rect 27065 24763 27123 24769
rect 27614 24760 27620 24772
rect 27672 24760 27678 24812
rect 28626 24800 28632 24812
rect 28587 24772 28632 24800
rect 28626 24760 28632 24772
rect 28684 24800 28690 24812
rect 29365 24803 29423 24809
rect 29365 24800 29377 24803
rect 28684 24772 29377 24800
rect 28684 24760 28690 24772
rect 29365 24769 29377 24772
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 25685 24735 25743 24741
rect 25685 24701 25697 24735
rect 25731 24732 25743 24735
rect 26234 24732 26240 24744
rect 25731 24704 26240 24732
rect 25731 24701 25743 24704
rect 25685 24695 25743 24701
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 27246 24732 27252 24744
rect 27207 24704 27252 24732
rect 27246 24692 27252 24704
rect 27304 24732 27310 24744
rect 27522 24732 27528 24744
rect 27304 24704 27528 24732
rect 27304 24692 27310 24704
rect 27522 24692 27528 24704
rect 27580 24692 27586 24744
rect 24670 24664 24676 24676
rect 24320 24636 24676 24664
rect 24670 24624 24676 24636
rect 24728 24664 24734 24676
rect 29472 24664 29500 24840
rect 29549 24803 29607 24809
rect 29549 24769 29561 24803
rect 29595 24800 29607 24803
rect 30098 24800 30104 24812
rect 29595 24772 30104 24800
rect 29595 24769 29607 24772
rect 29549 24763 29607 24769
rect 30098 24760 30104 24772
rect 30156 24760 30162 24812
rect 30377 24803 30435 24809
rect 30377 24769 30389 24803
rect 30423 24769 30435 24803
rect 30377 24763 30435 24769
rect 29825 24735 29883 24741
rect 29825 24701 29837 24735
rect 29871 24732 29883 24735
rect 30190 24732 30196 24744
rect 29871 24704 30196 24732
rect 29871 24701 29883 24704
rect 29825 24695 29883 24701
rect 30190 24692 30196 24704
rect 30248 24692 30254 24744
rect 30392 24732 30420 24763
rect 30466 24760 30472 24812
rect 30524 24800 30530 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 30524 24772 30573 24800
rect 30524 24760 30530 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30668 24800 30696 24840
rect 31220 24800 31248 24908
rect 32490 24896 32496 24908
rect 32548 24896 32554 24948
rect 33502 24936 33508 24948
rect 33415 24908 33508 24936
rect 33502 24896 33508 24908
rect 33560 24936 33566 24948
rect 34054 24936 34060 24948
rect 33560 24908 34060 24936
rect 33560 24896 33566 24908
rect 34054 24896 34060 24908
rect 34112 24896 34118 24948
rect 31294 24828 31300 24880
rect 31352 24868 31358 24880
rect 38010 24868 38016 24880
rect 31352 24840 33180 24868
rect 31352 24828 31358 24840
rect 32140 24809 32168 24840
rect 33152 24812 33180 24840
rect 37108 24840 38016 24868
rect 30668 24772 31248 24800
rect 32125 24803 32183 24809
rect 30561 24763 30619 24769
rect 32125 24769 32137 24803
rect 32171 24769 32183 24803
rect 32125 24763 32183 24769
rect 32401 24803 32459 24809
rect 32401 24769 32413 24803
rect 32447 24800 32459 24803
rect 32858 24800 32864 24812
rect 32447 24772 32864 24800
rect 32447 24769 32459 24772
rect 32401 24763 32459 24769
rect 32858 24760 32864 24772
rect 32916 24760 32922 24812
rect 33134 24800 33140 24812
rect 33095 24772 33140 24800
rect 33134 24760 33140 24772
rect 33192 24760 33198 24812
rect 33321 24803 33379 24809
rect 33321 24769 33333 24803
rect 33367 24800 33379 24803
rect 33686 24800 33692 24812
rect 33367 24772 33692 24800
rect 33367 24769 33379 24772
rect 33321 24763 33379 24769
rect 31754 24732 31760 24744
rect 30392 24704 31760 24732
rect 31754 24692 31760 24704
rect 31812 24692 31818 24744
rect 31938 24692 31944 24744
rect 31996 24732 32002 24744
rect 32217 24735 32275 24741
rect 32217 24732 32229 24735
rect 31996 24704 32229 24732
rect 31996 24692 32002 24704
rect 32217 24701 32229 24704
rect 32263 24701 32275 24735
rect 32217 24695 32275 24701
rect 32306 24692 32312 24744
rect 32364 24732 32370 24744
rect 33336 24732 33364 24763
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 34698 24760 34704 24812
rect 34756 24800 34762 24812
rect 37108 24800 37136 24840
rect 38010 24828 38016 24840
rect 38068 24828 38074 24880
rect 37274 24800 37280 24812
rect 34756 24772 37136 24800
rect 37235 24772 37280 24800
rect 34756 24760 34762 24772
rect 37274 24760 37280 24772
rect 37332 24760 37338 24812
rect 46014 24760 46020 24812
rect 46072 24800 46078 24812
rect 46477 24803 46535 24809
rect 46477 24800 46489 24803
rect 46072 24772 46489 24800
rect 46072 24760 46078 24772
rect 46477 24769 46489 24772
rect 46523 24769 46535 24803
rect 46477 24763 46535 24769
rect 47118 24760 47124 24812
rect 47176 24800 47182 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47176 24772 47593 24800
rect 47176 24760 47182 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 32364 24704 33364 24732
rect 32364 24692 32370 24704
rect 36998 24692 37004 24744
rect 37056 24732 37062 24744
rect 37553 24735 37611 24741
rect 37553 24732 37565 24735
rect 37056 24704 37565 24732
rect 37056 24692 37062 24704
rect 37553 24701 37565 24704
rect 37599 24732 37611 24735
rect 38746 24732 38752 24744
rect 37599 24704 38752 24732
rect 37599 24701 37611 24704
rect 37553 24695 37611 24701
rect 38746 24692 38752 24704
rect 38804 24692 38810 24744
rect 46198 24732 46204 24744
rect 46159 24704 46204 24732
rect 46198 24692 46204 24704
rect 46256 24692 46262 24744
rect 24728 24636 29500 24664
rect 24728 24624 24734 24636
rect 29914 24624 29920 24676
rect 29972 24664 29978 24676
rect 46750 24664 46756 24676
rect 29972 24636 46756 24664
rect 29972 24624 29978 24636
rect 46750 24624 46756 24636
rect 46808 24624 46814 24676
rect 24946 24596 24952 24608
rect 23768 24568 24952 24596
rect 24946 24556 24952 24568
rect 25004 24596 25010 24608
rect 26142 24596 26148 24608
rect 25004 24568 26148 24596
rect 25004 24556 25010 24568
rect 26142 24556 26148 24568
rect 26200 24556 26206 24608
rect 26326 24596 26332 24608
rect 26287 24568 26332 24596
rect 26326 24556 26332 24568
rect 26384 24556 26390 24608
rect 26510 24556 26516 24608
rect 26568 24596 26574 24608
rect 27982 24596 27988 24608
rect 26568 24568 27988 24596
rect 26568 24556 26574 24568
rect 27982 24556 27988 24568
rect 28040 24556 28046 24608
rect 28810 24596 28816 24608
rect 28771 24568 28816 24596
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 30006 24556 30012 24608
rect 30064 24596 30070 24608
rect 30469 24599 30527 24605
rect 30469 24596 30481 24599
rect 30064 24568 30481 24596
rect 30064 24556 30070 24568
rect 30469 24565 30481 24568
rect 30515 24565 30527 24599
rect 30469 24559 30527 24565
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 32306 24596 32312 24608
rect 31352 24568 32312 24596
rect 31352 24556 31358 24568
rect 32306 24556 32312 24568
rect 32364 24556 32370 24608
rect 32398 24556 32404 24608
rect 32456 24596 32462 24608
rect 32585 24599 32643 24605
rect 32585 24596 32597 24599
rect 32456 24568 32597 24596
rect 32456 24556 32462 24568
rect 32585 24565 32597 24568
rect 32631 24565 32643 24599
rect 32585 24559 32643 24565
rect 32950 24556 32956 24608
rect 33008 24596 33014 24608
rect 33137 24599 33195 24605
rect 33137 24596 33149 24599
rect 33008 24568 33149 24596
rect 33008 24556 33014 24568
rect 33137 24565 33149 24568
rect 33183 24565 33195 24599
rect 33137 24559 33195 24565
rect 36722 24556 36728 24608
rect 36780 24596 36786 24608
rect 37369 24599 37427 24605
rect 37369 24596 37381 24599
rect 36780 24568 37381 24596
rect 36780 24556 36786 24568
rect 37369 24565 37381 24568
rect 37415 24565 37427 24599
rect 37369 24559 37427 24565
rect 37458 24556 37464 24608
rect 37516 24596 37522 24608
rect 37516 24568 37561 24596
rect 37516 24556 37522 24568
rect 46474 24556 46480 24608
rect 46532 24596 46538 24608
rect 47673 24599 47731 24605
rect 47673 24596 47685 24599
rect 46532 24568 47685 24596
rect 46532 24556 46538 24568
rect 47673 24565 47685 24568
rect 47719 24565 47731 24599
rect 47673 24559 47731 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 12894 24392 12900 24404
rect 2746 24364 12900 24392
rect 1670 24284 1676 24336
rect 1728 24324 1734 24336
rect 2746 24324 2774 24364
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 13078 24392 13084 24404
rect 13035 24364 13084 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 21821 24395 21879 24401
rect 17236 24364 21404 24392
rect 1728 24296 2774 24324
rect 1728 24284 1734 24296
rect 8938 24284 8944 24336
rect 8996 24324 9002 24336
rect 9033 24327 9091 24333
rect 9033 24324 9045 24327
rect 8996 24296 9045 24324
rect 8996 24284 9002 24296
rect 9033 24293 9045 24296
rect 9079 24293 9091 24327
rect 9033 24287 9091 24293
rect 11790 24284 11796 24336
rect 11848 24324 11854 24336
rect 12345 24327 12403 24333
rect 12345 24324 12357 24327
rect 11848 24296 12357 24324
rect 11848 24284 11854 24296
rect 12345 24293 12357 24296
rect 12391 24293 12403 24327
rect 12345 24287 12403 24293
rect 1946 24216 1952 24268
rect 2004 24256 2010 24268
rect 17236 24256 17264 24364
rect 17497 24327 17555 24333
rect 17497 24293 17509 24327
rect 17543 24324 17555 24327
rect 17954 24324 17960 24336
rect 17543 24296 17960 24324
rect 17543 24293 17555 24296
rect 17497 24287 17555 24293
rect 17954 24284 17960 24296
rect 18012 24284 18018 24336
rect 21376 24324 21404 24364
rect 21821 24361 21833 24395
rect 21867 24392 21879 24395
rect 22002 24392 22008 24404
rect 21867 24364 22008 24392
rect 21867 24361 21879 24364
rect 21821 24355 21879 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 26234 24392 26240 24404
rect 22152 24364 22876 24392
rect 26195 24364 26240 24392
rect 22152 24352 22158 24364
rect 22738 24324 22744 24336
rect 21376 24296 22744 24324
rect 22738 24284 22744 24296
rect 22796 24284 22802 24336
rect 18138 24256 18144 24268
rect 2004 24228 17264 24256
rect 17328 24228 18144 24256
rect 2004 24216 2010 24228
rect 8941 24191 8999 24197
rect 8941 24157 8953 24191
rect 8987 24188 8999 24191
rect 9030 24188 9036 24200
rect 8987 24160 9036 24188
rect 8987 24157 8999 24160
rect 8941 24151 8999 24157
rect 9030 24148 9036 24160
rect 9088 24148 9094 24200
rect 9950 24188 9956 24200
rect 9911 24160 9956 24188
rect 9950 24148 9956 24160
rect 10008 24148 10014 24200
rect 12250 24188 12256 24200
rect 12211 24160 12256 24188
rect 12250 24148 12256 24160
rect 12308 24148 12314 24200
rect 12526 24148 12532 24200
rect 12584 24188 12590 24200
rect 12897 24191 12955 24197
rect 12897 24188 12909 24191
rect 12584 24160 12909 24188
rect 12584 24148 12590 24160
rect 12897 24157 12909 24160
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24188 16727 24191
rect 17328 24188 17356 24228
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 20073 24259 20131 24265
rect 20073 24225 20085 24259
rect 20119 24256 20131 24259
rect 22002 24256 22008 24268
rect 20119 24228 22008 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 22848 24197 22876 24364
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 28810 24392 28816 24404
rect 28771 24364 28816 24392
rect 28810 24352 28816 24364
rect 28868 24352 28874 24404
rect 28920 24364 30604 24392
rect 26145 24327 26203 24333
rect 26145 24293 26157 24327
rect 26191 24324 26203 24327
rect 26881 24327 26939 24333
rect 26881 24324 26893 24327
rect 26191 24296 26893 24324
rect 26191 24293 26203 24296
rect 26145 24287 26203 24293
rect 26881 24293 26893 24296
rect 26927 24293 26939 24327
rect 26881 24287 26939 24293
rect 26970 24284 26976 24336
rect 27028 24324 27034 24336
rect 28920 24324 28948 24364
rect 27028 24296 28948 24324
rect 28997 24327 29055 24333
rect 27028 24284 27034 24296
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 29687 24327 29745 24333
rect 29687 24324 29699 24327
rect 29043 24296 29699 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 29687 24293 29699 24296
rect 29733 24293 29745 24327
rect 29687 24287 29745 24293
rect 29825 24327 29883 24333
rect 29825 24293 29837 24327
rect 29871 24324 29883 24327
rect 30469 24327 30527 24333
rect 30469 24324 30481 24327
rect 29871 24296 30481 24324
rect 29871 24293 29883 24296
rect 29825 24287 29883 24293
rect 30469 24293 30481 24296
rect 30515 24293 30527 24327
rect 30576 24324 30604 24364
rect 30650 24352 30656 24404
rect 30708 24392 30714 24404
rect 31297 24395 31355 24401
rect 31297 24392 31309 24395
rect 30708 24364 31309 24392
rect 30708 24352 30714 24364
rect 31297 24361 31309 24364
rect 31343 24361 31355 24395
rect 31297 24355 31355 24361
rect 31757 24395 31815 24401
rect 31757 24361 31769 24395
rect 31803 24392 31815 24395
rect 31938 24392 31944 24404
rect 31803 24364 31944 24392
rect 31803 24361 31815 24364
rect 31757 24355 31815 24361
rect 31938 24352 31944 24364
rect 31996 24352 32002 24404
rect 35434 24352 35440 24404
rect 35492 24392 35498 24404
rect 36909 24395 36967 24401
rect 36909 24392 36921 24395
rect 35492 24364 36921 24392
rect 35492 24352 35498 24364
rect 36909 24361 36921 24364
rect 36955 24392 36967 24395
rect 37274 24392 37280 24404
rect 36955 24364 37280 24392
rect 36955 24361 36967 24364
rect 36909 24355 36967 24361
rect 37274 24352 37280 24364
rect 37332 24352 37338 24404
rect 37829 24395 37887 24401
rect 37829 24361 37841 24395
rect 37875 24392 37887 24395
rect 38286 24392 38292 24404
rect 37875 24364 38292 24392
rect 37875 24361 37887 24364
rect 37829 24355 37887 24361
rect 38286 24352 38292 24364
rect 38344 24352 38350 24404
rect 30742 24324 30748 24336
rect 30576 24296 30748 24324
rect 30469 24287 30527 24293
rect 30742 24284 30748 24296
rect 30800 24284 30806 24336
rect 32858 24324 32864 24336
rect 32140 24296 32864 24324
rect 23109 24259 23167 24265
rect 23109 24225 23121 24259
rect 23155 24256 23167 24259
rect 24026 24256 24032 24268
rect 23155 24228 24032 24256
rect 23155 24225 23167 24228
rect 23109 24219 23167 24225
rect 24026 24216 24032 24228
rect 24084 24216 24090 24268
rect 25866 24216 25872 24268
rect 25924 24256 25930 24268
rect 31481 24259 31539 24265
rect 25924 24228 27108 24256
rect 25924 24216 25930 24228
rect 16715 24160 17356 24188
rect 17405 24191 17463 24197
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 17405 24157 17417 24191
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 22833 24191 22891 24197
rect 19659 24160 20116 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 10134 24080 10140 24132
rect 10192 24120 10198 24132
rect 10229 24123 10287 24129
rect 10229 24120 10241 24123
rect 10192 24092 10241 24120
rect 10192 24080 10198 24092
rect 10229 24089 10241 24092
rect 10275 24089 10287 24123
rect 11606 24120 11612 24132
rect 11454 24092 11612 24120
rect 10229 24083 10287 24089
rect 11606 24080 11612 24092
rect 11664 24080 11670 24132
rect 17034 24080 17040 24132
rect 17092 24120 17098 24132
rect 17310 24120 17316 24132
rect 17092 24092 17316 24120
rect 17092 24080 17098 24092
rect 17310 24080 17316 24092
rect 17368 24120 17374 24132
rect 17420 24120 17448 24151
rect 17368 24092 17448 24120
rect 17368 24080 17374 24092
rect 9582 24012 9588 24064
rect 9640 24052 9646 24064
rect 11701 24055 11759 24061
rect 11701 24052 11713 24055
rect 9640 24024 11713 24052
rect 9640 24012 9646 24024
rect 11701 24021 11713 24024
rect 11747 24052 11759 24055
rect 12986 24052 12992 24064
rect 11747 24024 12992 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 16850 24052 16856 24064
rect 16763 24024 16856 24052
rect 16850 24012 16856 24024
rect 16908 24052 16914 24064
rect 17586 24052 17592 24064
rect 16908 24024 17592 24052
rect 16908 24012 16914 24024
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 19705 24055 19763 24061
rect 19705 24021 19717 24055
rect 19751 24052 19763 24055
rect 19978 24052 19984 24064
rect 19751 24024 19984 24052
rect 19751 24021 19763 24024
rect 19705 24015 19763 24021
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20088 24052 20116 24160
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 25958 24188 25964 24200
rect 25919 24160 25964 24188
rect 22833 24151 22891 24157
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26050 24148 26056 24200
rect 26108 24188 26114 24200
rect 26421 24191 26479 24197
rect 26108 24160 26153 24188
rect 26108 24148 26114 24160
rect 26421 24157 26433 24191
rect 26467 24157 26479 24191
rect 26878 24188 26884 24200
rect 26839 24160 26884 24188
rect 26421 24151 26479 24157
rect 20346 24120 20352 24132
rect 20307 24092 20352 24120
rect 20346 24080 20352 24092
rect 20404 24080 20410 24132
rect 21082 24080 21088 24132
rect 21140 24080 21146 24132
rect 21634 24080 21640 24132
rect 21692 24120 21698 24132
rect 26326 24120 26332 24132
rect 21692 24092 26332 24120
rect 21692 24080 21698 24092
rect 26326 24080 26332 24092
rect 26384 24080 26390 24132
rect 20990 24052 20996 24064
rect 20088 24024 20996 24052
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 22462 24052 22468 24064
rect 22423 24024 22468 24052
rect 22462 24012 22468 24024
rect 22520 24012 22526 24064
rect 22925 24055 22983 24061
rect 22925 24021 22937 24055
rect 22971 24052 22983 24055
rect 24394 24052 24400 24064
rect 22971 24024 24400 24052
rect 22971 24021 22983 24024
rect 22925 24015 22983 24021
rect 24394 24012 24400 24024
rect 24452 24012 24458 24064
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 25685 24055 25743 24061
rect 25685 24052 25697 24055
rect 25648 24024 25697 24052
rect 25648 24012 25654 24024
rect 25685 24021 25697 24024
rect 25731 24021 25743 24055
rect 25685 24015 25743 24021
rect 26142 24012 26148 24064
rect 26200 24052 26206 24064
rect 26436 24052 26464 24151
rect 26878 24148 26884 24160
rect 26936 24148 26942 24200
rect 27080 24197 27108 24228
rect 28644 24228 30880 24256
rect 27065 24191 27123 24197
rect 27065 24157 27077 24191
rect 27111 24157 27123 24191
rect 27065 24151 27123 24157
rect 28644 24129 28672 24228
rect 29454 24188 29460 24200
rect 28736 24160 29460 24188
rect 28629 24123 28687 24129
rect 28629 24089 28641 24123
rect 28675 24089 28687 24123
rect 28629 24083 28687 24089
rect 28736 24052 28764 24160
rect 29454 24148 29460 24160
rect 29512 24188 29518 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29512 24160 29561 24188
rect 29512 24148 29518 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 30006 24188 30012 24200
rect 29967 24160 30012 24188
rect 29549 24151 29607 24157
rect 30006 24148 30012 24160
rect 30064 24148 30070 24200
rect 30282 24188 30288 24200
rect 30116 24160 30288 24188
rect 28845 24123 28903 24129
rect 28845 24089 28857 24123
rect 28891 24120 28903 24123
rect 30116 24120 30144 24160
rect 30282 24148 30288 24160
rect 30340 24188 30346 24200
rect 30745 24191 30803 24197
rect 30745 24188 30757 24191
rect 30340 24160 30757 24188
rect 30340 24148 30346 24160
rect 30745 24157 30757 24160
rect 30791 24157 30803 24191
rect 30745 24151 30803 24157
rect 28891 24092 30144 24120
rect 30469 24123 30527 24129
rect 28891 24089 28903 24092
rect 28845 24083 28903 24089
rect 30469 24089 30481 24123
rect 30515 24120 30527 24123
rect 30852 24120 30880 24228
rect 31481 24225 31493 24259
rect 31527 24256 31539 24259
rect 32140 24256 32168 24296
rect 32858 24284 32864 24296
rect 32916 24324 32922 24336
rect 32916 24296 33180 24324
rect 32916 24284 32922 24296
rect 33045 24259 33103 24265
rect 33045 24256 33057 24259
rect 31527 24228 32168 24256
rect 32232 24228 33057 24256
rect 31527 24225 31539 24228
rect 31481 24219 31539 24225
rect 31294 24188 31300 24200
rect 31255 24160 31300 24188
rect 31294 24148 31300 24160
rect 31352 24148 31358 24200
rect 32232 24197 32260 24228
rect 33045 24225 33057 24228
rect 33091 24225 33103 24259
rect 33045 24219 33103 24225
rect 31573 24191 31631 24197
rect 31573 24182 31585 24191
rect 31496 24157 31585 24182
rect 31619 24157 31631 24191
rect 31496 24154 31631 24157
rect 31496 24120 31524 24154
rect 31573 24151 31631 24154
rect 32217 24191 32275 24197
rect 32217 24157 32229 24191
rect 32263 24157 32275 24191
rect 32398 24188 32404 24200
rect 32359 24160 32404 24188
rect 32217 24151 32275 24157
rect 32398 24148 32404 24160
rect 32456 24148 32462 24200
rect 32493 24191 32551 24197
rect 32493 24157 32505 24191
rect 32539 24188 32551 24191
rect 32766 24188 32772 24200
rect 32539 24160 32772 24188
rect 32539 24157 32551 24160
rect 32493 24151 32551 24157
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 33152 24197 33180 24296
rect 37090 24284 37096 24336
rect 37148 24324 37154 24336
rect 47762 24324 47768 24336
rect 37148 24296 37193 24324
rect 46308 24296 47768 24324
rect 37148 24284 37154 24296
rect 46308 24265 46336 24296
rect 47762 24284 47768 24296
rect 47820 24284 47826 24336
rect 36817 24259 36875 24265
rect 36817 24225 36829 24259
rect 36863 24225 36875 24259
rect 46293 24259 46351 24265
rect 36817 24219 36875 24225
rect 37568 24228 37872 24256
rect 32953 24191 33011 24197
rect 32953 24157 32965 24191
rect 32999 24157 33011 24191
rect 32953 24151 33011 24157
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24188 33195 24191
rect 33870 24188 33876 24200
rect 33183 24160 33876 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 30515 24092 30880 24120
rect 30515 24089 30527 24092
rect 30469 24083 30527 24089
rect 26200 24024 28764 24052
rect 26200 24012 26206 24024
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 29917 24055 29975 24061
rect 29917 24052 29929 24055
rect 29880 24024 29929 24052
rect 29880 24012 29886 24024
rect 29917 24021 29929 24024
rect 29963 24021 29975 24055
rect 29917 24015 29975 24021
rect 30653 24055 30711 24061
rect 30653 24021 30665 24055
rect 30699 24052 30711 24055
rect 30742 24052 30748 24064
rect 30699 24024 30748 24052
rect 30699 24021 30711 24024
rect 30653 24015 30711 24021
rect 30742 24012 30748 24024
rect 30800 24012 30806 24064
rect 30852 24052 30880 24092
rect 31312 24092 31524 24120
rect 31312 24064 31340 24092
rect 31662 24080 31668 24132
rect 31720 24120 31726 24132
rect 32416 24120 32444 24148
rect 31720 24092 32444 24120
rect 31720 24080 31726 24092
rect 31294 24052 31300 24064
rect 30852 24024 31300 24052
rect 31294 24012 31300 24024
rect 31352 24012 31358 24064
rect 32122 24012 32128 24064
rect 32180 24052 32186 24064
rect 32309 24055 32367 24061
rect 32309 24052 32321 24055
rect 32180 24024 32321 24052
rect 32180 24012 32186 24024
rect 32309 24021 32321 24024
rect 32355 24021 32367 24055
rect 32784 24052 32812 24148
rect 32968 24120 32996 24151
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 36173 24191 36231 24197
rect 36173 24157 36185 24191
rect 36219 24188 36231 24191
rect 36219 24160 36768 24188
rect 36219 24157 36231 24160
rect 36173 24151 36231 24157
rect 36740 24132 36768 24160
rect 33502 24120 33508 24132
rect 32968 24092 33508 24120
rect 33502 24080 33508 24092
rect 33560 24080 33566 24132
rect 35894 24120 35900 24132
rect 35855 24092 35900 24120
rect 35894 24080 35900 24092
rect 35952 24080 35958 24132
rect 36078 24120 36084 24132
rect 36004 24092 36084 24120
rect 36004 24052 36032 24092
rect 36078 24080 36084 24092
rect 36136 24120 36142 24132
rect 36136 24092 36229 24120
rect 36136 24080 36142 24092
rect 36354 24080 36360 24132
rect 36412 24120 36418 24132
rect 36633 24123 36691 24129
rect 36633 24120 36645 24123
rect 36412 24092 36645 24120
rect 36412 24080 36418 24092
rect 36633 24089 36645 24092
rect 36679 24089 36691 24123
rect 36633 24083 36691 24089
rect 36722 24080 36728 24132
rect 36780 24080 36786 24132
rect 36170 24052 36176 24064
rect 32784 24024 36032 24052
rect 36131 24024 36176 24052
rect 32309 24015 32367 24021
rect 36170 24012 36176 24024
rect 36228 24012 36234 24064
rect 36538 24012 36544 24064
rect 36596 24052 36602 24064
rect 36832 24052 36860 24219
rect 36998 24197 37004 24200
rect 36949 24191 37004 24197
rect 36949 24157 36961 24191
rect 36995 24157 37004 24191
rect 36949 24151 37004 24157
rect 36998 24148 37004 24151
rect 37056 24148 37062 24200
rect 37568 24052 37596 24228
rect 37844 24197 37872 24228
rect 46293 24225 46305 24259
rect 46339 24225 46351 24259
rect 46474 24256 46480 24268
rect 46435 24228 46480 24256
rect 46293 24219 46351 24225
rect 46474 24216 46480 24228
rect 46532 24216 46538 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 37650 24191 37708 24197
rect 37650 24157 37662 24191
rect 37696 24188 37708 24191
rect 37829 24191 37887 24197
rect 37696 24160 37780 24188
rect 37696 24157 37708 24160
rect 37650 24151 37708 24157
rect 37752 24132 37780 24160
rect 37829 24157 37841 24191
rect 37875 24188 37887 24191
rect 38562 24188 38568 24200
rect 37875 24160 38568 24188
rect 37875 24157 37887 24160
rect 37829 24151 37887 24157
rect 38562 24148 38568 24160
rect 38620 24148 38626 24200
rect 37734 24080 37740 24132
rect 37792 24120 37798 24132
rect 38194 24120 38200 24132
rect 37792 24092 38200 24120
rect 37792 24080 37798 24092
rect 38194 24080 38200 24092
rect 38252 24080 38258 24132
rect 36596 24024 37596 24052
rect 36596 24012 36602 24024
rect 37918 24012 37924 24064
rect 37976 24052 37982 24064
rect 38013 24055 38071 24061
rect 38013 24052 38025 24055
rect 37976 24024 38025 24052
rect 37976 24012 37982 24024
rect 38013 24021 38025 24024
rect 38059 24021 38071 24055
rect 38013 24015 38071 24021
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1946 23848 1952 23860
rect 1907 23820 1952 23848
rect 1946 23808 1952 23820
rect 2004 23808 2010 23860
rect 10134 23848 10140 23860
rect 10095 23820 10140 23848
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 15102 23848 15108 23860
rect 11572 23820 15108 23848
rect 11572 23808 11578 23820
rect 15102 23808 15108 23820
rect 15160 23808 15166 23860
rect 18432 23820 25544 23848
rect 12710 23780 12716 23792
rect 9876 23752 12716 23780
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 9582 23712 9588 23724
rect 8812 23684 9588 23712
rect 8812 23672 8818 23684
rect 9582 23672 9588 23684
rect 9640 23712 9646 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9640 23684 9781 23712
rect 9640 23672 9646 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9876 23653 9904 23752
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 14274 23740 14280 23792
rect 14332 23740 14338 23792
rect 15120 23780 15148 23808
rect 15120 23752 17724 23780
rect 11514 23712 11520 23724
rect 11475 23684 11520 23712
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 12250 23712 12256 23724
rect 11716 23684 12256 23712
rect 9861 23647 9919 23653
rect 9861 23613 9873 23647
rect 9907 23613 9919 23647
rect 9861 23607 9919 23613
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11716 23517 11744 23684
rect 12250 23672 12256 23684
rect 12308 23712 12314 23724
rect 12437 23715 12495 23721
rect 12437 23712 12449 23715
rect 12308 23684 12449 23712
rect 12308 23672 12314 23684
rect 12437 23681 12449 23684
rect 12483 23681 12495 23715
rect 12437 23675 12495 23681
rect 15010 23672 15016 23724
rect 15068 23712 15074 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 15068 23684 16681 23712
rect 15068 23672 15074 23684
rect 16669 23681 16681 23684
rect 16715 23712 16727 23715
rect 17494 23712 17500 23724
rect 16715 23684 17500 23712
rect 16715 23681 16727 23684
rect 16669 23675 16727 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 17696 23721 17724 23752
rect 18432 23721 18460 23820
rect 19978 23780 19984 23792
rect 19918 23752 19984 23780
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 22738 23740 22744 23792
rect 22796 23780 22802 23792
rect 22796 23752 24532 23780
rect 22796 23740 22802 23752
rect 17681 23715 17739 23721
rect 17681 23681 17693 23715
rect 17727 23681 17739 23715
rect 17681 23675 17739 23681
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23681 18475 23715
rect 22462 23712 22468 23724
rect 22423 23684 22468 23712
rect 18417 23675 18475 23681
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 12575 23616 13461 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 13449 23613 13461 23616
rect 13495 23613 13507 23647
rect 13449 23607 13507 23613
rect 13725 23647 13783 23653
rect 13725 23613 13737 23647
rect 13771 23644 13783 23647
rect 14458 23644 14464 23656
rect 13771 23616 14464 23644
rect 13771 23613 13783 23616
rect 13725 23607 13783 23613
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 17696 23576 17724 23675
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 24029 23715 24087 23721
rect 24029 23681 24041 23715
rect 24075 23681 24087 23715
rect 24029 23675 24087 23681
rect 18693 23647 18751 23653
rect 18693 23613 18705 23647
rect 18739 23644 18751 23647
rect 19242 23644 19248 23656
rect 18739 23616 19248 23644
rect 18739 23613 18751 23616
rect 18693 23607 18751 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 17696 23548 18184 23576
rect 11701 23511 11759 23517
rect 11701 23508 11713 23511
rect 11020 23480 11713 23508
rect 11020 23468 11026 23480
rect 11701 23477 11713 23480
rect 11747 23477 11759 23511
rect 11701 23471 11759 23477
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 13814 23508 13820 23520
rect 12400 23480 13820 23508
rect 12400 23468 12406 23480
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 14366 23508 14372 23520
rect 13872 23480 14372 23508
rect 13872 23468 13878 23480
rect 14366 23468 14372 23480
rect 14424 23468 14430 23520
rect 15194 23508 15200 23520
rect 15155 23480 15200 23508
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 16758 23508 16764 23520
rect 16719 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 17865 23511 17923 23517
rect 17865 23477 17877 23511
rect 17911 23508 17923 23511
rect 18046 23508 18052 23520
rect 17911 23480 18052 23508
rect 17911 23477 17923 23480
rect 17865 23471 17923 23477
rect 18046 23468 18052 23480
rect 18104 23468 18110 23520
rect 18156 23508 18184 23548
rect 20165 23511 20223 23517
rect 20165 23508 20177 23511
rect 18156 23480 20177 23508
rect 20165 23477 20177 23480
rect 20211 23477 20223 23511
rect 22278 23508 22284 23520
rect 22239 23480 22284 23508
rect 20165 23471 20223 23477
rect 22278 23468 22284 23480
rect 22336 23468 22342 23520
rect 23750 23468 23756 23520
rect 23808 23508 23814 23520
rect 24044 23508 24072 23675
rect 24121 23647 24179 23653
rect 24121 23613 24133 23647
rect 24167 23613 24179 23647
rect 24394 23644 24400 23656
rect 24355 23616 24400 23644
rect 24121 23607 24179 23613
rect 24136 23576 24164 23607
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 24504 23644 24532 23752
rect 25516 23712 25544 23820
rect 26050 23808 26056 23860
rect 26108 23848 26114 23860
rect 26329 23851 26387 23857
rect 26329 23848 26341 23851
rect 26108 23820 26341 23848
rect 26108 23808 26114 23820
rect 26329 23817 26341 23820
rect 26375 23817 26387 23851
rect 26329 23811 26387 23817
rect 26418 23808 26424 23860
rect 26476 23848 26482 23860
rect 26878 23848 26884 23860
rect 26476 23820 26884 23848
rect 26476 23808 26482 23820
rect 26878 23808 26884 23820
rect 26936 23808 26942 23860
rect 31110 23848 31116 23860
rect 27172 23820 31116 23848
rect 25866 23740 25872 23792
rect 25924 23780 25930 23792
rect 27065 23783 27123 23789
rect 27065 23780 27077 23783
rect 25924 23752 27077 23780
rect 25924 23740 25930 23752
rect 26142 23712 26148 23724
rect 25516 23684 26148 23712
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23712 26295 23715
rect 26326 23712 26332 23724
rect 26283 23684 26332 23712
rect 26283 23681 26295 23684
rect 26237 23675 26295 23681
rect 26326 23672 26332 23684
rect 26384 23672 26390 23724
rect 26436 23721 26464 23752
rect 27065 23749 27077 23752
rect 27111 23749 27123 23783
rect 27065 23743 27123 23749
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23681 26479 23715
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26421 23675 26479 23681
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27172 23644 27200 23820
rect 31110 23808 31116 23820
rect 31168 23808 31174 23860
rect 31294 23848 31300 23860
rect 31255 23820 31300 23848
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 31846 23808 31852 23860
rect 31904 23848 31910 23860
rect 31904 23820 32260 23848
rect 31904 23808 31910 23820
rect 29822 23780 29828 23792
rect 29783 23752 29828 23780
rect 29822 23740 29828 23752
rect 29880 23740 29886 23792
rect 31202 23780 31208 23792
rect 31050 23752 31208 23780
rect 31202 23740 31208 23752
rect 31260 23740 31266 23792
rect 27522 23672 27528 23724
rect 27580 23712 27586 23724
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 27580 23684 29561 23712
rect 27580 23672 27586 23684
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 31846 23712 31852 23724
rect 29549 23675 29607 23681
rect 31036 23684 31852 23712
rect 24504 23616 27200 23644
rect 30190 23604 30196 23656
rect 30248 23644 30254 23656
rect 31036 23644 31064 23684
rect 31846 23672 31852 23684
rect 31904 23672 31910 23724
rect 32122 23712 32128 23724
rect 32083 23684 32128 23712
rect 32122 23672 32128 23684
rect 32180 23672 32186 23724
rect 32232 23712 32260 23820
rect 32306 23808 32312 23860
rect 32364 23848 32370 23860
rect 32364 23820 32444 23848
rect 32364 23808 32370 23820
rect 32416 23780 32444 23820
rect 32490 23808 32496 23860
rect 32548 23848 32554 23860
rect 34701 23851 34759 23857
rect 34701 23848 34713 23851
rect 32548 23820 34713 23848
rect 32548 23808 32554 23820
rect 34701 23817 34713 23820
rect 34747 23848 34759 23851
rect 34790 23848 34796 23860
rect 34747 23820 34796 23848
rect 34747 23817 34759 23820
rect 34701 23811 34759 23817
rect 34790 23808 34796 23820
rect 34848 23808 34854 23860
rect 35894 23808 35900 23860
rect 35952 23848 35958 23860
rect 38473 23851 38531 23857
rect 38473 23848 38485 23851
rect 35952 23820 38485 23848
rect 35952 23808 35958 23820
rect 38473 23817 38485 23820
rect 38519 23817 38531 23851
rect 38473 23811 38531 23817
rect 32416 23752 35848 23780
rect 32309 23715 32367 23721
rect 32309 23712 32321 23715
rect 32232 23684 32321 23712
rect 32309 23681 32321 23684
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 32401 23715 32459 23721
rect 32401 23681 32413 23715
rect 32447 23712 32459 23715
rect 32447 23684 32628 23712
rect 32447 23681 32459 23684
rect 32401 23675 32459 23681
rect 30248 23616 31064 23644
rect 30248 23604 30254 23616
rect 31110 23604 31116 23656
rect 31168 23644 31174 23656
rect 32493 23647 32551 23653
rect 32493 23644 32505 23647
rect 31168 23616 32505 23644
rect 31168 23604 31174 23616
rect 32493 23613 32505 23616
rect 32539 23613 32551 23647
rect 32600 23644 32628 23684
rect 32674 23672 32680 23724
rect 32732 23712 32738 23724
rect 32732 23684 32777 23712
rect 32732 23672 32738 23684
rect 32858 23672 32864 23724
rect 32916 23712 32922 23724
rect 34698 23712 34704 23724
rect 32916 23684 34704 23712
rect 32916 23672 32922 23684
rect 34698 23672 34704 23684
rect 34756 23672 34762 23724
rect 35434 23712 35440 23724
rect 35395 23684 35440 23712
rect 35434 23672 35440 23684
rect 35492 23672 35498 23724
rect 35820 23712 35848 23752
rect 36170 23740 36176 23792
rect 36228 23780 36234 23792
rect 36228 23752 37780 23780
rect 36228 23740 36234 23752
rect 36354 23712 36360 23724
rect 35820 23684 36360 23712
rect 36354 23672 36360 23684
rect 36412 23672 36418 23724
rect 36538 23712 36544 23724
rect 36499 23684 36544 23712
rect 36538 23672 36544 23684
rect 36596 23672 36602 23724
rect 36722 23712 36728 23724
rect 36683 23684 36728 23712
rect 36722 23672 36728 23684
rect 36780 23672 36786 23724
rect 37550 23712 37556 23724
rect 37511 23684 37556 23712
rect 37550 23672 37556 23684
rect 37608 23672 37614 23724
rect 37752 23721 37780 23752
rect 38304 23752 41414 23780
rect 37645 23715 37703 23721
rect 37645 23681 37657 23715
rect 37691 23681 37703 23715
rect 37645 23675 37703 23681
rect 37737 23715 37795 23721
rect 37737 23681 37749 23715
rect 37783 23681 37795 23715
rect 37918 23712 37924 23724
rect 37879 23684 37924 23712
rect 37737 23675 37795 23681
rect 33870 23644 33876 23656
rect 32600 23616 33876 23644
rect 32493 23607 32551 23613
rect 33870 23604 33876 23616
rect 33928 23604 33934 23656
rect 35529 23647 35587 23653
rect 35529 23613 35541 23647
rect 35575 23644 35587 23647
rect 36740 23644 36768 23672
rect 37274 23644 37280 23656
rect 35575 23616 36768 23644
rect 37235 23616 37280 23644
rect 35575 23613 35587 23616
rect 35529 23607 35587 23613
rect 37274 23604 37280 23616
rect 37332 23604 37338 23656
rect 37660 23644 37688 23675
rect 37918 23672 37924 23684
rect 37976 23672 37982 23724
rect 38304 23644 38332 23752
rect 38381 23715 38439 23721
rect 38381 23681 38393 23715
rect 38427 23681 38439 23715
rect 38562 23712 38568 23724
rect 38523 23684 38568 23712
rect 38381 23675 38439 23681
rect 37660 23616 38332 23644
rect 28810 23576 28816 23588
rect 24136 23548 28816 23576
rect 28810 23536 28816 23548
rect 28868 23536 28874 23588
rect 32214 23576 32220 23588
rect 30852 23548 32220 23576
rect 30852 23508 30880 23548
rect 32214 23536 32220 23548
rect 32272 23536 32278 23588
rect 32324 23548 35848 23576
rect 23808 23480 30880 23508
rect 23808 23468 23814 23480
rect 31754 23468 31760 23520
rect 31812 23508 31818 23520
rect 32324 23508 32352 23548
rect 31812 23480 32352 23508
rect 31812 23468 31818 23480
rect 32398 23468 32404 23520
rect 32456 23508 32462 23520
rect 32861 23511 32919 23517
rect 32861 23508 32873 23511
rect 32456 23480 32873 23508
rect 32456 23468 32462 23480
rect 32861 23477 32873 23480
rect 32907 23477 32919 23511
rect 35710 23508 35716 23520
rect 35671 23480 35716 23508
rect 32861 23471 32919 23477
rect 35710 23468 35716 23480
rect 35768 23468 35774 23520
rect 35820 23508 35848 23548
rect 36354 23536 36360 23588
rect 36412 23576 36418 23588
rect 38396 23576 38424 23675
rect 38562 23672 38568 23684
rect 38620 23672 38626 23724
rect 41386 23644 41414 23752
rect 45186 23712 45192 23724
rect 45147 23684 45192 23712
rect 45186 23672 45192 23684
rect 45244 23672 45250 23724
rect 47578 23712 47584 23724
rect 47539 23684 47584 23712
rect 47578 23672 47584 23684
rect 47636 23672 47642 23724
rect 44082 23644 44088 23656
rect 41386 23616 44088 23644
rect 44082 23604 44088 23616
rect 44140 23604 44146 23656
rect 45373 23647 45431 23653
rect 45373 23613 45385 23647
rect 45419 23644 45431 23647
rect 46566 23644 46572 23656
rect 45419 23616 46572 23644
rect 45419 23613 45431 23616
rect 45373 23607 45431 23613
rect 46566 23604 46572 23616
rect 46624 23604 46630 23656
rect 46842 23644 46848 23656
rect 46803 23616 46848 23644
rect 46842 23604 46848 23616
rect 46900 23604 46906 23656
rect 47946 23576 47952 23588
rect 36412 23548 38424 23576
rect 41386 23548 47952 23576
rect 36412 23536 36418 23548
rect 41386 23508 41414 23548
rect 47946 23536 47952 23548
rect 48004 23536 48010 23588
rect 47670 23508 47676 23520
rect 35820 23480 41414 23508
rect 47631 23480 47676 23508
rect 47670 23468 47676 23480
rect 47728 23468 47734 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 14458 23264 14464 23316
rect 14516 23304 14522 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14516 23276 14657 23304
rect 14516 23264 14522 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 19334 23304 19340 23316
rect 19295 23276 19340 23304
rect 14645 23267 14703 23273
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 23750 23304 23756 23316
rect 23711 23276 23756 23304
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 26970 23264 26976 23316
rect 27028 23304 27034 23316
rect 27065 23307 27123 23313
rect 27065 23304 27077 23307
rect 27028 23276 27077 23304
rect 27028 23264 27034 23276
rect 27065 23273 27077 23276
rect 27111 23304 27123 23307
rect 27525 23307 27583 23313
rect 27525 23304 27537 23307
rect 27111 23276 27537 23304
rect 27111 23273 27123 23276
rect 27065 23267 27123 23273
rect 27525 23273 27537 23276
rect 27571 23273 27583 23307
rect 27525 23267 27583 23273
rect 27985 23307 28043 23313
rect 27985 23273 27997 23307
rect 28031 23304 28043 23307
rect 28902 23304 28908 23316
rect 28031 23276 28908 23304
rect 28031 23273 28043 23276
rect 27985 23267 28043 23273
rect 28902 23264 28908 23276
rect 28960 23264 28966 23316
rect 30282 23304 30288 23316
rect 30243 23276 30288 23304
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 31202 23304 31208 23316
rect 31163 23276 31208 23304
rect 31202 23264 31208 23276
rect 31260 23264 31266 23316
rect 31846 23264 31852 23316
rect 31904 23304 31910 23316
rect 36446 23304 36452 23316
rect 31904 23276 36452 23304
rect 31904 23264 31910 23276
rect 36446 23264 36452 23276
rect 36504 23264 36510 23316
rect 38473 23307 38531 23313
rect 38473 23273 38485 23307
rect 38519 23304 38531 23307
rect 38562 23304 38568 23316
rect 38519 23276 38568 23304
rect 38519 23273 38531 23276
rect 38473 23267 38531 23273
rect 38562 23264 38568 23276
rect 38620 23264 38626 23316
rect 2746 23208 17080 23236
rect 14 22992 20 23044
rect 72 23032 78 23044
rect 2746 23032 2774 23208
rect 14366 23168 14372 23180
rect 11440 23140 14228 23168
rect 14327 23140 14372 23168
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 11330 23100 11336 23112
rect 10459 23072 11336 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 72 23004 2774 23032
rect 72 22992 78 23004
rect 9950 22992 9956 23044
rect 10008 23032 10014 23044
rect 10781 23035 10839 23041
rect 10781 23032 10793 23035
rect 10008 23004 10793 23032
rect 10008 22992 10014 23004
rect 10781 23001 10793 23004
rect 10827 23032 10839 23035
rect 11440 23032 11468 23140
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 10827 23004 11468 23032
rect 10827 23001 10839 23004
rect 10781 22995 10839 23001
rect 10318 22924 10324 22976
rect 10376 22964 10382 22976
rect 10962 22964 10968 22976
rect 10376 22936 10968 22964
rect 10376 22924 10382 22936
rect 10962 22924 10968 22936
rect 11020 22964 11026 22976
rect 11532 22964 11560 23063
rect 12360 23032 12388 23063
rect 12802 23060 12808 23112
rect 12860 23100 12866 23112
rect 13265 23103 13323 23109
rect 13265 23100 13277 23103
rect 12860 23072 13277 23100
rect 12860 23060 12866 23072
rect 13265 23069 13277 23072
rect 13311 23100 13323 23103
rect 13354 23100 13360 23112
rect 13311 23072 13360 23100
rect 13311 23069 13323 23072
rect 13265 23063 13323 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 14200 23032 14228 23140
rect 14366 23128 14372 23140
rect 14424 23128 14430 23180
rect 15194 23168 15200 23180
rect 14476 23140 15200 23168
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14476 23100 14504 23140
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 16758 23168 16764 23180
rect 16719 23140 16764 23168
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 17052 23177 17080 23208
rect 17037 23171 17095 23177
rect 17037 23137 17049 23171
rect 17083 23137 17095 23171
rect 22002 23168 22008 23180
rect 21963 23140 22008 23168
rect 17037 23131 17095 23137
rect 22002 23128 22008 23140
rect 22060 23168 22066 23180
rect 22370 23168 22376 23180
rect 22060 23140 22376 23168
rect 22060 23128 22066 23140
rect 22370 23128 22376 23140
rect 22428 23168 22434 23180
rect 25317 23171 25375 23177
rect 25317 23168 25329 23171
rect 22428 23140 25329 23168
rect 22428 23128 22434 23140
rect 25317 23137 25329 23140
rect 25363 23137 25375 23171
rect 25590 23168 25596 23180
rect 25551 23140 25596 23168
rect 25317 23131 25375 23137
rect 25590 23128 25596 23140
rect 25648 23128 25654 23180
rect 26786 23128 26792 23180
rect 26844 23168 26850 23180
rect 30374 23168 30380 23180
rect 26844 23140 27844 23168
rect 30287 23140 30380 23168
rect 26844 23128 26850 23140
rect 15102 23100 15108 23112
rect 14323 23072 14504 23100
rect 15063 23072 15108 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23100 19303 23103
rect 19978 23100 19984 23112
rect 19291 23072 19984 23100
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 16592 23032 16620 23063
rect 19978 23060 19984 23072
rect 20036 23100 20042 23112
rect 20530 23100 20536 23112
rect 20036 23072 20536 23100
rect 20036 23060 20042 23072
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20714 23100 20720 23112
rect 20671 23072 20720 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 27706 23100 27712 23112
rect 27667 23072 27712 23100
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 27816 23109 27844 23140
rect 30300 23109 30328 23140
rect 30374 23128 30380 23140
rect 30432 23168 30438 23180
rect 31662 23168 31668 23180
rect 30432 23140 31668 23168
rect 30432 23128 30438 23140
rect 31662 23128 31668 23140
rect 31720 23128 31726 23180
rect 34790 23128 34796 23180
rect 34848 23168 34854 23180
rect 35253 23171 35311 23177
rect 35253 23168 35265 23171
rect 34848 23140 35265 23168
rect 34848 23128 34854 23140
rect 35253 23137 35265 23140
rect 35299 23137 35311 23171
rect 35253 23131 35311 23137
rect 46477 23171 46535 23177
rect 46477 23137 46489 23171
rect 46523 23168 46535 23171
rect 47670 23168 47676 23180
rect 46523 23140 47676 23168
rect 46523 23137 46535 23140
rect 46477 23131 46535 23137
rect 47670 23128 47676 23140
rect 47728 23128 47734 23180
rect 27801 23103 27859 23109
rect 27801 23069 27813 23103
rect 27847 23069 27859 23103
rect 27801 23063 27859 23069
rect 30285 23103 30343 23109
rect 30285 23069 30297 23103
rect 30331 23069 30343 23103
rect 30285 23063 30343 23069
rect 30466 23060 30472 23112
rect 30524 23100 30530 23112
rect 30650 23100 30656 23112
rect 30524 23072 30656 23100
rect 30524 23060 30530 23072
rect 30650 23060 30656 23072
rect 30708 23060 30714 23112
rect 31113 23103 31171 23109
rect 31113 23069 31125 23103
rect 31159 23100 31171 23103
rect 32953 23103 33011 23109
rect 32953 23100 32965 23103
rect 31159 23072 32965 23100
rect 31159 23069 31171 23072
rect 31113 23063 31171 23069
rect 32953 23069 32965 23072
rect 32999 23100 33011 23103
rect 33226 23100 33232 23112
rect 32999 23072 33232 23100
rect 32999 23069 33011 23072
rect 32953 23063 33011 23069
rect 33226 23060 33232 23072
rect 33284 23060 33290 23112
rect 34698 23060 34704 23112
rect 34756 23100 34762 23112
rect 36725 23103 36783 23109
rect 36725 23100 36737 23103
rect 34756 23072 36737 23100
rect 34756 23060 34762 23072
rect 36725 23069 36737 23072
rect 36771 23069 36783 23103
rect 41414 23100 41420 23112
rect 41375 23072 41420 23100
rect 36725 23063 36783 23069
rect 41414 23060 41420 23072
rect 41472 23060 41478 23112
rect 42153 23103 42211 23109
rect 42153 23069 42165 23103
rect 42199 23069 42211 23103
rect 46290 23100 46296 23112
rect 46251 23072 46296 23100
rect 42153 23063 42211 23069
rect 18414 23032 18420 23044
rect 12360 23004 13492 23032
rect 14200 23004 15424 23032
rect 16592 23004 18420 23032
rect 11698 22964 11704 22976
rect 11020 22936 11560 22964
rect 11659 22936 11704 22964
rect 11020 22924 11026 22936
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 12434 22924 12440 22976
rect 12492 22964 12498 22976
rect 13464 22973 13492 23004
rect 13449 22967 13507 22973
rect 12492 22936 12537 22964
rect 12492 22924 12498 22936
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 14182 22964 14188 22976
rect 13495 22936 14188 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14182 22924 14188 22936
rect 14240 22924 14246 22976
rect 15286 22964 15292 22976
rect 15247 22936 15292 22964
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 15396 22964 15424 23004
rect 18414 22992 18420 23004
rect 18472 22992 18478 23044
rect 22278 23032 22284 23044
rect 22239 23004 22284 23032
rect 22278 22992 22284 23004
rect 22336 22992 22342 23044
rect 26326 22992 26332 23044
rect 26384 22992 26390 23044
rect 27062 22992 27068 23044
rect 27120 23032 27126 23044
rect 27525 23035 27583 23041
rect 27525 23032 27537 23035
rect 27120 23004 27537 23032
rect 27120 22992 27126 23004
rect 27525 23001 27537 23004
rect 27571 23001 27583 23035
rect 27525 22995 27583 23001
rect 35161 23035 35219 23041
rect 35161 23001 35173 23035
rect 35207 23032 35219 23035
rect 35710 23032 35716 23044
rect 35207 23004 35716 23032
rect 35207 23001 35219 23004
rect 35161 22995 35219 23001
rect 35710 22992 35716 23004
rect 35768 22992 35774 23044
rect 37001 23035 37059 23041
rect 37001 23001 37013 23035
rect 37047 23032 37059 23035
rect 37274 23032 37280 23044
rect 37047 23004 37280 23032
rect 37047 23001 37059 23004
rect 37001 22995 37059 23001
rect 37274 22992 37280 23004
rect 37332 22992 37338 23044
rect 37458 22992 37464 23044
rect 37516 22992 37522 23044
rect 41322 22992 41328 23044
rect 41380 23032 41386 23044
rect 42168 23032 42196 23063
rect 46290 23060 46296 23072
rect 46348 23060 46354 23112
rect 41380 23004 42196 23032
rect 42429 23035 42487 23041
rect 41380 22992 41386 23004
rect 42429 23001 42441 23035
rect 42475 23032 42487 23035
rect 47118 23032 47124 23044
rect 42475 23004 47124 23032
rect 42475 23001 42487 23004
rect 42429 22995 42487 23001
rect 47118 22992 47124 23004
rect 47176 22992 47182 23044
rect 48133 23035 48191 23041
rect 48133 23001 48145 23035
rect 48179 23032 48191 23035
rect 48222 23032 48228 23044
rect 48179 23004 48228 23032
rect 48179 23001 48191 23004
rect 48133 22995 48191 23001
rect 48222 22992 48228 23004
rect 48280 22992 48286 23044
rect 19058 22964 19064 22976
rect 15396 22936 19064 22964
rect 19058 22924 19064 22936
rect 19116 22924 19122 22976
rect 20438 22964 20444 22976
rect 20399 22936 20444 22964
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 33045 22967 33103 22973
rect 33045 22933 33057 22967
rect 33091 22964 33103 22967
rect 33134 22964 33140 22976
rect 33091 22936 33140 22964
rect 33091 22933 33103 22936
rect 33045 22927 33103 22933
rect 33134 22924 33140 22936
rect 33192 22924 33198 22976
rect 34606 22924 34612 22976
rect 34664 22964 34670 22976
rect 34701 22967 34759 22973
rect 34701 22964 34713 22967
rect 34664 22936 34713 22964
rect 34664 22924 34670 22936
rect 34701 22933 34713 22936
rect 34747 22933 34759 22967
rect 34701 22927 34759 22933
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 35069 22967 35127 22973
rect 35069 22964 35081 22967
rect 34848 22936 35081 22964
rect 34848 22924 34854 22936
rect 35069 22933 35081 22936
rect 35115 22933 35127 22967
rect 41598 22964 41604 22976
rect 41559 22936 41604 22964
rect 35069 22927 35127 22933
rect 41598 22924 41604 22936
rect 41656 22924 41662 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 13078 22760 13084 22772
rect 8680 22732 13084 22760
rect 8018 22624 8024 22636
rect 7979 22596 8024 22624
rect 8018 22584 8024 22596
rect 8076 22584 8082 22636
rect 8680 22633 8708 22732
rect 13078 22720 13084 22732
rect 13136 22760 13142 22772
rect 13265 22763 13323 22769
rect 13265 22760 13277 22763
rect 13136 22732 13277 22760
rect 13136 22720 13142 22732
rect 13265 22729 13277 22732
rect 13311 22729 13323 22763
rect 14274 22760 14280 22772
rect 14235 22732 14280 22760
rect 13265 22723 13323 22729
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 18414 22760 18420 22772
rect 18375 22732 18420 22760
rect 18414 22720 18420 22732
rect 18472 22720 18478 22772
rect 22066 22732 46520 22760
rect 11698 22692 11704 22704
rect 11532 22664 11704 22692
rect 11532 22633 11560 22664
rect 11698 22652 11704 22664
rect 11756 22652 11762 22704
rect 12434 22652 12440 22704
rect 12492 22652 12498 22704
rect 13354 22652 13360 22704
rect 13412 22692 13418 22704
rect 13412 22664 15884 22692
rect 13412 22652 13418 22664
rect 8665 22627 8723 22633
rect 8665 22593 8677 22627
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22593 11575 22627
rect 14182 22624 14188 22636
rect 14095 22596 14188 22624
rect 11517 22587 11575 22593
rect 14182 22584 14188 22596
rect 14240 22624 14246 22636
rect 14734 22624 14740 22636
rect 14240 22596 14740 22624
rect 14240 22584 14246 22596
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 15856 22633 15884 22664
rect 16850 22652 16856 22704
rect 16908 22692 16914 22704
rect 16945 22695 17003 22701
rect 16945 22692 16957 22695
rect 16908 22664 16957 22692
rect 16908 22652 16914 22664
rect 16945 22661 16957 22664
rect 16991 22661 17003 22695
rect 18969 22695 19027 22701
rect 18969 22692 18981 22695
rect 18170 22664 18981 22692
rect 16945 22655 17003 22661
rect 18969 22661 18981 22664
rect 19015 22661 19027 22695
rect 18969 22655 19027 22661
rect 19058 22652 19064 22704
rect 19116 22692 19122 22704
rect 22066 22692 22094 22732
rect 23382 22692 23388 22704
rect 19116 22664 22094 22692
rect 23343 22664 23388 22692
rect 19116 22652 19122 22664
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 26326 22692 26332 22704
rect 26287 22664 26332 22692
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 27614 22692 27620 22704
rect 26804 22664 27620 22692
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 18877 22627 18935 22633
rect 18877 22593 18889 22627
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 20530 22624 20536 22636
rect 20491 22596 20536 22624
rect 19705 22587 19763 22593
rect 8846 22556 8852 22568
rect 8807 22528 8852 22556
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 9125 22559 9183 22565
rect 9125 22525 9137 22559
rect 9171 22525 9183 22559
rect 11790 22556 11796 22568
rect 11751 22528 11796 22556
rect 9125 22519 9183 22525
rect 3786 22448 3792 22500
rect 3844 22488 3850 22500
rect 9140 22488 9168 22519
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 16666 22556 16672 22568
rect 16627 22528 16672 22556
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 18892 22556 18920 22587
rect 16776 22528 18920 22556
rect 3844 22460 9168 22488
rect 16025 22491 16083 22497
rect 3844 22448 3850 22460
rect 16025 22457 16037 22491
rect 16071 22488 16083 22491
rect 16574 22488 16580 22500
rect 16071 22460 16580 22488
rect 16071 22457 16083 22460
rect 16025 22451 16083 22457
rect 16574 22448 16580 22460
rect 16632 22488 16638 22500
rect 16776 22488 16804 22528
rect 19720 22500 19748 22587
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 23106 22584 23112 22636
rect 23164 22624 23170 22636
rect 23293 22627 23351 22633
rect 23293 22624 23305 22627
rect 23164 22596 23305 22624
rect 23164 22584 23170 22596
rect 23293 22593 23305 22596
rect 23339 22593 23351 22627
rect 23293 22587 23351 22593
rect 26142 22584 26148 22636
rect 26200 22624 26206 22636
rect 26237 22627 26295 22633
rect 26237 22624 26249 22627
rect 26200 22596 26249 22624
rect 26200 22584 26206 22596
rect 26237 22593 26249 22596
rect 26283 22624 26295 22627
rect 26804 22624 26832 22664
rect 27614 22652 27620 22664
rect 27672 22692 27678 22704
rect 28166 22692 28172 22704
rect 27672 22664 28172 22692
rect 27672 22652 27678 22664
rect 28166 22652 28172 22664
rect 28224 22652 28230 22704
rect 32398 22692 32404 22704
rect 32359 22664 32404 22692
rect 32398 22652 32404 22664
rect 32456 22652 32462 22704
rect 33134 22652 33140 22704
rect 33192 22652 33198 22704
rect 34606 22652 34612 22704
rect 34664 22692 34670 22704
rect 35161 22695 35219 22701
rect 35161 22692 35173 22695
rect 34664 22664 35173 22692
rect 34664 22652 34670 22664
rect 35161 22661 35173 22664
rect 35207 22661 35219 22695
rect 36446 22692 36452 22704
rect 35161 22655 35219 22661
rect 35544 22664 36452 22692
rect 26283 22596 26832 22624
rect 26973 22627 27031 22633
rect 26283 22593 26295 22596
rect 26237 22587 26295 22593
rect 26973 22593 26985 22627
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 26786 22516 26792 22568
rect 26844 22556 26850 22568
rect 26988 22556 27016 22587
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 35069 22627 35127 22633
rect 27120 22596 27165 22624
rect 27120 22584 27126 22596
rect 35069 22593 35081 22627
rect 35115 22624 35127 22627
rect 35434 22624 35440 22636
rect 35115 22596 35440 22624
rect 35115 22593 35127 22596
rect 35069 22587 35127 22593
rect 35434 22584 35440 22596
rect 35492 22584 35498 22636
rect 26844 22528 27016 22556
rect 27249 22559 27307 22565
rect 26844 22516 26850 22528
rect 27249 22525 27261 22559
rect 27295 22556 27307 22559
rect 27706 22556 27712 22568
rect 27295 22528 27712 22556
rect 27295 22525 27307 22528
rect 27249 22519 27307 22525
rect 27706 22516 27712 22528
rect 27764 22516 27770 22568
rect 32122 22556 32128 22568
rect 32083 22528 32128 22556
rect 32122 22516 32128 22528
rect 32180 22516 32186 22568
rect 33870 22556 33876 22568
rect 33831 22528 33876 22556
rect 33870 22516 33876 22528
rect 33928 22516 33934 22568
rect 35345 22559 35403 22565
rect 35345 22525 35357 22559
rect 35391 22556 35403 22559
rect 35544 22556 35572 22664
rect 36446 22652 36452 22664
rect 36504 22652 36510 22704
rect 37369 22695 37427 22701
rect 37369 22661 37381 22695
rect 37415 22692 37427 22695
rect 37458 22692 37464 22704
rect 37415 22664 37464 22692
rect 37415 22661 37427 22664
rect 37369 22655 37427 22661
rect 37458 22652 37464 22664
rect 37516 22652 37522 22704
rect 41414 22652 41420 22704
rect 41472 22692 41478 22704
rect 41509 22695 41567 22701
rect 41509 22692 41521 22695
rect 41472 22664 41521 22692
rect 41472 22652 41478 22664
rect 41509 22661 41521 22664
rect 41555 22661 41567 22695
rect 41509 22655 41567 22661
rect 45373 22695 45431 22701
rect 45373 22661 45385 22695
rect 45419 22692 45431 22695
rect 46014 22692 46020 22704
rect 45419 22664 46020 22692
rect 45419 22661 45431 22664
rect 45373 22655 45431 22661
rect 46014 22652 46020 22664
rect 46072 22652 46078 22704
rect 46492 22692 46520 22732
rect 46566 22720 46572 22772
rect 46624 22760 46630 22772
rect 47673 22763 47731 22769
rect 47673 22760 47685 22763
rect 46624 22732 47685 22760
rect 46624 22720 46630 22732
rect 47673 22729 47685 22732
rect 47719 22729 47731 22763
rect 47673 22723 47731 22729
rect 46492 22664 47624 22692
rect 47596 22636 47624 22664
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22593 36139 22627
rect 37274 22624 37280 22636
rect 37235 22596 37280 22624
rect 36081 22587 36139 22593
rect 35391 22528 35572 22556
rect 35391 22525 35403 22528
rect 35345 22519 35403 22525
rect 16632 22460 16804 22488
rect 16632 22448 16638 22460
rect 19702 22448 19708 22500
rect 19760 22488 19766 22500
rect 20898 22488 20904 22500
rect 19760 22460 20904 22488
rect 19760 22448 19766 22460
rect 20898 22448 20904 22460
rect 20956 22448 20962 22500
rect 26878 22448 26884 22500
rect 26936 22488 26942 22500
rect 26973 22491 27031 22497
rect 26973 22488 26985 22491
rect 26936 22460 26985 22488
rect 26936 22448 26942 22460
rect 26973 22457 26985 22460
rect 27019 22488 27031 22491
rect 27338 22488 27344 22500
rect 27019 22460 27344 22488
rect 27019 22457 27031 22460
rect 26973 22451 27031 22457
rect 27338 22448 27344 22460
rect 27396 22448 27402 22500
rect 34701 22491 34759 22497
rect 34701 22457 34713 22491
rect 34747 22488 34759 22491
rect 36096 22488 36124 22587
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 47578 22624 47584 22636
rect 47491 22596 47584 22624
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 42426 22556 42432 22568
rect 42387 22528 42432 22556
rect 42426 22516 42432 22528
rect 42484 22516 42490 22568
rect 42610 22556 42616 22568
rect 42571 22528 42616 22556
rect 42610 22516 42616 22528
rect 42668 22516 42674 22568
rect 43990 22556 43996 22568
rect 43951 22528 43996 22556
rect 43990 22516 43996 22528
rect 44048 22516 44054 22568
rect 45189 22559 45247 22565
rect 45189 22525 45201 22559
rect 45235 22556 45247 22559
rect 45235 22528 45554 22556
rect 45235 22525 45247 22528
rect 45189 22519 45247 22525
rect 34747 22460 36124 22488
rect 45526 22488 45554 22528
rect 45646 22516 45652 22568
rect 45704 22556 45710 22568
rect 47854 22556 47860 22568
rect 45704 22528 47860 22556
rect 45704 22516 45710 22528
rect 47854 22516 47860 22528
rect 47912 22516 47918 22568
rect 47394 22488 47400 22500
rect 45526 22460 47400 22488
rect 34747 22457 34759 22460
rect 34701 22451 34759 22457
rect 47394 22448 47400 22460
rect 47452 22448 47458 22500
rect 8113 22423 8171 22429
rect 8113 22389 8125 22423
rect 8159 22420 8171 22423
rect 9122 22420 9128 22432
rect 8159 22392 9128 22420
rect 8159 22389 8171 22392
rect 8113 22383 8171 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 19981 22423 20039 22429
rect 19981 22389 19993 22423
rect 20027 22420 20039 22423
rect 20162 22420 20168 22432
rect 20027 22392 20168 22420
rect 20027 22389 20039 22392
rect 19981 22383 20039 22389
rect 20162 22380 20168 22392
rect 20220 22380 20226 22432
rect 20717 22423 20775 22429
rect 20717 22389 20729 22423
rect 20763 22420 20775 22423
rect 20806 22420 20812 22432
rect 20763 22392 20812 22420
rect 20763 22389 20775 22392
rect 20717 22383 20775 22389
rect 20806 22380 20812 22392
rect 20864 22380 20870 22432
rect 35342 22380 35348 22432
rect 35400 22420 35406 22432
rect 35897 22423 35955 22429
rect 35897 22420 35909 22423
rect 35400 22392 35909 22420
rect 35400 22380 35406 22392
rect 35897 22389 35909 22392
rect 35943 22389 35955 22423
rect 35897 22383 35955 22389
rect 38194 22380 38200 22432
rect 38252 22420 38258 22432
rect 41322 22420 41328 22432
rect 38252 22392 41328 22420
rect 38252 22380 38258 22392
rect 41322 22380 41328 22392
rect 41380 22420 41386 22432
rect 41601 22423 41659 22429
rect 41601 22420 41613 22423
rect 41380 22392 41613 22420
rect 41380 22380 41386 22392
rect 41601 22389 41613 22392
rect 41647 22389 41659 22423
rect 41601 22383 41659 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8846 22216 8852 22228
rect 8343 22188 8852 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8846 22176 8852 22188
rect 8904 22176 8910 22228
rect 14829 22219 14887 22225
rect 14829 22185 14841 22219
rect 14875 22216 14887 22219
rect 15930 22216 15936 22228
rect 14875 22188 15936 22216
rect 14875 22185 14887 22188
rect 14829 22179 14887 22185
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 20790 22219 20848 22225
rect 20790 22216 20802 22219
rect 20496 22188 20802 22216
rect 20496 22176 20502 22188
rect 20790 22185 20802 22188
rect 20836 22185 20848 22219
rect 20790 22179 20848 22185
rect 20898 22176 20904 22228
rect 20956 22216 20962 22228
rect 38194 22216 38200 22228
rect 20956 22188 38200 22216
rect 20956 22176 20962 22188
rect 38194 22176 38200 22188
rect 38252 22176 38258 22228
rect 41417 22219 41475 22225
rect 41417 22185 41429 22219
rect 41463 22216 41475 22219
rect 42610 22216 42616 22228
rect 41463 22188 42616 22216
rect 41463 22185 41475 22188
rect 41417 22179 41475 22185
rect 42610 22176 42616 22188
rect 42668 22176 42674 22228
rect 46290 22176 46296 22228
rect 46348 22216 46354 22228
rect 47949 22219 48007 22225
rect 47949 22216 47961 22219
rect 46348 22188 47961 22216
rect 46348 22176 46354 22188
rect 47949 22185 47961 22188
rect 47995 22185 48007 22219
rect 47949 22179 48007 22185
rect 12618 22148 12624 22160
rect 12579 22120 12624 22148
rect 12618 22108 12624 22120
rect 12676 22108 12682 22160
rect 17034 22148 17040 22160
rect 16995 22120 17040 22148
rect 17034 22108 17040 22120
rect 17092 22108 17098 22160
rect 23109 22151 23167 22157
rect 23109 22148 23121 22151
rect 22480 22120 23121 22148
rect 8938 22080 8944 22092
rect 8899 22052 8944 22080
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 9122 22080 9128 22092
rect 9083 22052 9128 22080
rect 9122 22040 9128 22052
rect 9180 22040 9186 22092
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9401 22083 9459 22089
rect 9401 22080 9413 22083
rect 9364 22052 9413 22080
rect 9364 22040 9370 22052
rect 9401 22049 9413 22052
rect 9447 22049 9459 22083
rect 16117 22083 16175 22089
rect 9401 22043 9459 22049
rect 11348 22052 16068 22080
rect 11348 22024 11376 22052
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 21981 8263 22015
rect 11330 22012 11336 22024
rect 11291 21984 11336 22012
rect 8205 21975 8263 21981
rect 8220 21944 8248 21975
rect 11330 21972 11336 21984
rect 11388 21972 11394 22024
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13320 21984 14780 22012
rect 13320 21972 13326 21984
rect 8220 21916 9628 21944
rect 9600 21888 9628 21916
rect 12986 21904 12992 21956
rect 13044 21944 13050 21956
rect 14645 21947 14703 21953
rect 14645 21944 14657 21947
rect 13044 21916 14657 21944
rect 13044 21904 13050 21916
rect 14645 21913 14657 21916
rect 14691 21913 14703 21947
rect 14752 21944 14780 21984
rect 15286 21972 15292 22024
rect 15344 22012 15350 22024
rect 15562 22012 15568 22024
rect 15344 21984 15568 22012
rect 15344 21972 15350 21984
rect 15562 21972 15568 21984
rect 15620 22012 15626 22024
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15620 21984 15853 22012
rect 15620 21972 15626 21984
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 16040 22012 16068 22052
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 16666 22080 16672 22092
rect 16163 22052 16672 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 20533 22083 20591 22089
rect 20533 22049 20545 22083
rect 20579 22080 20591 22083
rect 20806 22080 20812 22092
rect 20579 22052 20812 22080
rect 20579 22049 20591 22052
rect 20533 22043 20591 22049
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 16040 21984 17785 22012
rect 15841 21975 15899 21981
rect 17773 21981 17785 21984
rect 17819 22012 17831 22015
rect 19702 22012 19708 22024
rect 17819 21984 19708 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 22480 22012 22508 22120
rect 23109 22117 23121 22120
rect 23155 22117 23167 22151
rect 27982 22148 27988 22160
rect 27943 22120 27988 22148
rect 23109 22111 23167 22117
rect 27982 22108 27988 22120
rect 28040 22108 28046 22160
rect 32766 22148 32772 22160
rect 32679 22120 32772 22148
rect 32766 22108 32772 22120
rect 32824 22148 32830 22160
rect 33226 22148 33232 22160
rect 32824 22120 33232 22148
rect 32824 22108 32830 22120
rect 33226 22108 33232 22120
rect 33284 22108 33290 22160
rect 26970 22080 26976 22092
rect 26160 22052 26976 22080
rect 26160 22021 26188 22052
rect 21942 21984 22508 22012
rect 23017 22015 23075 22021
rect 20073 21975 20131 21981
rect 23017 21981 23029 22015
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 26145 22015 26203 22021
rect 26145 21981 26157 22015
rect 26191 21981 26203 22015
rect 26145 21975 26203 21981
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 22012 26387 22015
rect 26602 22012 26608 22024
rect 26375 21984 26608 22012
rect 26375 21981 26387 21984
rect 26329 21975 26387 21981
rect 16669 21947 16727 21953
rect 16669 21944 16681 21947
rect 14752 21916 16681 21944
rect 14645 21907 14703 21913
rect 16669 21913 16681 21916
rect 16715 21944 16727 21947
rect 17218 21944 17224 21956
rect 16715 21916 17224 21944
rect 16715 21913 16727 21916
rect 16669 21907 16727 21913
rect 17218 21904 17224 21916
rect 17276 21904 17282 21956
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 18598 21944 18604 21956
rect 18371 21916 18604 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 18598 21904 18604 21916
rect 18656 21904 18662 21956
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 19904 21944 19932 21975
rect 19392 21916 19932 21944
rect 20088 21944 20116 21975
rect 20806 21944 20812 21956
rect 20088 21916 20812 21944
rect 19392 21904 19398 21916
rect 20806 21904 20812 21916
rect 20864 21904 20870 21956
rect 22557 21947 22615 21953
rect 22557 21913 22569 21947
rect 22603 21944 22615 21947
rect 22646 21944 22652 21956
rect 22603 21916 22652 21944
rect 22603 21913 22615 21916
rect 22557 21907 22615 21913
rect 5442 21836 5448 21888
rect 5500 21876 5506 21888
rect 9306 21876 9312 21888
rect 5500 21848 9312 21876
rect 5500 21836 5506 21848
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9582 21836 9588 21888
rect 9640 21876 9646 21888
rect 11425 21879 11483 21885
rect 11425 21876 11437 21879
rect 9640 21848 11437 21876
rect 9640 21836 9646 21848
rect 11425 21845 11437 21848
rect 11471 21845 11483 21879
rect 11425 21839 11483 21845
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 12805 21879 12863 21885
rect 12805 21876 12817 21879
rect 12032 21848 12817 21876
rect 12032 21836 12038 21848
rect 12805 21845 12817 21848
rect 12851 21845 12863 21879
rect 12805 21839 12863 21845
rect 14458 21836 14464 21888
rect 14516 21876 14522 21888
rect 14845 21879 14903 21885
rect 14845 21876 14857 21879
rect 14516 21848 14857 21876
rect 14516 21836 14522 21848
rect 14845 21845 14857 21848
rect 14891 21845 14903 21879
rect 14845 21839 14903 21845
rect 15013 21879 15071 21885
rect 15013 21845 15025 21879
rect 15059 21876 15071 21879
rect 15746 21876 15752 21888
rect 15059 21848 15752 21876
rect 15059 21845 15071 21848
rect 15013 21839 15071 21845
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 16942 21836 16948 21888
rect 17000 21876 17006 21888
rect 17129 21879 17187 21885
rect 17129 21876 17141 21879
rect 17000 21848 17141 21876
rect 17000 21836 17006 21848
rect 17129 21845 17141 21848
rect 17175 21845 17187 21879
rect 17129 21839 17187 21845
rect 20073 21879 20131 21885
rect 20073 21845 20085 21879
rect 20119 21876 20131 21879
rect 20438 21876 20444 21888
rect 20119 21848 20444 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20438 21836 20444 21848
rect 20496 21836 20502 21888
rect 20530 21836 20536 21888
rect 20588 21876 20594 21888
rect 22572 21876 22600 21907
rect 22646 21904 22652 21916
rect 22704 21904 22710 21956
rect 23032 21944 23060 21975
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 26804 22021 26832 22052
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 30466 22080 30472 22092
rect 27080 22052 29960 22080
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 21981 26847 22015
rect 27080 22012 27108 22052
rect 27706 22012 27712 22024
rect 26789 21975 26847 21981
rect 26896 21984 27108 22012
rect 27667 21984 27712 22012
rect 23106 21944 23112 21956
rect 23032 21916 23112 21944
rect 23106 21904 23112 21916
rect 23164 21944 23170 21956
rect 23382 21944 23388 21956
rect 23164 21916 23388 21944
rect 23164 21904 23170 21916
rect 23382 21904 23388 21916
rect 23440 21944 23446 21956
rect 26896 21944 26924 21984
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 21981 27859 22015
rect 27801 21975 27859 21981
rect 23440 21916 26924 21944
rect 23440 21904 23446 21916
rect 26970 21904 26976 21956
rect 27028 21944 27034 21956
rect 27816 21944 27844 21975
rect 28166 21972 28172 22024
rect 28224 22012 28230 22024
rect 28445 22015 28503 22021
rect 28445 22012 28457 22015
rect 28224 21984 28457 22012
rect 28224 21972 28230 21984
rect 28445 21981 28457 21984
rect 28491 21981 28503 22015
rect 29822 22012 29828 22024
rect 29783 21984 29828 22012
rect 28445 21975 28503 21981
rect 29822 21972 29828 21984
rect 29880 21972 29886 22024
rect 29178 21944 29184 21956
rect 27028 21916 27073 21944
rect 27172 21916 27844 21944
rect 28368 21916 29184 21944
rect 27028 21904 27034 21916
rect 27172 21888 27200 21916
rect 20588 21848 22600 21876
rect 26329 21879 26387 21885
rect 20588 21836 20594 21848
rect 26329 21845 26341 21879
rect 26375 21876 26387 21879
rect 26418 21876 26424 21888
rect 26375 21848 26424 21876
rect 26375 21845 26387 21848
rect 26329 21839 26387 21845
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 27154 21876 27160 21888
rect 27115 21848 27160 21876
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27246 21836 27252 21888
rect 27304 21876 27310 21888
rect 28368 21876 28396 21916
rect 29178 21904 29184 21916
rect 29236 21904 29242 21956
rect 29641 21947 29699 21953
rect 29641 21913 29653 21947
rect 29687 21944 29699 21947
rect 29730 21944 29736 21956
rect 29687 21916 29736 21944
rect 29687 21913 29699 21916
rect 29641 21907 29699 21913
rect 29730 21904 29736 21916
rect 29788 21904 29794 21956
rect 29932 21944 29960 22052
rect 30024 22052 30472 22080
rect 30024 22021 30052 22052
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 31726 22052 32076 22080
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 21981 30067 22015
rect 30009 21975 30067 21981
rect 30098 21972 30104 22024
rect 30156 22012 30162 22024
rect 30156 21984 30201 22012
rect 30156 21972 30162 21984
rect 31726 21944 31754 22052
rect 29932 21916 31754 21944
rect 28534 21876 28540 21888
rect 27304 21848 28396 21876
rect 28495 21848 28540 21876
rect 27304 21836 27310 21848
rect 28534 21836 28540 21848
rect 28592 21836 28598 21888
rect 29454 21836 29460 21888
rect 29512 21876 29518 21888
rect 30098 21876 30104 21888
rect 29512 21848 30104 21876
rect 29512 21836 29518 21848
rect 30098 21836 30104 21848
rect 30156 21836 30162 21888
rect 32048 21876 32076 22052
rect 32122 22040 32128 22092
rect 32180 22080 32186 22092
rect 33042 22080 33048 22092
rect 32180 22052 33048 22080
rect 32180 22040 32186 22052
rect 33042 22040 33048 22052
rect 33100 22080 33106 22092
rect 34698 22080 34704 22092
rect 33100 22052 34704 22080
rect 33100 22040 33106 22052
rect 34698 22040 34704 22052
rect 34756 22040 34762 22092
rect 34977 22083 35035 22089
rect 34977 22049 34989 22083
rect 35023 22080 35035 22083
rect 35342 22080 35348 22092
rect 35023 22052 35348 22080
rect 35023 22049 35035 22052
rect 34977 22043 35035 22049
rect 35342 22040 35348 22052
rect 35400 22040 35406 22092
rect 35434 22040 35440 22092
rect 35492 22080 35498 22092
rect 36449 22083 36507 22089
rect 36449 22080 36461 22083
rect 35492 22052 36461 22080
rect 35492 22040 35498 22052
rect 36449 22049 36461 22052
rect 36495 22049 36507 22083
rect 42702 22080 42708 22092
rect 42663 22052 42708 22080
rect 36449 22043 36507 22049
rect 42702 22040 42708 22052
rect 42760 22040 42766 22092
rect 46658 22080 46664 22092
rect 46619 22052 46664 22080
rect 46658 22040 46664 22052
rect 46716 22040 46722 22092
rect 32585 22015 32643 22021
rect 32585 21981 32597 22015
rect 32631 22012 32643 22015
rect 33413 22015 33471 22021
rect 33413 22012 33425 22015
rect 32631 21984 33425 22012
rect 32631 21981 32643 21984
rect 32585 21975 32643 21981
rect 33413 21981 33425 21984
rect 33459 22012 33471 22015
rect 33962 22012 33968 22024
rect 33459 21984 33968 22012
rect 33459 21981 33471 21984
rect 33413 21975 33471 21981
rect 33962 21972 33968 21984
rect 34020 21972 34026 22024
rect 38841 22015 38899 22021
rect 38841 21981 38853 22015
rect 38887 21981 38899 22015
rect 38841 21975 38899 21981
rect 41325 22015 41383 22021
rect 41325 21981 41337 22015
rect 41371 22012 41383 22015
rect 41598 22012 41604 22024
rect 41371 21984 41604 22012
rect 41371 21981 41383 21984
rect 41325 21975 41383 21981
rect 35618 21904 35624 21956
rect 35676 21904 35682 21956
rect 38856 21944 38884 21975
rect 41598 21972 41604 21984
rect 41656 22012 41662 22024
rect 42153 22015 42211 22021
rect 42153 22012 42165 22015
rect 41656 21984 42165 22012
rect 41656 21972 41662 21984
rect 42153 21981 42165 21984
rect 42199 22012 42211 22015
rect 42610 22012 42616 22024
rect 42199 21984 42616 22012
rect 42199 21981 42211 21984
rect 42153 21975 42211 21981
rect 42610 21972 42616 21984
rect 42668 21972 42674 22024
rect 45462 22012 45468 22024
rect 45423 21984 45468 22012
rect 45462 21972 45468 21984
rect 45520 21972 45526 22024
rect 42794 21944 42800 21956
rect 38856 21916 42800 21944
rect 42794 21904 42800 21916
rect 42852 21904 42858 21956
rect 45646 21944 45652 21956
rect 45607 21916 45652 21944
rect 45646 21904 45652 21916
rect 45704 21904 45710 21956
rect 33502 21876 33508 21888
rect 32048 21848 33508 21876
rect 33502 21836 33508 21848
rect 33560 21836 33566 21888
rect 38930 21876 38936 21888
rect 38891 21848 38936 21876
rect 38930 21836 38936 21848
rect 38988 21836 38994 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 11790 21672 11796 21684
rect 11751 21644 11796 21672
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12618 21672 12624 21684
rect 12579 21644 12624 21672
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 12989 21675 13047 21681
rect 12989 21672 13001 21675
rect 12952 21644 13001 21672
rect 12952 21632 12958 21644
rect 12989 21641 13001 21644
rect 13035 21641 13047 21675
rect 12989 21635 13047 21641
rect 16761 21675 16819 21681
rect 16761 21641 16773 21675
rect 16807 21672 16819 21675
rect 16850 21672 16856 21684
rect 16807 21644 16856 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 17034 21632 17040 21684
rect 17092 21672 17098 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 17092 21644 17417 21672
rect 17092 21632 17098 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 20772 21644 20821 21672
rect 20772 21632 20778 21644
rect 20809 21641 20821 21644
rect 20855 21641 20867 21675
rect 20809 21635 20867 21641
rect 26329 21675 26387 21681
rect 26329 21641 26341 21675
rect 26375 21672 26387 21675
rect 27154 21672 27160 21684
rect 26375 21644 27160 21672
rect 26375 21641 26387 21644
rect 26329 21635 26387 21641
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 29178 21672 29184 21684
rect 27264 21644 29184 21672
rect 3510 21564 3516 21616
rect 3568 21604 3574 21616
rect 15565 21607 15623 21613
rect 15565 21604 15577 21607
rect 3568 21576 15577 21604
rect 3568 21564 3574 21576
rect 15565 21573 15577 21576
rect 15611 21573 15623 21607
rect 18230 21604 18236 21616
rect 15565 21567 15623 21573
rect 17696 21576 18236 21604
rect 8754 21496 8760 21548
rect 8812 21536 8818 21548
rect 8849 21539 8907 21545
rect 8849 21536 8861 21539
rect 8812 21508 8861 21536
rect 8812 21496 8818 21508
rect 8849 21505 8861 21508
rect 8895 21505 8907 21539
rect 11974 21536 11980 21548
rect 11935 21508 11980 21536
rect 8849 21499 8907 21505
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21536 12863 21539
rect 12986 21536 12992 21548
rect 12851 21508 12992 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 13722 21536 13728 21548
rect 13096 21508 13728 21536
rect 9033 21471 9091 21477
rect 9033 21437 9045 21471
rect 9079 21468 9091 21471
rect 9122 21468 9128 21480
rect 9079 21440 9128 21468
rect 9079 21437 9091 21440
rect 9033 21431 9091 21437
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21437 9367 21471
rect 9309 21431 9367 21437
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 9324 21400 9352 21431
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12768 21440 12909 21468
rect 12768 21428 12774 21440
rect 12897 21437 12909 21440
rect 12943 21468 12955 21471
rect 13096 21468 13124 21508
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17696 21545 17724 21576
rect 18230 21564 18236 21576
rect 18288 21564 18294 21616
rect 18414 21604 18420 21616
rect 18375 21576 18420 21604
rect 18414 21564 18420 21576
rect 18472 21564 18478 21616
rect 18506 21564 18512 21616
rect 18564 21604 18570 21616
rect 18617 21607 18675 21613
rect 18617 21604 18629 21607
rect 18564 21576 18629 21604
rect 18564 21564 18570 21576
rect 18617 21573 18629 21576
rect 18663 21573 18675 21607
rect 18617 21567 18675 21573
rect 19797 21607 19855 21613
rect 19797 21573 19809 21607
rect 19843 21604 19855 21607
rect 19843 21576 20852 21604
rect 19843 21573 19855 21576
rect 19797 21567 19855 21573
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21536 17923 21539
rect 18432 21536 18460 21564
rect 20824 21548 20852 21576
rect 22646 21564 22652 21616
rect 22704 21604 22710 21616
rect 27264 21604 27292 21644
rect 29178 21632 29184 21644
rect 29236 21632 29242 21684
rect 32122 21672 32128 21684
rect 29656 21644 32128 21672
rect 22704 21576 27292 21604
rect 22704 21564 22710 21576
rect 28534 21564 28540 21616
rect 28592 21564 28598 21616
rect 19610 21536 19616 21548
rect 17911 21508 18460 21536
rect 19571 21508 19616 21536
rect 17911 21505 17923 21508
rect 17865 21499 17923 21505
rect 19610 21496 19616 21508
rect 19668 21496 19674 21548
rect 20438 21536 20444 21548
rect 20399 21508 20444 21536
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 12943 21440 13124 21468
rect 13173 21471 13231 21477
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13173 21437 13185 21471
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 6972 21372 9352 21400
rect 6972 21360 6978 21372
rect 13078 21360 13084 21412
rect 13136 21400 13142 21412
rect 13188 21400 13216 21431
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 13909 21471 13967 21477
rect 13320 21440 13365 21468
rect 13320 21428 13326 21440
rect 13909 21437 13921 21471
rect 13955 21468 13967 21471
rect 14918 21468 14924 21480
rect 13955 21440 14924 21468
rect 13955 21437 13967 21440
rect 13909 21431 13967 21437
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21468 17831 21471
rect 18322 21468 18328 21480
rect 17819 21440 18328 21468
rect 17819 21437 17831 21440
rect 17773 21431 17831 21437
rect 13136 21372 13216 21400
rect 17604 21400 17632 21431
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 19981 21471 20039 21477
rect 19981 21437 19993 21471
rect 20027 21468 20039 21471
rect 20640 21468 20668 21499
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22554 21536 22560 21548
rect 22515 21508 22560 21536
rect 22373 21499 22431 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 20027 21440 20668 21468
rect 20027 21437 20039 21440
rect 19981 21431 20039 21437
rect 21726 21428 21732 21480
rect 21784 21468 21790 21480
rect 23032 21468 23060 21499
rect 23382 21496 23388 21548
rect 23440 21536 23446 21548
rect 23661 21539 23719 21545
rect 23661 21536 23673 21539
rect 23440 21508 23673 21536
rect 23440 21496 23446 21508
rect 23661 21505 23673 21508
rect 23707 21505 23719 21539
rect 23661 21499 23719 21505
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21536 25375 21539
rect 26142 21536 26148 21548
rect 25363 21508 26148 21536
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 26142 21496 26148 21508
rect 26200 21496 26206 21548
rect 26418 21496 26424 21548
rect 26476 21536 26482 21548
rect 29656 21536 29684 21644
rect 32122 21632 32128 21644
rect 32180 21632 32186 21684
rect 35618 21672 35624 21684
rect 35579 21644 35624 21672
rect 35618 21632 35624 21644
rect 35676 21632 35682 21684
rect 44082 21632 44088 21684
rect 44140 21672 44146 21684
rect 44913 21675 44971 21681
rect 44913 21672 44925 21675
rect 44140 21644 44925 21672
rect 44140 21632 44146 21644
rect 44913 21641 44925 21644
rect 44959 21641 44971 21675
rect 45646 21672 45652 21684
rect 45607 21644 45652 21672
rect 44913 21635 44971 21641
rect 45646 21632 45652 21644
rect 45704 21632 45710 21684
rect 29730 21564 29736 21616
rect 29788 21604 29794 21616
rect 30101 21607 30159 21613
rect 30101 21604 30113 21607
rect 29788 21576 30113 21604
rect 29788 21564 29794 21576
rect 30101 21573 30113 21576
rect 30147 21573 30159 21607
rect 32217 21607 32275 21613
rect 32217 21604 32229 21607
rect 31326 21576 32229 21604
rect 30101 21567 30159 21573
rect 32217 21573 32229 21576
rect 32263 21573 32275 21607
rect 38930 21604 38936 21616
rect 38891 21576 38936 21604
rect 32217 21567 32275 21573
rect 38930 21564 38936 21576
rect 38988 21564 38994 21616
rect 42702 21564 42708 21616
rect 42760 21604 42766 21616
rect 42760 21576 47624 21604
rect 42760 21564 42766 21576
rect 29825 21539 29883 21545
rect 29825 21536 29837 21539
rect 26476 21508 26521 21536
rect 29656 21508 29837 21536
rect 26476 21496 26482 21508
rect 29825 21505 29837 21508
rect 29871 21505 29883 21539
rect 29825 21499 29883 21505
rect 32125 21539 32183 21545
rect 32125 21505 32137 21539
rect 32171 21536 32183 21539
rect 32766 21536 32772 21548
rect 32171 21508 32772 21536
rect 32171 21505 32183 21508
rect 32125 21499 32183 21505
rect 32766 21496 32772 21508
rect 32824 21496 32830 21548
rect 33502 21496 33508 21548
rect 33560 21536 33566 21548
rect 35529 21539 35587 21545
rect 35529 21536 35541 21539
rect 33560 21508 35541 21536
rect 33560 21496 33566 21508
rect 35529 21505 35541 21508
rect 35575 21536 35587 21539
rect 37274 21536 37280 21548
rect 35575 21508 37280 21536
rect 35575 21505 35587 21508
rect 35529 21499 35587 21505
rect 37274 21496 37280 21508
rect 37332 21496 37338 21548
rect 42610 21536 42616 21548
rect 42571 21508 42616 21536
rect 42610 21496 42616 21508
rect 42668 21496 42674 21548
rect 45097 21539 45155 21545
rect 45097 21505 45109 21539
rect 45143 21505 45155 21539
rect 45097 21499 45155 21505
rect 45557 21539 45615 21545
rect 45557 21505 45569 21539
rect 45603 21536 45615 21539
rect 45738 21536 45744 21548
rect 45603 21508 45744 21536
rect 45603 21505 45615 21508
rect 45557 21499 45615 21505
rect 21784 21440 23060 21468
rect 25961 21471 26019 21477
rect 21784 21428 21790 21440
rect 25961 21437 25973 21471
rect 26007 21468 26019 21471
rect 27246 21468 27252 21480
rect 26007 21440 27252 21468
rect 26007 21437 26019 21440
rect 25961 21431 26019 21437
rect 27246 21428 27252 21440
rect 27304 21428 27310 21480
rect 27522 21468 27528 21480
rect 27483 21440 27528 21468
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21468 27859 21471
rect 28258 21468 28264 21480
rect 27847 21440 28264 21468
rect 27847 21437 27859 21440
rect 27801 21431 27859 21437
rect 28258 21428 28264 21440
rect 28316 21428 28322 21480
rect 38749 21471 38807 21477
rect 38749 21468 38761 21471
rect 28828 21440 38761 21468
rect 18506 21400 18512 21412
rect 17604 21372 18512 21400
rect 13136 21360 13142 21372
rect 18506 21360 18512 21372
rect 18564 21360 18570 21412
rect 21450 21360 21456 21412
rect 21508 21400 21514 21412
rect 23014 21400 23020 21412
rect 21508 21372 23020 21400
rect 21508 21360 21514 21372
rect 23014 21360 23020 21372
rect 23072 21360 23078 21412
rect 23109 21403 23167 21409
rect 23109 21369 23121 21403
rect 23155 21400 23167 21403
rect 23155 21372 27660 21400
rect 23155 21369 23167 21372
rect 23109 21363 23167 21369
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 18601 21335 18659 21341
rect 18601 21332 18613 21335
rect 18288 21304 18613 21332
rect 18288 21292 18294 21304
rect 18601 21301 18613 21304
rect 18647 21301 18659 21335
rect 18782 21332 18788 21344
rect 18743 21304 18788 21332
rect 18601 21295 18659 21301
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 22370 21332 22376 21344
rect 22331 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 23750 21332 23756 21344
rect 23711 21304 23756 21332
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 25406 21332 25412 21344
rect 25367 21304 25412 21332
rect 25406 21292 25412 21304
rect 25464 21292 25470 21344
rect 26050 21292 26056 21344
rect 26108 21332 26114 21344
rect 26145 21335 26203 21341
rect 26145 21332 26157 21335
rect 26108 21304 26157 21332
rect 26108 21292 26114 21304
rect 26145 21301 26157 21304
rect 26191 21301 26203 21335
rect 27632 21332 27660 21372
rect 28828 21332 28856 21440
rect 38749 21437 38761 21440
rect 38795 21437 38807 21471
rect 38749 21431 38807 21437
rect 39114 21428 39120 21480
rect 39172 21468 39178 21480
rect 39209 21471 39267 21477
rect 39209 21468 39221 21471
rect 39172 21440 39221 21468
rect 39172 21428 39178 21440
rect 39209 21437 39221 21440
rect 39255 21437 39267 21471
rect 42794 21468 42800 21480
rect 42755 21440 42800 21468
rect 39209 21431 39267 21437
rect 42794 21428 42800 21440
rect 42852 21428 42858 21480
rect 45112 21468 45140 21499
rect 45738 21496 45744 21508
rect 45796 21496 45802 21548
rect 46198 21536 46204 21548
rect 46159 21508 46204 21536
rect 46198 21496 46204 21508
rect 46256 21496 46262 21548
rect 47486 21536 47492 21548
rect 46308 21508 47492 21536
rect 46106 21468 46112 21480
rect 45112 21440 46112 21468
rect 46106 21428 46112 21440
rect 46164 21428 46170 21480
rect 42812 21400 42840 21428
rect 43254 21400 43260 21412
rect 42812 21372 43260 21400
rect 43254 21360 43260 21372
rect 43312 21400 43318 21412
rect 43312 21372 45554 21400
rect 43312 21360 43318 21372
rect 27632 21304 28856 21332
rect 26145 21295 26203 21301
rect 28902 21292 28908 21344
rect 28960 21332 28966 21344
rect 29273 21335 29331 21341
rect 29273 21332 29285 21335
rect 28960 21304 29285 21332
rect 28960 21292 28966 21304
rect 29273 21301 29285 21304
rect 29319 21301 29331 21335
rect 29273 21295 29331 21301
rect 30466 21292 30472 21344
rect 30524 21332 30530 21344
rect 31573 21335 31631 21341
rect 31573 21332 31585 21335
rect 30524 21304 31585 21332
rect 30524 21292 30530 21304
rect 31573 21301 31585 21304
rect 31619 21301 31631 21335
rect 45526 21332 45554 21372
rect 46308 21332 46336 21508
rect 47486 21496 47492 21508
rect 47544 21496 47550 21548
rect 47596 21545 47624 21576
rect 47581 21539 47639 21545
rect 47581 21505 47593 21539
rect 47627 21505 47639 21539
rect 47581 21499 47639 21505
rect 46477 21471 46535 21477
rect 46477 21437 46489 21471
rect 46523 21468 46535 21471
rect 46658 21468 46664 21480
rect 46523 21440 46664 21468
rect 46523 21437 46535 21440
rect 46477 21431 46535 21437
rect 46658 21428 46664 21440
rect 46716 21428 46722 21480
rect 45526 21304 46336 21332
rect 31573 21295 31631 21301
rect 46474 21292 46480 21344
rect 46532 21332 46538 21344
rect 47673 21335 47731 21341
rect 47673 21332 47685 21335
rect 46532 21304 47685 21332
rect 46532 21292 46538 21304
rect 47673 21301 47685 21304
rect 47719 21301 47731 21335
rect 47673 21295 47731 21301
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 9122 21128 9128 21140
rect 9083 21100 9128 21128
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 12710 21128 12716 21140
rect 12671 21100 12716 21128
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 12952 21100 14289 21128
rect 12952 21088 12958 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 14458 21128 14464 21140
rect 14419 21100 14464 21128
rect 14277 21091 14335 21097
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14918 21088 14924 21140
rect 14976 21128 14982 21140
rect 15013 21131 15071 21137
rect 15013 21128 15025 21131
rect 14976 21100 15025 21128
rect 14976 21088 14982 21100
rect 15013 21097 15025 21100
rect 15059 21097 15071 21131
rect 17218 21128 17224 21140
rect 17179 21100 17224 21128
rect 15013 21091 15071 21097
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 21913 21131 21971 21137
rect 21913 21097 21925 21131
rect 21959 21128 21971 21131
rect 22186 21128 22192 21140
rect 21959 21100 22192 21128
rect 21959 21097 21971 21100
rect 21913 21091 21971 21097
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 23014 21088 23020 21140
rect 23072 21128 23078 21140
rect 28258 21128 28264 21140
rect 23072 21100 26188 21128
rect 28219 21100 28264 21128
rect 23072 21088 23078 21100
rect 21542 21020 21548 21072
rect 21600 21060 21606 21072
rect 26160 21060 26188 21100
rect 28258 21088 28264 21100
rect 28316 21088 28322 21140
rect 28350 21088 28356 21140
rect 28408 21128 28414 21140
rect 45462 21128 45468 21140
rect 28408 21100 45468 21128
rect 28408 21088 28414 21100
rect 45462 21088 45468 21100
rect 45520 21088 45526 21140
rect 21600 21032 24532 21060
rect 26160 21032 29040 21060
rect 21600 21020 21606 21032
rect 15930 20952 15936 21004
rect 15988 20992 15994 21004
rect 18782 20992 18788 21004
rect 15988 20964 18788 20992
rect 15988 20952 15994 20964
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 9033 20927 9091 20933
rect 9033 20924 9045 20927
rect 8352 20896 9045 20924
rect 8352 20884 8358 20896
rect 9033 20893 9045 20896
rect 9079 20924 9091 20927
rect 9582 20924 9588 20936
rect 9079 20896 9588 20924
rect 9079 20893 9091 20896
rect 9033 20887 9091 20893
rect 9582 20884 9588 20896
rect 9640 20924 9646 20936
rect 9677 20927 9735 20933
rect 9677 20924 9689 20927
rect 9640 20896 9689 20924
rect 9640 20884 9646 20896
rect 9677 20893 9689 20896
rect 9723 20893 9735 20927
rect 10318 20924 10324 20936
rect 10279 20896 10324 20924
rect 9677 20887 9735 20893
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20924 10471 20927
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 10459 20896 10977 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 15102 20924 15108 20936
rect 14967 20896 15108 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 17310 20924 17316 20936
rect 15611 20896 17316 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 17310 20884 17316 20896
rect 17368 20884 17374 20936
rect 17420 20933 17448 20964
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 20530 20992 20536 21004
rect 20491 20964 20536 20992
rect 20530 20952 20536 20964
rect 20588 20952 20594 21004
rect 21726 20992 21732 21004
rect 20640 20964 21732 20992
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20893 17463 20927
rect 17586 20924 17592 20936
rect 17547 20896 17592 20924
rect 17405 20887 17463 20893
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 17681 20927 17739 20933
rect 17681 20893 17693 20927
rect 17727 20893 17739 20927
rect 17681 20887 17739 20893
rect 18141 20927 18199 20933
rect 18141 20893 18153 20927
rect 18187 20924 18199 20927
rect 18506 20924 18512 20936
rect 18187 20896 18512 20924
rect 18187 20893 18199 20896
rect 18141 20887 18199 20893
rect 11238 20856 11244 20868
rect 11199 20828 11244 20856
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11698 20816 11704 20868
rect 11756 20816 11762 20868
rect 13722 20816 13728 20868
rect 13780 20856 13786 20868
rect 14093 20859 14151 20865
rect 14093 20856 14105 20859
rect 13780 20828 14105 20856
rect 13780 20816 13786 20828
rect 14093 20825 14105 20828
rect 14139 20825 14151 20859
rect 17696 20856 17724 20887
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 19392 20896 19901 20924
rect 19392 20884 19398 20896
rect 19889 20893 19901 20896
rect 19935 20924 19947 20927
rect 20640 20924 20668 20964
rect 21726 20952 21732 20964
rect 21784 20992 21790 21004
rect 21784 20964 22232 20992
rect 21784 20952 21790 20964
rect 20806 20924 20812 20936
rect 19935 20896 20668 20924
rect 20719 20896 20812 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 20806 20884 20812 20896
rect 20864 20924 20870 20936
rect 21818 20924 21824 20936
rect 20864 20896 21824 20924
rect 20864 20884 20870 20896
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 22002 20884 22008 20936
rect 22060 20924 22066 20936
rect 22204 20933 22232 20964
rect 22097 20927 22155 20933
rect 22097 20924 22109 20927
rect 22060 20896 22109 20924
rect 22060 20884 22066 20896
rect 22097 20893 22109 20896
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 22189 20927 22247 20933
rect 22189 20893 22201 20927
rect 22235 20893 22247 20927
rect 22189 20887 22247 20893
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 17696 20828 18368 20856
rect 14093 20819 14151 20825
rect 9766 20788 9772 20800
rect 9727 20760 9772 20788
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 14274 20748 14280 20800
rect 14332 20797 14338 20800
rect 14332 20791 14351 20797
rect 14339 20757 14351 20791
rect 14332 20751 14351 20757
rect 14332 20748 14338 20751
rect 15286 20748 15292 20800
rect 15344 20788 15350 20800
rect 15657 20791 15715 20797
rect 15657 20788 15669 20791
rect 15344 20760 15669 20788
rect 15344 20748 15350 20760
rect 15657 20757 15669 20760
rect 15703 20757 15715 20791
rect 15657 20751 15715 20757
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 18233 20791 18291 20797
rect 18233 20788 18245 20791
rect 18012 20760 18245 20788
rect 18012 20748 18018 20760
rect 18233 20757 18245 20760
rect 18279 20757 18291 20791
rect 18340 20788 18368 20828
rect 18414 20816 18420 20868
rect 18472 20856 18478 20868
rect 19610 20856 19616 20868
rect 18472 20828 19616 20856
rect 18472 20816 18478 20828
rect 19610 20816 19616 20828
rect 19668 20856 19674 20868
rect 19705 20859 19763 20865
rect 19705 20856 19717 20859
rect 19668 20828 19717 20856
rect 19668 20816 19674 20828
rect 19705 20825 19717 20828
rect 19751 20825 19763 20859
rect 20070 20856 20076 20868
rect 19705 20819 19763 20825
rect 19904 20828 20076 20856
rect 19904 20788 19932 20828
rect 20070 20816 20076 20828
rect 20128 20816 20134 20868
rect 20714 20816 20720 20868
rect 20772 20856 20778 20868
rect 21542 20856 21548 20868
rect 20772 20828 21548 20856
rect 20772 20816 20778 20828
rect 21542 20816 21548 20828
rect 21600 20856 21606 20868
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 21600 20828 21925 20856
rect 21600 20816 21606 20828
rect 21913 20825 21925 20828
rect 21959 20825 21971 20859
rect 22664 20856 22692 20887
rect 21913 20819 21971 20825
rect 22066 20828 22692 20856
rect 18340 20760 19932 20788
rect 18233 20751 18291 20757
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 22066 20788 22094 20828
rect 24504 20800 24532 21032
rect 24857 20995 24915 21001
rect 24857 20961 24869 20995
rect 24903 20992 24915 20995
rect 27522 20992 27528 21004
rect 24903 20964 27528 20992
rect 24903 20961 24915 20964
rect 24857 20955 24915 20961
rect 27522 20952 27528 20964
rect 27580 20952 27586 21004
rect 27614 20924 27620 20936
rect 27575 20896 27620 20924
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 27706 20884 27712 20936
rect 27764 20924 27770 20936
rect 27764 20896 27809 20924
rect 27764 20884 27770 20896
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 27948 20896 27993 20924
rect 27948 20884 27954 20896
rect 28074 20884 28080 20936
rect 28132 20933 28138 20936
rect 28132 20924 28140 20933
rect 28132 20896 28177 20924
rect 28132 20887 28140 20896
rect 28132 20884 28138 20887
rect 25130 20856 25136 20868
rect 25091 20828 25136 20856
rect 25130 20816 25136 20828
rect 25188 20816 25194 20868
rect 25406 20816 25412 20868
rect 25464 20856 25470 20868
rect 25464 20828 25622 20856
rect 26436 20828 26740 20856
rect 25464 20816 25470 20828
rect 20036 20760 22094 20788
rect 20036 20748 20042 20760
rect 22462 20748 22468 20800
rect 22520 20788 22526 20800
rect 22833 20791 22891 20797
rect 22833 20788 22845 20791
rect 22520 20760 22845 20788
rect 22520 20748 22526 20760
rect 22833 20757 22845 20760
rect 22879 20757 22891 20791
rect 22833 20751 22891 20757
rect 24486 20748 24492 20800
rect 24544 20788 24550 20800
rect 26436 20788 26464 20828
rect 26602 20788 26608 20800
rect 24544 20760 26464 20788
rect 26563 20760 26608 20788
rect 24544 20748 24550 20760
rect 26602 20748 26608 20760
rect 26660 20748 26666 20800
rect 26712 20788 26740 20828
rect 27798 20816 27804 20868
rect 27856 20856 27862 20868
rect 27985 20859 28043 20865
rect 27985 20856 27997 20859
rect 27856 20828 27997 20856
rect 27856 20816 27862 20828
rect 27985 20825 27997 20828
rect 28031 20856 28043 20859
rect 28902 20856 28908 20868
rect 28031 20828 28908 20856
rect 28031 20825 28043 20828
rect 27985 20819 28043 20825
rect 28902 20816 28908 20828
rect 28960 20816 28966 20868
rect 29012 20856 29040 21032
rect 29178 21020 29184 21072
rect 29236 21060 29242 21072
rect 42426 21060 42432 21072
rect 29236 21032 42432 21060
rect 29236 21020 29242 21032
rect 42426 21020 42432 21032
rect 42484 21020 42490 21072
rect 30374 20992 30380 21004
rect 30335 20964 30380 20992
rect 30374 20952 30380 20964
rect 30432 20952 30438 21004
rect 42061 20995 42119 21001
rect 42061 20992 42073 20995
rect 35866 20964 42073 20992
rect 30466 20924 30472 20936
rect 30427 20896 30472 20924
rect 30466 20884 30472 20896
rect 30524 20884 30530 20936
rect 35866 20856 35894 20964
rect 42061 20961 42073 20964
rect 42107 20992 42119 20995
rect 42518 20992 42524 21004
rect 42107 20964 42524 20992
rect 42107 20961 42119 20964
rect 42061 20955 42119 20961
rect 42518 20952 42524 20964
rect 42576 20952 42582 21004
rect 46474 20992 46480 21004
rect 46435 20964 46480 20992
rect 46474 20952 46480 20964
rect 46532 20952 46538 21004
rect 48130 20992 48136 21004
rect 48091 20964 48136 20992
rect 48130 20952 48136 20964
rect 48188 20952 48194 21004
rect 41877 20927 41935 20933
rect 41877 20893 41889 20927
rect 41923 20924 41935 20927
rect 42610 20924 42616 20936
rect 41923 20896 42616 20924
rect 41923 20893 41935 20896
rect 41877 20887 41935 20893
rect 42610 20884 42616 20896
rect 42668 20884 42674 20936
rect 45833 20927 45891 20933
rect 45833 20893 45845 20927
rect 45879 20924 45891 20927
rect 46293 20927 46351 20933
rect 46293 20924 46305 20927
rect 45879 20896 46305 20924
rect 45879 20893 45891 20896
rect 45833 20887 45891 20893
rect 46293 20893 46305 20896
rect 46339 20893 46351 20927
rect 46293 20887 46351 20893
rect 29012 20828 35894 20856
rect 28350 20788 28356 20800
rect 26712 20760 28356 20788
rect 28350 20748 28356 20760
rect 28408 20748 28414 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 30837 20791 30895 20797
rect 30837 20788 30849 20791
rect 29052 20760 30849 20788
rect 29052 20748 29058 20760
rect 30837 20757 30849 20760
rect 30883 20757 30895 20791
rect 30837 20751 30895 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 9398 20584 9404 20596
rect 8812 20556 9404 20584
rect 8812 20544 8818 20556
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 11698 20584 11704 20596
rect 11659 20556 11704 20584
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 14734 20584 14740 20596
rect 12406 20556 14740 20584
rect 8205 20519 8263 20525
rect 8205 20485 8217 20519
rect 8251 20516 8263 20519
rect 8941 20519 8999 20525
rect 8941 20516 8953 20519
rect 8251 20488 8953 20516
rect 8251 20485 8263 20488
rect 8205 20479 8263 20485
rect 8941 20485 8953 20488
rect 8987 20485 8999 20519
rect 12406 20516 12434 20556
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 17586 20544 17592 20596
rect 17644 20584 17650 20596
rect 17644 20556 19104 20584
rect 17644 20544 17650 20556
rect 13170 20516 13176 20528
rect 8941 20479 8999 20485
rect 11624 20488 12434 20516
rect 12544 20488 13176 20516
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8294 20448 8300 20460
rect 8159 20420 8300 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 11624 20457 11652 20488
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20417 11667 20451
rect 11609 20411 11667 20417
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20448 12495 20451
rect 12544 20448 12572 20488
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 17770 20516 17776 20528
rect 17328 20488 17776 20516
rect 12483 20420 12572 20448
rect 12621 20451 12679 20457
rect 12483 20417 12495 20420
rect 12437 20411 12495 20417
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 12894 20448 12900 20460
rect 12667 20420 12900 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 12894 20408 12900 20420
rect 12952 20448 12958 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12952 20420 13277 20448
rect 12952 20408 12958 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13722 20448 13728 20460
rect 13495 20420 13728 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 12530 20383 12588 20389
rect 12530 20349 12542 20383
rect 12576 20380 12588 20383
rect 12713 20383 12771 20389
rect 12576 20352 12664 20380
rect 12576 20349 12588 20352
rect 12530 20343 12588 20349
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 9232 20312 9260 20343
rect 12636 20324 12664 20352
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 13464 20380 13492 20411
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16574 20448 16580 20460
rect 15979 20420 16580 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 17328 20457 17356 20488
rect 17770 20476 17776 20488
rect 17828 20476 17834 20528
rect 18414 20476 18420 20528
rect 18472 20516 18478 20528
rect 18472 20488 18552 20516
rect 18472 20476 18478 20488
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20448 17647 20451
rect 17954 20448 17960 20460
rect 17635 20420 17960 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 18322 20448 18328 20460
rect 18283 20420 18328 20448
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 18524 20457 18552 20488
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18230 20380 18236 20392
rect 12759 20352 13492 20380
rect 18191 20352 18236 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 18230 20340 18236 20352
rect 18288 20340 18294 20392
rect 18417 20383 18475 20389
rect 18417 20349 18429 20383
rect 18463 20380 18475 20383
rect 18690 20380 18696 20392
rect 18463 20352 18696 20380
rect 18463 20349 18475 20352
rect 18417 20343 18475 20349
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 4028 20284 9260 20312
rect 4028 20272 4034 20284
rect 12618 20272 12624 20324
rect 12676 20312 12682 20324
rect 13078 20312 13084 20324
rect 12676 20284 13084 20312
rect 12676 20272 12682 20284
rect 13078 20272 13084 20284
rect 13136 20312 13142 20324
rect 14274 20312 14280 20324
rect 13136 20284 14280 20312
rect 13136 20272 13142 20284
rect 14274 20272 14280 20284
rect 14332 20272 14338 20324
rect 17310 20272 17316 20324
rect 17368 20312 17374 20324
rect 17497 20315 17555 20321
rect 17497 20312 17509 20315
rect 17368 20284 17509 20312
rect 17368 20272 17374 20284
rect 17497 20281 17509 20284
rect 17543 20312 17555 20315
rect 18966 20312 18972 20324
rect 17543 20284 18972 20312
rect 17543 20281 17555 20284
rect 17497 20275 17555 20281
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 19076 20312 19104 20556
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20772 20556 20821 20584
rect 20772 20544 20778 20556
rect 20809 20553 20821 20556
rect 20855 20553 20867 20587
rect 20809 20547 20867 20553
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 25501 20587 25559 20593
rect 25501 20584 25513 20587
rect 25188 20556 25513 20584
rect 25188 20544 25194 20556
rect 25501 20553 25513 20556
rect 25547 20553 25559 20587
rect 25501 20547 25559 20553
rect 27525 20587 27583 20593
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 27706 20584 27712 20596
rect 27571 20556 27712 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 27706 20544 27712 20556
rect 27764 20544 27770 20596
rect 29270 20584 29276 20596
rect 29104 20556 29276 20584
rect 20898 20516 20904 20528
rect 20859 20488 20904 20516
rect 20898 20476 20904 20488
rect 20956 20476 20962 20528
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 22428 20488 22753 20516
rect 22428 20476 22434 20488
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 22741 20479 22799 20485
rect 23750 20476 23756 20528
rect 23808 20476 23814 20528
rect 24486 20516 24492 20528
rect 24447 20488 24492 20516
rect 24486 20476 24492 20488
rect 24544 20476 24550 20528
rect 26602 20516 26608 20528
rect 25792 20488 26608 20516
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20448 19763 20451
rect 20717 20451 20775 20457
rect 19751 20420 20668 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20070 20380 20076 20392
rect 20027 20352 20076 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 20438 20380 20444 20392
rect 20399 20352 20444 20380
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 20640 20380 20668 20420
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 20806 20448 20812 20460
rect 20763 20420 20812 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 22462 20448 22468 20460
rect 22423 20420 22468 20448
rect 22462 20408 22468 20420
rect 22520 20408 22526 20460
rect 25792 20457 25820 20488
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 27338 20516 27344 20528
rect 27299 20488 27344 20516
rect 27338 20476 27344 20488
rect 27396 20476 27402 20528
rect 29104 20525 29132 20556
rect 29270 20544 29276 20556
rect 29328 20544 29334 20596
rect 29457 20587 29515 20593
rect 29457 20553 29469 20587
rect 29503 20584 29515 20587
rect 29822 20584 29828 20596
rect 29503 20556 29828 20584
rect 29503 20553 29515 20556
rect 29457 20547 29515 20553
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 45557 20587 45615 20593
rect 45557 20553 45569 20587
rect 45603 20584 45615 20587
rect 45922 20584 45928 20596
rect 45603 20556 45928 20584
rect 45603 20553 45615 20556
rect 45557 20547 45615 20553
rect 45922 20544 45928 20556
rect 45980 20544 45986 20596
rect 29089 20519 29147 20525
rect 29089 20485 29101 20519
rect 29135 20485 29147 20519
rect 29089 20479 29147 20485
rect 42610 20476 42616 20528
rect 42668 20516 42674 20528
rect 42889 20519 42947 20525
rect 42889 20516 42901 20519
rect 42668 20488 42901 20516
rect 42668 20476 42674 20488
rect 42889 20485 42901 20488
rect 42935 20485 42947 20519
rect 42889 20479 42947 20485
rect 43162 20476 43168 20528
rect 43220 20516 43226 20528
rect 43220 20488 47624 20516
rect 43220 20476 43226 20488
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20417 25835 20451
rect 25958 20448 25964 20460
rect 25919 20420 25964 20448
rect 25777 20411 25835 20417
rect 21082 20380 21088 20392
rect 20640 20352 21088 20380
rect 21082 20340 21088 20352
rect 21140 20340 21146 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20349 21235 20383
rect 25700 20380 25728 20411
rect 25958 20408 25964 20420
rect 26016 20408 26022 20460
rect 26050 20408 26056 20460
rect 26108 20448 26114 20460
rect 27157 20451 27215 20457
rect 26108 20420 26153 20448
rect 26108 20408 26114 20420
rect 27157 20417 27169 20451
rect 27203 20448 27215 20451
rect 27982 20448 27988 20460
rect 27203 20420 27988 20448
rect 27203 20417 27215 20420
rect 27157 20411 27215 20417
rect 27982 20408 27988 20420
rect 28040 20408 28046 20460
rect 28905 20451 28963 20457
rect 28905 20417 28917 20451
rect 28951 20448 28963 20451
rect 28994 20448 29000 20460
rect 28951 20420 29000 20448
rect 28951 20417 28963 20420
rect 28905 20411 28963 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29178 20448 29184 20460
rect 29139 20420 29184 20448
rect 29178 20408 29184 20420
rect 29236 20408 29242 20460
rect 29270 20408 29276 20460
rect 29328 20448 29334 20460
rect 45462 20448 45468 20460
rect 29328 20420 29373 20448
rect 45423 20420 45468 20448
rect 29328 20408 29334 20420
rect 45462 20408 45468 20420
rect 45520 20408 45526 20460
rect 46014 20448 46020 20460
rect 45975 20420 46020 20448
rect 46014 20408 46020 20420
rect 46072 20408 46078 20460
rect 47596 20457 47624 20488
rect 47581 20451 47639 20457
rect 47581 20417 47593 20451
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 28074 20380 28080 20392
rect 25700 20352 28080 20380
rect 21177 20343 21235 20349
rect 20088 20312 20116 20340
rect 21192 20312 21220 20343
rect 28074 20340 28080 20352
rect 28132 20380 28138 20392
rect 29454 20380 29460 20392
rect 28132 20352 29460 20380
rect 28132 20340 28138 20352
rect 29454 20340 29460 20352
rect 29512 20340 29518 20392
rect 45738 20340 45744 20392
rect 45796 20380 45802 20392
rect 46293 20383 46351 20389
rect 46293 20380 46305 20383
rect 45796 20352 46305 20380
rect 45796 20340 45802 20352
rect 46293 20349 46305 20352
rect 46339 20349 46351 20383
rect 46293 20343 46351 20349
rect 19076 20284 19932 20312
rect 20088 20284 21220 20312
rect 12066 20204 12072 20256
rect 12124 20244 12130 20256
rect 12253 20247 12311 20253
rect 12253 20244 12265 20247
rect 12124 20216 12265 20244
rect 12124 20204 12130 20216
rect 12253 20213 12265 20216
rect 12299 20213 12311 20247
rect 12253 20207 12311 20213
rect 12342 20204 12348 20256
rect 12400 20244 12406 20256
rect 13357 20247 13415 20253
rect 13357 20244 13369 20247
rect 12400 20216 13369 20244
rect 12400 20204 12406 20216
rect 13357 20213 13369 20216
rect 13403 20213 13415 20247
rect 16022 20244 16028 20256
rect 15983 20216 16028 20244
rect 13357 20207 13415 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 18049 20247 18107 20253
rect 18049 20213 18061 20247
rect 18095 20244 18107 20247
rect 18138 20244 18144 20256
rect 18095 20216 18144 20244
rect 18095 20213 18107 20216
rect 18049 20207 18107 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19904 20253 19932 20284
rect 19521 20247 19579 20253
rect 19521 20244 19533 20247
rect 19484 20216 19533 20244
rect 19484 20204 19490 20216
rect 19521 20213 19533 20216
rect 19567 20213 19579 20247
rect 19521 20207 19579 20213
rect 19889 20247 19947 20253
rect 19889 20213 19901 20247
rect 19935 20244 19947 20247
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 19935 20216 21097 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 21085 20213 21097 20216
rect 21131 20244 21143 20247
rect 21634 20244 21640 20256
rect 21131 20216 21640 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 43162 20244 43168 20256
rect 43123 20216 43168 20244
rect 43162 20204 43168 20216
rect 43220 20204 43226 20256
rect 46474 20204 46480 20256
rect 46532 20244 46538 20256
rect 47673 20247 47731 20253
rect 47673 20244 47685 20247
rect 46532 20216 47685 20244
rect 46532 20204 46538 20216
rect 47673 20213 47685 20216
rect 47719 20213 47731 20247
rect 47673 20207 47731 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 11238 20000 11244 20052
rect 11296 20040 11302 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11296 20012 11897 20040
rect 11296 20000 11302 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 19886 20000 19892 20052
rect 19944 20040 19950 20052
rect 20530 20040 20536 20052
rect 19944 20012 20536 20040
rect 19944 20000 19950 20012
rect 20530 20000 20536 20012
rect 20588 20040 20594 20052
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 20588 20012 20913 20040
rect 20588 20000 20594 20012
rect 20901 20009 20913 20012
rect 20947 20009 20959 20043
rect 21082 20040 21088 20052
rect 21043 20012 21088 20040
rect 20901 20003 20959 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 22002 20040 22008 20052
rect 21963 20012 22008 20040
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22189 20043 22247 20049
rect 22189 20009 22201 20043
rect 22235 20040 22247 20043
rect 22554 20040 22560 20052
rect 22235 20012 22560 20040
rect 22235 20009 22247 20012
rect 22189 20003 22247 20009
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 24857 20043 24915 20049
rect 24857 20009 24869 20043
rect 24903 20040 24915 20043
rect 25222 20040 25228 20052
rect 24903 20012 25228 20040
rect 24903 20009 24915 20012
rect 24857 20003 24915 20009
rect 25222 20000 25228 20012
rect 25280 20000 25286 20052
rect 25685 20043 25743 20049
rect 25685 20009 25697 20043
rect 25731 20040 25743 20043
rect 25958 20040 25964 20052
rect 25731 20012 25964 20040
rect 25731 20009 25743 20012
rect 25685 20003 25743 20009
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 27614 20000 27620 20052
rect 27672 20040 27678 20052
rect 28169 20043 28227 20049
rect 28169 20040 28181 20043
rect 27672 20012 28181 20040
rect 27672 20000 27678 20012
rect 28169 20009 28181 20012
rect 28215 20009 28227 20043
rect 28169 20003 28227 20009
rect 40678 20000 40684 20052
rect 40736 20040 40742 20052
rect 45554 20040 45560 20052
rect 40736 20012 45560 20040
rect 40736 20000 40742 20012
rect 45554 20000 45560 20012
rect 45612 20000 45618 20052
rect 17954 19932 17960 19984
rect 18012 19972 18018 19984
rect 18690 19972 18696 19984
rect 18012 19944 18696 19972
rect 18012 19932 18018 19944
rect 18690 19932 18696 19944
rect 18748 19932 18754 19984
rect 45462 19972 45468 19984
rect 44284 19944 45468 19972
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 9585 19907 9643 19913
rect 9585 19904 9597 19907
rect 9272 19876 9597 19904
rect 9272 19864 9278 19876
rect 9585 19873 9597 19876
rect 9631 19873 9643 19907
rect 9766 19904 9772 19916
rect 9727 19876 9772 19904
rect 9585 19867 9643 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12805 19907 12863 19913
rect 12805 19873 12817 19907
rect 12851 19904 12863 19907
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 12851 19876 14197 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 14185 19867 14243 19873
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1820 19808 2053 19836
rect 1820 19796 1826 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 12066 19836 12072 19848
rect 12027 19808 12072 19836
rect 2041 19799 2099 19805
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 12250 19836 12256 19848
rect 12211 19808 12256 19836
rect 12250 19796 12256 19808
rect 12308 19836 12314 19848
rect 12820 19836 12848 19867
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19904 17739 19907
rect 18414 19904 18420 19916
rect 17727 19876 18420 19904
rect 17727 19873 17739 19876
rect 17681 19867 17739 19873
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 19058 19864 19064 19916
rect 19116 19904 19122 19916
rect 19116 19876 20576 19904
rect 19116 19864 19122 19876
rect 12986 19836 12992 19848
rect 12308 19808 12848 19836
rect 12947 19808 12992 19836
rect 12308 19796 12314 19808
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13262 19796 13268 19848
rect 13320 19836 13326 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13320 19808 14105 19836
rect 13320 19796 13326 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 14093 19799 14151 19805
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 11425 19771 11483 19777
rect 11425 19737 11437 19771
rect 11471 19768 11483 19771
rect 11606 19768 11612 19780
rect 11471 19740 11612 19768
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 12894 19728 12900 19780
rect 12952 19768 12958 19780
rect 14826 19768 14832 19780
rect 12952 19740 14832 19768
rect 12952 19728 12958 19740
rect 14826 19728 14832 19740
rect 14884 19768 14890 19780
rect 15120 19768 15148 19799
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 18233 19839 18291 19845
rect 18233 19836 18245 19839
rect 17276 19808 18245 19836
rect 17276 19796 17282 19808
rect 18233 19805 18245 19808
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 18932 19808 20269 19836
rect 18932 19796 18938 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20548 19836 20576 19876
rect 21726 19864 21732 19916
rect 21784 19904 21790 19916
rect 21784 19876 22094 19904
rect 21784 19864 21790 19876
rect 20898 19836 20904 19848
rect 20548 19808 20904 19836
rect 20257 19799 20315 19805
rect 14884 19740 15148 19768
rect 14884 19728 14890 19740
rect 16850 19728 16856 19780
rect 16908 19768 16914 19780
rect 16945 19771 17003 19777
rect 16945 19768 16957 19771
rect 16908 19740 16957 19768
rect 16908 19728 16914 19740
rect 16945 19737 16957 19740
rect 16991 19737 17003 19771
rect 17862 19768 17868 19780
rect 17823 19740 17868 19768
rect 16945 19731 17003 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 17957 19771 18015 19777
rect 17957 19737 17969 19771
rect 18003 19768 18015 19771
rect 18322 19768 18328 19780
rect 18003 19740 18328 19768
rect 18003 19737 18015 19740
rect 17957 19731 18015 19737
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19058 19728 19064 19780
rect 19116 19768 19122 19780
rect 19705 19771 19763 19777
rect 19705 19768 19717 19771
rect 19116 19740 19717 19768
rect 19116 19728 19122 19740
rect 19705 19737 19717 19740
rect 19751 19737 19763 19771
rect 19886 19768 19892 19780
rect 19847 19740 19892 19768
rect 19705 19731 19763 19737
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 20732 19777 20760 19808
rect 20898 19796 20904 19808
rect 20956 19836 20962 19848
rect 20956 19808 21956 19836
rect 22066 19811 22094 19876
rect 24394 19864 24400 19916
rect 24452 19904 24458 19916
rect 24489 19907 24547 19913
rect 24489 19904 24501 19907
rect 24452 19876 24501 19904
rect 24452 19864 24458 19876
rect 24489 19873 24501 19876
rect 24535 19904 24547 19907
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 24535 19876 25329 19904
rect 24535 19873 24547 19876
rect 24489 19867 24547 19873
rect 25317 19873 25329 19876
rect 25363 19904 25375 19907
rect 27801 19907 27859 19913
rect 27801 19904 27813 19907
rect 25363 19876 27813 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 27801 19873 27813 19876
rect 27847 19904 27859 19907
rect 29178 19904 29184 19916
rect 27847 19876 29184 19904
rect 27847 19873 27859 19876
rect 27801 19867 27859 19873
rect 29178 19864 29184 19876
rect 29236 19904 29242 19916
rect 30193 19907 30251 19913
rect 30193 19904 30205 19907
rect 29236 19876 30205 19904
rect 29236 19864 29242 19876
rect 30193 19873 30205 19876
rect 30239 19873 30251 19907
rect 30193 19867 30251 19873
rect 24670 19836 24676 19848
rect 20956 19796 20962 19808
rect 19981 19771 20039 19777
rect 19981 19737 19993 19771
rect 20027 19768 20039 19771
rect 20717 19771 20775 19777
rect 20027 19740 20668 19768
rect 20027 19737 20039 19740
rect 19981 19731 20039 19737
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 13173 19703 13231 19709
rect 13173 19700 13185 19703
rect 12860 19672 13185 19700
rect 12860 19660 12866 19672
rect 13173 19669 13185 19672
rect 13219 19669 13231 19703
rect 13173 19663 13231 19669
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 18230 19700 18236 19712
rect 18095 19672 18236 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 18230 19660 18236 19672
rect 18288 19700 18294 19712
rect 18874 19700 18880 19712
rect 18288 19672 18880 19700
rect 18288 19660 18294 19672
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 20070 19700 20076 19712
rect 20031 19672 20076 19700
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20640 19700 20668 19740
rect 20717 19737 20729 19771
rect 20763 19737 20775 19771
rect 20717 19731 20775 19737
rect 20806 19728 20812 19780
rect 20864 19768 20870 19780
rect 21821 19771 21879 19777
rect 21821 19768 21833 19771
rect 20864 19740 21833 19768
rect 20864 19728 20870 19740
rect 21821 19737 21833 19740
rect 21867 19737 21879 19771
rect 21821 19731 21879 19737
rect 20898 19700 20904 19712
rect 20956 19709 20962 19712
rect 20956 19703 20975 19709
rect 20640 19672 20904 19700
rect 20898 19660 20904 19672
rect 20963 19669 20975 19703
rect 21928 19700 21956 19808
rect 22051 19805 22109 19811
rect 24631 19808 24676 19836
rect 22051 19771 22063 19805
rect 22097 19771 22109 19805
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19805 25559 19839
rect 25501 19799 25559 19805
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19836 28043 19839
rect 28442 19836 28448 19848
rect 28031 19808 28448 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 22051 19765 22109 19771
rect 25130 19728 25136 19780
rect 25188 19768 25194 19780
rect 25516 19768 25544 19799
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 30006 19836 30012 19848
rect 29967 19808 30012 19836
rect 30006 19796 30012 19808
rect 30064 19796 30070 19848
rect 44284 19845 44312 19944
rect 45462 19932 45468 19944
rect 45520 19932 45526 19984
rect 46106 19932 46112 19984
rect 46164 19972 46170 19984
rect 46164 19944 46980 19972
rect 46164 19932 46170 19944
rect 45833 19907 45891 19913
rect 45833 19904 45845 19907
rect 44468 19876 45845 19904
rect 44468 19845 44496 19876
rect 45833 19873 45845 19876
rect 45879 19873 45891 19907
rect 46474 19904 46480 19916
rect 46435 19876 46480 19904
rect 45833 19867 45891 19873
rect 46474 19864 46480 19876
rect 46532 19864 46538 19916
rect 46952 19913 46980 19944
rect 46937 19907 46995 19913
rect 46937 19873 46949 19907
rect 46983 19873 46995 19907
rect 46937 19867 46995 19873
rect 44269 19839 44327 19845
rect 44269 19805 44281 19839
rect 44315 19805 44327 19839
rect 44269 19799 44327 19805
rect 44453 19839 44511 19845
rect 44453 19805 44465 19839
rect 44499 19805 44511 19839
rect 44453 19799 44511 19805
rect 45465 19839 45523 19845
rect 45465 19805 45477 19839
rect 45511 19805 45523 19839
rect 45465 19799 45523 19805
rect 25188 19740 25544 19768
rect 45480 19768 45508 19799
rect 45554 19796 45560 19848
rect 45612 19836 45618 19848
rect 45649 19839 45707 19845
rect 45649 19836 45661 19839
rect 45612 19808 45661 19836
rect 45612 19796 45618 19808
rect 45649 19805 45661 19808
rect 45695 19805 45707 19839
rect 45649 19799 45707 19805
rect 46198 19796 46204 19848
rect 46256 19836 46262 19848
rect 46293 19839 46351 19845
rect 46293 19836 46305 19839
rect 46256 19808 46305 19836
rect 46256 19796 46262 19808
rect 46293 19805 46305 19808
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 45922 19768 45928 19780
rect 45480 19740 45928 19768
rect 25188 19728 25194 19740
rect 45922 19728 45928 19740
rect 45980 19768 45986 19780
rect 47302 19768 47308 19780
rect 45980 19740 47308 19768
rect 45980 19728 45986 19740
rect 47302 19728 47308 19740
rect 47360 19728 47366 19780
rect 22462 19700 22468 19712
rect 21928 19672 22468 19700
rect 20956 19663 20975 19669
rect 20956 19660 20962 19663
rect 22462 19660 22468 19672
rect 22520 19660 22526 19712
rect 44361 19703 44419 19709
rect 44361 19669 44373 19703
rect 44407 19700 44419 19703
rect 46106 19700 46112 19712
rect 44407 19672 46112 19700
rect 44407 19669 44419 19672
rect 44361 19663 44419 19669
rect 46106 19660 46112 19672
rect 46164 19660 46170 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12986 19496 12992 19508
rect 12483 19468 12992 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12986 19456 12992 19468
rect 13044 19456 13050 19508
rect 14090 19496 14096 19508
rect 13188 19468 14096 19496
rect 9398 19428 9404 19440
rect 9359 19400 9404 19428
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 12069 19431 12127 19437
rect 12069 19397 12081 19431
rect 12115 19428 12127 19431
rect 13078 19428 13084 19440
rect 12115 19400 13084 19428
rect 12115 19397 12127 19400
rect 12069 19391 12127 19397
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 9582 19360 9588 19372
rect 9355 19332 9588 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 12253 19363 12311 19369
rect 12253 19329 12265 19363
rect 12299 19360 12311 19363
rect 12618 19360 12624 19372
rect 12299 19332 12624 19360
rect 12299 19329 12333 19332
rect 12253 19323 12333 19329
rect 12268 19306 12333 19323
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13188 19369 13216 19468
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16080 19468 17172 19496
rect 16080 19456 16086 19468
rect 14918 19428 14924 19440
rect 14674 19400 14924 19428
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 17034 19428 17040 19440
rect 16991 19400 17040 19428
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 17144 19428 17172 19468
rect 17770 19456 17776 19508
rect 17828 19496 17834 19508
rect 18230 19496 18236 19508
rect 17828 19468 18236 19496
rect 17828 19456 17834 19468
rect 18230 19456 18236 19468
rect 18288 19496 18294 19508
rect 18417 19499 18475 19505
rect 18417 19496 18429 19499
rect 18288 19468 18429 19496
rect 18288 19456 18294 19468
rect 18417 19465 18429 19468
rect 18463 19465 18475 19499
rect 18966 19496 18972 19508
rect 18927 19468 18972 19496
rect 18417 19459 18475 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 45281 19499 45339 19505
rect 45281 19465 45293 19499
rect 45327 19496 45339 19499
rect 45462 19496 45468 19508
rect 45327 19468 45468 19496
rect 45327 19465 45339 19468
rect 45281 19459 45339 19465
rect 45462 19456 45468 19468
rect 45520 19456 45526 19508
rect 45922 19456 45928 19508
rect 45980 19456 45986 19508
rect 40678 19428 40684 19440
rect 17144 19400 17434 19428
rect 35866 19400 40684 19428
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 15562 19360 15568 19372
rect 14884 19332 14964 19360
rect 15523 19332 15568 19360
rect 14884 19320 14890 19332
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 12268 19292 12296 19306
rect 13446 19292 13452 19304
rect 9272 19264 12296 19292
rect 12406 19264 13124 19292
rect 13407 19264 13452 19292
rect 9272 19252 9278 19264
rect 3878 19184 3884 19236
rect 3936 19224 3942 19236
rect 12406 19224 12434 19264
rect 3936 19196 12434 19224
rect 3936 19184 3942 19196
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 12986 19156 12992 19168
rect 3476 19128 12992 19156
rect 3476 19116 3482 19128
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 13096 19156 13124 19264
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 14936 19301 14964 19332
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 18874 19360 18880 19372
rect 18835 19332 18880 19360
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19334 19360 19340 19372
rect 19107 19332 19340 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 22462 19360 22468 19372
rect 22423 19332 22468 19360
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 24578 19360 24584 19372
rect 24351 19332 24584 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 24578 19320 24584 19332
rect 24636 19320 24642 19372
rect 27525 19363 27583 19369
rect 27525 19329 27537 19363
rect 27571 19360 27583 19363
rect 35866 19360 35894 19400
rect 40678 19388 40684 19400
rect 40736 19388 40742 19440
rect 45554 19428 45560 19440
rect 45204 19400 45560 19428
rect 27571 19332 35894 19360
rect 42429 19363 42487 19369
rect 27571 19329 27583 19332
rect 27525 19323 27583 19329
rect 42429 19329 42441 19363
rect 42475 19360 42487 19363
rect 43162 19360 43168 19372
rect 42475 19332 43168 19360
rect 42475 19329 42487 19332
rect 42429 19323 42487 19329
rect 43162 19320 43168 19332
rect 43220 19360 43226 19372
rect 43898 19360 43904 19372
rect 43220 19332 43904 19360
rect 43220 19320 43226 19332
rect 43898 19320 43904 19332
rect 43956 19320 43962 19372
rect 45204 19369 45232 19400
rect 45554 19388 45560 19400
rect 45612 19388 45618 19440
rect 45940 19428 45968 19456
rect 45664 19400 45968 19428
rect 45189 19363 45247 19369
rect 45189 19329 45201 19363
rect 45235 19329 45247 19363
rect 45189 19323 45247 19329
rect 45373 19363 45431 19369
rect 45373 19329 45385 19363
rect 45419 19360 45431 19363
rect 45664 19360 45692 19400
rect 45419 19332 45692 19360
rect 45419 19329 45431 19332
rect 45373 19323 45431 19329
rect 45738 19320 45744 19372
rect 45796 19360 45802 19372
rect 45925 19363 45983 19369
rect 45925 19360 45937 19363
rect 45796 19332 45937 19360
rect 45796 19320 45802 19332
rect 45925 19329 45937 19332
rect 45971 19329 45983 19363
rect 46106 19360 46112 19372
rect 46067 19332 46112 19360
rect 45925 19323 45983 19329
rect 46106 19320 46112 19332
rect 46164 19320 46170 19372
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15841 19295 15899 19301
rect 15841 19261 15853 19295
rect 15887 19292 15899 19295
rect 16669 19295 16727 19301
rect 16669 19292 16681 19295
rect 15887 19264 16681 19292
rect 15887 19261 15899 19264
rect 15841 19255 15899 19261
rect 16669 19261 16681 19264
rect 16715 19261 16727 19295
rect 22370 19292 22376 19304
rect 16669 19255 16727 19261
rect 16776 19264 22376 19292
rect 16776 19224 16804 19264
rect 22370 19252 22376 19264
rect 22428 19252 22434 19304
rect 22554 19292 22560 19304
rect 22515 19264 22560 19292
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 46198 19252 46204 19304
rect 46256 19292 46262 19304
rect 46845 19295 46903 19301
rect 46845 19292 46857 19295
rect 46256 19264 46857 19292
rect 46256 19252 46262 19264
rect 46845 19261 46857 19264
rect 46891 19261 46903 19295
rect 46845 19255 46903 19261
rect 14476 19196 16804 19224
rect 14476 19156 14504 19196
rect 17954 19184 17960 19236
rect 18012 19224 18018 19236
rect 18012 19196 19104 19224
rect 18012 19184 18018 19196
rect 13096 19128 14504 19156
rect 17494 19116 17500 19168
rect 17552 19156 17558 19168
rect 18138 19156 18144 19168
rect 17552 19128 18144 19156
rect 17552 19116 17558 19128
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 19076 19156 19104 19196
rect 22066 19196 35894 19224
rect 22066 19156 22094 19196
rect 19076 19128 22094 19156
rect 22833 19159 22891 19165
rect 22833 19125 22845 19159
rect 22879 19156 22891 19159
rect 23014 19156 23020 19168
rect 22879 19128 23020 19156
rect 22879 19125 22891 19128
rect 22833 19119 22891 19125
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 24489 19159 24547 19165
rect 24489 19156 24501 19159
rect 24452 19128 24501 19156
rect 24452 19116 24458 19128
rect 24489 19125 24501 19128
rect 24535 19125 24547 19159
rect 27614 19156 27620 19168
rect 27575 19128 27620 19156
rect 24489 19119 24547 19125
rect 27614 19116 27620 19128
rect 27672 19116 27678 19168
rect 35866 19156 35894 19196
rect 41322 19156 41328 19168
rect 35866 19128 41328 19156
rect 41322 19116 41328 19128
rect 41380 19116 41386 19168
rect 41414 19116 41420 19168
rect 41472 19156 41478 19168
rect 42521 19159 42579 19165
rect 42521 19156 42533 19159
rect 41472 19128 42533 19156
rect 41472 19116 41478 19128
rect 42521 19125 42533 19128
rect 42567 19125 42579 19159
rect 47762 19156 47768 19168
rect 47723 19128 47768 19156
rect 42521 19119 42579 19125
rect 47762 19116 47768 19128
rect 47820 19116 47826 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1946 18912 1952 18964
rect 2004 18952 2010 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2004 18924 2237 18952
rect 2004 18912 2010 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 2314 18912 2320 18964
rect 2372 18952 2378 18964
rect 12621 18955 12679 18961
rect 2372 18924 12434 18952
rect 2372 18912 2378 18924
rect 4798 18844 4804 18896
rect 4856 18884 4862 18896
rect 4856 18856 9720 18884
rect 4856 18844 4862 18856
rect 9214 18816 9220 18828
rect 9175 18788 9220 18816
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 9398 18816 9404 18828
rect 9359 18788 9404 18816
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9692 18825 9720 18856
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18785 9735 18819
rect 12250 18816 12256 18828
rect 12211 18788 12256 18816
rect 9677 18779 9735 18785
rect 12250 18776 12256 18788
rect 12308 18776 12314 18828
rect 12406 18816 12434 18924
rect 12621 18921 12633 18955
rect 12667 18952 12679 18955
rect 13446 18952 13452 18964
rect 12667 18924 13452 18952
rect 12667 18921 12679 18924
rect 12621 18915 12679 18921
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 14918 18952 14924 18964
rect 14879 18924 14924 18952
rect 14918 18912 14924 18924
rect 14976 18912 14982 18964
rect 17954 18952 17960 18964
rect 15028 18924 17960 18952
rect 12986 18844 12992 18896
rect 13044 18884 13050 18896
rect 15028 18884 15056 18924
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18322 18952 18328 18964
rect 18283 18924 18328 18952
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18506 18952 18512 18964
rect 18467 18924 18512 18952
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 19978 18952 19984 18964
rect 19939 18924 19984 18952
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 20717 18955 20775 18961
rect 20717 18952 20729 18955
rect 20312 18924 20729 18952
rect 20312 18912 20318 18924
rect 20717 18921 20729 18924
rect 20763 18921 20775 18955
rect 20898 18952 20904 18964
rect 20859 18924 20904 18952
rect 20717 18915 20775 18921
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 32490 18952 32496 18964
rect 22066 18924 32496 18952
rect 17494 18884 17500 18896
rect 13044 18856 15056 18884
rect 17455 18856 17500 18884
rect 13044 18844 13050 18856
rect 17494 18844 17500 18856
rect 17552 18844 17558 18896
rect 22066 18884 22094 18924
rect 32490 18912 32496 18924
rect 32548 18912 32554 18964
rect 45649 18955 45707 18961
rect 45649 18921 45661 18955
rect 45695 18952 45707 18955
rect 46014 18952 46020 18964
rect 45695 18924 46020 18952
rect 45695 18921 45707 18924
rect 45649 18915 45707 18921
rect 46014 18912 46020 18924
rect 46072 18912 46078 18964
rect 17604 18856 22094 18884
rect 17604 18816 17632 18856
rect 22370 18844 22376 18896
rect 22428 18884 22434 18896
rect 28166 18884 28172 18896
rect 22428 18856 28172 18884
rect 22428 18844 22434 18856
rect 28166 18844 28172 18856
rect 28224 18844 28230 18896
rect 28445 18887 28503 18893
rect 28445 18853 28457 18887
rect 28491 18884 28503 18887
rect 28491 18856 35894 18884
rect 28491 18853 28503 18856
rect 28445 18847 28503 18853
rect 12406 18788 17632 18816
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18785 17739 18819
rect 26145 18819 26203 18825
rect 26145 18816 26157 18819
rect 17681 18779 17739 18785
rect 22066 18788 26157 18816
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 6546 18748 6552 18760
rect 2188 18720 6552 18748
rect 2188 18708 2194 18720
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 11701 18751 11759 18757
rect 10612 18720 11652 18748
rect 2038 18640 2044 18692
rect 2096 18680 2102 18692
rect 10612 18680 10640 18720
rect 2096 18652 10640 18680
rect 2096 18640 2102 18652
rect 11514 18612 11520 18624
rect 11475 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 11624 18612 11652 18720
rect 11701 18717 11713 18751
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12894 18748 12900 18760
rect 12391 18720 12900 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 11716 18680 11744 18711
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13403 18720 14289 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 14277 18717 14289 18720
rect 14323 18748 14335 18751
rect 14458 18748 14464 18760
rect 14323 18720 14464 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 16761 18751 16819 18757
rect 14884 18720 14929 18748
rect 14884 18708 14890 18720
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 17696 18748 17724 18779
rect 22066 18748 22094 18788
rect 26145 18785 26157 18788
rect 26191 18785 26203 18819
rect 26145 18779 26203 18785
rect 26510 18776 26516 18828
rect 26568 18816 26574 18828
rect 27522 18816 27528 18828
rect 26568 18788 27528 18816
rect 26568 18776 26574 18788
rect 27522 18776 27528 18788
rect 27580 18776 27586 18828
rect 16807 18720 17724 18748
rect 17788 18720 22094 18748
rect 22373 18751 22431 18757
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 12802 18680 12808 18692
rect 11716 18652 12808 18680
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 17218 18680 17224 18692
rect 13188 18652 13492 18680
rect 13188 18612 13216 18652
rect 13354 18612 13360 18624
rect 11624 18584 13216 18612
rect 13315 18584 13360 18612
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 13464 18612 13492 18652
rect 16500 18652 17080 18680
rect 17179 18652 17224 18680
rect 16500 18612 16528 18652
rect 13464 18584 16528 18612
rect 16577 18615 16635 18621
rect 16577 18581 16589 18615
rect 16623 18612 16635 18615
rect 16942 18612 16948 18624
rect 16623 18584 16948 18612
rect 16623 18581 16635 18584
rect 16577 18575 16635 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17052 18612 17080 18652
rect 17218 18640 17224 18652
rect 17276 18640 17282 18692
rect 17788 18612 17816 18720
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 24394 18748 24400 18760
rect 24355 18720 24400 18748
rect 22373 18711 22431 18717
rect 18138 18680 18144 18692
rect 18099 18652 18144 18680
rect 18138 18640 18144 18652
rect 18196 18640 18202 18692
rect 19705 18683 19763 18689
rect 19705 18680 19717 18683
rect 18248 18652 19717 18680
rect 17052 18584 17816 18612
rect 18046 18572 18052 18624
rect 18104 18612 18110 18624
rect 18248 18612 18276 18652
rect 19705 18649 19717 18652
rect 19751 18649 19763 18683
rect 19705 18643 19763 18649
rect 20533 18683 20591 18689
rect 20533 18649 20545 18683
rect 20579 18680 20591 18683
rect 20622 18680 20628 18692
rect 20579 18652 20628 18680
rect 20579 18649 20591 18652
rect 20533 18643 20591 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 20714 18640 20720 18692
rect 20772 18689 20778 18692
rect 20772 18683 20791 18689
rect 20779 18649 20791 18683
rect 20772 18643 20791 18649
rect 20772 18640 20778 18643
rect 18104 18584 18276 18612
rect 18351 18615 18409 18621
rect 18104 18572 18110 18584
rect 18351 18581 18363 18615
rect 18397 18612 18409 18615
rect 18690 18612 18696 18624
rect 18397 18584 18696 18612
rect 18397 18581 18409 18584
rect 18351 18575 18409 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19978 18572 19984 18624
rect 20036 18612 20042 18624
rect 20990 18612 20996 18624
rect 20036 18584 20996 18612
rect 20036 18572 20042 18584
rect 20990 18572 20996 18584
rect 21048 18612 21054 18624
rect 22388 18612 22416 18711
rect 24394 18708 24400 18720
rect 24452 18708 24458 18760
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18717 26019 18751
rect 28258 18748 28264 18760
rect 28219 18720 28264 18748
rect 25961 18711 26019 18717
rect 25976 18680 26004 18711
rect 28258 18708 28264 18720
rect 28316 18708 28322 18760
rect 35866 18748 35894 18856
rect 41322 18844 41328 18896
rect 41380 18884 41386 18896
rect 41380 18856 41736 18884
rect 41380 18844 41386 18856
rect 41414 18816 41420 18828
rect 41375 18788 41420 18816
rect 41414 18776 41420 18788
rect 41472 18776 41478 18828
rect 41708 18825 41736 18856
rect 41693 18819 41751 18825
rect 41693 18785 41705 18819
rect 41739 18785 41751 18819
rect 41693 18779 41751 18785
rect 45830 18776 45836 18828
rect 45888 18816 45894 18828
rect 46014 18816 46020 18828
rect 45888 18788 46020 18816
rect 45888 18776 45894 18788
rect 46014 18776 46020 18788
rect 46072 18776 46078 18828
rect 46293 18819 46351 18825
rect 46293 18785 46305 18819
rect 46339 18816 46351 18819
rect 47762 18816 47768 18828
rect 46339 18788 47768 18816
rect 46339 18785 46351 18788
rect 46293 18779 46351 18785
rect 47762 18776 47768 18788
rect 47820 18776 47826 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 41230 18748 41236 18760
rect 35866 18720 41236 18748
rect 41230 18708 41236 18720
rect 41288 18708 41294 18760
rect 45554 18708 45560 18760
rect 45612 18748 45618 18760
rect 45741 18751 45799 18757
rect 45612 18720 45657 18748
rect 45612 18708 45618 18720
rect 45741 18717 45753 18751
rect 45787 18748 45799 18751
rect 45922 18748 45928 18760
rect 45787 18720 45928 18748
rect 45787 18717 45799 18720
rect 45741 18711 45799 18717
rect 45922 18708 45928 18720
rect 45980 18708 45986 18760
rect 27706 18680 27712 18692
rect 25976 18652 27712 18680
rect 27706 18640 27712 18652
rect 27764 18640 27770 18692
rect 29641 18683 29699 18689
rect 29641 18680 29653 18683
rect 27816 18652 29653 18680
rect 21048 18584 22416 18612
rect 22557 18615 22615 18621
rect 21048 18572 21054 18584
rect 22557 18581 22569 18615
rect 22603 18612 22615 18615
rect 22738 18612 22744 18624
rect 22603 18584 22744 18612
rect 22603 18581 22615 18584
rect 22557 18575 22615 18581
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 24486 18612 24492 18624
rect 24447 18584 24492 18612
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 27816 18612 27844 18652
rect 29641 18649 29653 18652
rect 29687 18649 29699 18683
rect 29641 18643 29699 18649
rect 29733 18683 29791 18689
rect 29733 18649 29745 18683
rect 29779 18649 29791 18683
rect 30650 18680 30656 18692
rect 30611 18652 30656 18680
rect 29733 18643 29791 18649
rect 24820 18584 27844 18612
rect 24820 18572 24826 18584
rect 29086 18572 29092 18624
rect 29144 18612 29150 18624
rect 29748 18612 29776 18643
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 47670 18680 47676 18692
rect 46523 18652 47676 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 47670 18640 47676 18652
rect 47728 18640 47734 18692
rect 29144 18584 29776 18612
rect 29144 18572 29150 18584
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 2314 18408 2320 18420
rect 1627 18380 2320 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 2314 18368 2320 18380
rect 2372 18368 2378 18420
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 25682 18408 25688 18420
rect 5040 18380 25688 18408
rect 5040 18368 5046 18380
rect 25682 18368 25688 18380
rect 25740 18408 25746 18420
rect 30650 18408 30656 18420
rect 25740 18380 26280 18408
rect 25740 18368 25746 18380
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 12897 18343 12955 18349
rect 12897 18340 12909 18343
rect 11572 18312 12909 18340
rect 11572 18300 11578 18312
rect 12897 18309 12909 18312
rect 12943 18309 12955 18343
rect 14182 18340 14188 18352
rect 14122 18312 14188 18340
rect 12897 18303 12955 18309
rect 14182 18300 14188 18312
rect 14240 18300 14246 18352
rect 16942 18340 16948 18352
rect 16903 18312 16948 18340
rect 16942 18300 16948 18312
rect 17000 18300 17006 18352
rect 17954 18300 17960 18352
rect 18012 18300 18018 18352
rect 20530 18340 20536 18352
rect 19536 18312 20536 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 14458 18232 14464 18284
rect 14516 18272 14522 18284
rect 15562 18272 15568 18284
rect 14516 18244 15568 18272
rect 14516 18232 14522 18244
rect 15562 18232 15568 18244
rect 15620 18272 15626 18284
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15620 18244 15669 18272
rect 15620 18232 15626 18244
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 19334 18272 19340 18284
rect 19295 18244 19340 18272
rect 15657 18235 15715 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 19536 18281 19564 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 23014 18340 23020 18352
rect 22975 18312 23020 18340
rect 23014 18300 23020 18312
rect 23072 18300 23078 18352
rect 24486 18340 24492 18352
rect 24242 18312 24492 18340
rect 24486 18300 24492 18312
rect 24544 18300 24550 18352
rect 26252 18349 26280 18380
rect 27356 18380 30656 18408
rect 26237 18343 26295 18349
rect 26237 18309 26249 18343
rect 26283 18309 26295 18343
rect 27356 18340 27384 18380
rect 30650 18368 30656 18380
rect 30708 18408 30714 18420
rect 40218 18408 40224 18420
rect 30708 18380 40224 18408
rect 30708 18368 30714 18380
rect 40218 18368 40224 18380
rect 40276 18368 40282 18420
rect 47670 18408 47676 18420
rect 47631 18380 47676 18408
rect 47670 18368 47676 18380
rect 47728 18368 47734 18420
rect 26237 18303 26295 18309
rect 27264 18312 27384 18340
rect 27433 18343 27491 18349
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19484 18244 19533 18272
rect 19484 18232 19490 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19978 18232 19984 18284
rect 20036 18272 20042 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20036 18244 20177 18272
rect 20036 18232 20042 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20990 18272 20996 18284
rect 20951 18244 20996 18272
rect 20165 18235 20223 18241
rect 20990 18232 20996 18244
rect 21048 18232 21054 18284
rect 21818 18272 21824 18284
rect 21731 18244 21824 18272
rect 21818 18232 21824 18244
rect 21876 18272 21882 18284
rect 22738 18272 22744 18284
rect 21876 18244 22600 18272
rect 22699 18244 22744 18272
rect 21876 18232 21882 18244
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 13354 18204 13360 18216
rect 12667 18176 13360 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 14274 18164 14280 18216
rect 14332 18204 14338 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14332 18176 14381 18204
rect 14332 18164 14338 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 15933 18207 15991 18213
rect 15933 18173 15945 18207
rect 15979 18204 15991 18207
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 15979 18176 16681 18204
rect 15979 18173 15991 18176
rect 15933 18167 15991 18173
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18204 20315 18207
rect 20438 18204 20444 18216
rect 20303 18176 20444 18204
rect 20303 18173 20315 18176
rect 20257 18167 20315 18173
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 22572 18204 22600 18244
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 25498 18232 25504 18284
rect 25556 18272 25562 18284
rect 26053 18275 26111 18281
rect 26053 18272 26065 18275
rect 25556 18244 26065 18272
rect 25556 18232 25562 18244
rect 26053 18241 26065 18244
rect 26099 18272 26111 18275
rect 27264 18272 27292 18312
rect 27433 18309 27445 18343
rect 27479 18340 27491 18343
rect 27614 18340 27620 18352
rect 27479 18312 27620 18340
rect 27479 18309 27491 18312
rect 27433 18303 27491 18309
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 46382 18272 46388 18284
rect 26099 18244 27292 18272
rect 46343 18244 46388 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 46382 18232 46388 18244
rect 46440 18232 46446 18284
rect 47118 18232 47124 18284
rect 47176 18272 47182 18284
rect 47486 18272 47492 18284
rect 47176 18244 47492 18272
rect 47176 18232 47182 18244
rect 47486 18232 47492 18244
rect 47544 18272 47550 18284
rect 47581 18275 47639 18281
rect 47581 18272 47593 18275
rect 47544 18244 47593 18272
rect 47544 18232 47550 18244
rect 47581 18241 47593 18244
rect 47627 18241 47639 18275
rect 47581 18235 47639 18241
rect 24394 18204 24400 18216
rect 22572 18176 24400 18204
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 24765 18207 24823 18213
rect 24765 18173 24777 18207
rect 24811 18173 24823 18207
rect 24765 18167 24823 18173
rect 27249 18207 27307 18213
rect 27249 18173 27261 18207
rect 27295 18204 27307 18207
rect 28074 18204 28080 18216
rect 27295 18176 28080 18204
rect 27295 18173 27307 18176
rect 27249 18167 27307 18173
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 18380 18040 18429 18068
rect 18380 18028 18386 18040
rect 18417 18037 18429 18040
rect 18463 18068 18475 18071
rect 18506 18068 18512 18080
rect 18463 18040 18512 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19426 18068 19432 18080
rect 19383 18040 19432 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 20533 18071 20591 18077
rect 20533 18037 20545 18071
rect 20579 18068 20591 18071
rect 20806 18068 20812 18080
rect 20579 18040 20812 18068
rect 20579 18037 20591 18040
rect 20533 18031 20591 18037
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21910 18068 21916 18080
rect 21871 18040 21916 18068
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 24780 18068 24808 18167
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 28166 18164 28172 18216
rect 28224 18204 28230 18216
rect 28224 18176 28269 18204
rect 28224 18164 28230 18176
rect 22520 18040 24808 18068
rect 26421 18071 26479 18077
rect 22520 18028 22526 18040
rect 26421 18037 26433 18071
rect 26467 18068 26479 18071
rect 27154 18068 27160 18080
rect 26467 18040 27160 18068
rect 26467 18037 26479 18040
rect 26421 18031 26479 18037
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 46201 18071 46259 18077
rect 46201 18037 46213 18071
rect 46247 18068 46259 18071
rect 46842 18068 46848 18080
rect 46247 18040 46848 18068
rect 46247 18037 46259 18040
rect 46201 18031 46259 18037
rect 46842 18028 46848 18040
rect 46900 18028 46906 18080
rect 47026 18068 47032 18080
rect 46987 18040 47032 18068
rect 47026 18028 47032 18040
rect 47084 18028 47090 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 14182 17864 14188 17876
rect 14143 17836 14188 17864
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 16945 17867 17003 17873
rect 16945 17833 16957 17867
rect 16991 17864 17003 17867
rect 17954 17864 17960 17876
rect 16991 17836 17960 17864
rect 16991 17833 17003 17836
rect 16945 17827 17003 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 19392 17836 19809 17864
rect 19392 17824 19398 17836
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 20990 17864 20996 17876
rect 19797 17827 19855 17833
rect 20548 17836 20996 17864
rect 20548 17737 20576 17836
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 46658 17796 46664 17808
rect 39960 17768 46664 17796
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17697 20591 17731
rect 20806 17728 20812 17740
rect 20767 17700 20812 17728
rect 20533 17691 20591 17697
rect 20806 17688 20812 17700
rect 20864 17688 20870 17740
rect 39960 17737 39988 17768
rect 46658 17756 46664 17768
rect 46716 17756 46722 17808
rect 39945 17731 40003 17737
rect 39945 17697 39957 17731
rect 39991 17697 40003 17731
rect 40218 17728 40224 17740
rect 40179 17700 40224 17728
rect 39945 17691 40003 17697
rect 40218 17688 40224 17700
rect 40276 17688 40282 17740
rect 46477 17731 46535 17737
rect 46477 17697 46489 17731
rect 46523 17728 46535 17731
rect 48038 17728 48044 17740
rect 46523 17700 48044 17728
rect 46523 17697 46535 17700
rect 46477 17691 46535 17697
rect 48038 17688 48044 17700
rect 48096 17688 48102 17740
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14826 17660 14832 17672
rect 14139 17632 14832 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16632 17632 16865 17660
rect 16632 17620 16638 17632
rect 16853 17629 16865 17632
rect 16899 17660 16911 17663
rect 17678 17660 17684 17672
rect 16899 17632 17684 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18104 17632 18245 17660
rect 18104 17620 18110 17632
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20438 17660 20444 17672
rect 20119 17632 20444 17660
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 21910 17620 21916 17672
rect 21968 17620 21974 17672
rect 25498 17660 25504 17672
rect 25459 17632 25504 17660
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 25682 17660 25688 17672
rect 25643 17632 25688 17660
rect 25682 17620 25688 17632
rect 25740 17620 25746 17672
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17660 25927 17663
rect 26418 17660 26424 17672
rect 25915 17632 26424 17660
rect 25915 17629 25927 17632
rect 25869 17623 25927 17629
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 27062 17660 27068 17672
rect 27023 17632 27068 17660
rect 27062 17620 27068 17632
rect 27120 17620 27126 17672
rect 45462 17620 45468 17672
rect 45520 17660 45526 17672
rect 46293 17663 46351 17669
rect 46293 17660 46305 17663
rect 45520 17632 46305 17660
rect 45520 17620 45526 17632
rect 46293 17629 46305 17632
rect 46339 17629 46351 17663
rect 46293 17623 46351 17629
rect 47854 17620 47860 17672
rect 47912 17660 47918 17672
rect 48133 17663 48191 17669
rect 48133 17660 48145 17663
rect 47912 17632 48145 17660
rect 47912 17620 47918 17632
rect 48056 17604 48084 17632
rect 48133 17629 48145 17632
rect 48179 17629 48191 17663
rect 48133 17623 48191 17629
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19797 17595 19855 17601
rect 19797 17592 19809 17595
rect 19392 17564 19809 17592
rect 19392 17552 19398 17564
rect 19797 17561 19809 17564
rect 19843 17561 19855 17595
rect 28074 17592 28080 17604
rect 27922 17564 28080 17592
rect 19797 17555 19855 17561
rect 28074 17552 28080 17564
rect 28132 17552 28138 17604
rect 40037 17595 40095 17601
rect 40037 17561 40049 17595
rect 40083 17592 40095 17595
rect 40402 17592 40408 17604
rect 40083 17564 40408 17592
rect 40083 17561 40095 17564
rect 40037 17555 40095 17561
rect 40402 17552 40408 17564
rect 40460 17552 40466 17604
rect 48038 17552 48044 17604
rect 48096 17552 48102 17604
rect 18414 17524 18420 17536
rect 18327 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17524 18478 17536
rect 19150 17524 19156 17536
rect 18472 17496 19156 17524
rect 18472 17484 18478 17496
rect 19150 17484 19156 17496
rect 19208 17484 19214 17536
rect 19978 17524 19984 17536
rect 19891 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17524 20042 17536
rect 20254 17524 20260 17536
rect 20036 17496 20260 17524
rect 20036 17484 20042 17496
rect 20254 17484 20260 17496
rect 20312 17524 20318 17536
rect 20714 17524 20720 17536
rect 20312 17496 20720 17524
rect 20312 17484 20318 17496
rect 20714 17484 20720 17496
rect 20772 17524 20778 17536
rect 22281 17527 22339 17533
rect 22281 17524 22293 17527
rect 20772 17496 22293 17524
rect 20772 17484 20778 17496
rect 22281 17493 22293 17496
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 20622 17320 20628 17332
rect 19392 17292 20628 17320
rect 19392 17280 19398 17292
rect 20622 17280 20628 17292
rect 20680 17320 20686 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 20680 17292 21281 17320
rect 20680 17280 20686 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 21269 17283 21327 17289
rect 27341 17323 27399 17329
rect 27341 17289 27353 17323
rect 27387 17320 27399 17323
rect 28258 17320 28264 17332
rect 27387 17292 28264 17320
rect 27387 17289 27399 17292
rect 27341 17283 27399 17289
rect 28258 17280 28264 17292
rect 28316 17280 28322 17332
rect 45526 17292 46796 17320
rect 45526 17264 45554 17292
rect 18414 17252 18420 17264
rect 17144 17224 18420 17252
rect 17144 17193 17172 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 19797 17255 19855 17261
rect 19797 17252 19809 17255
rect 19484 17224 19809 17252
rect 19484 17212 19490 17224
rect 19797 17221 19809 17224
rect 19843 17221 19855 17255
rect 21913 17255 21971 17261
rect 21913 17252 21925 17255
rect 21022 17224 21925 17252
rect 19797 17215 19855 17221
rect 21913 17221 21925 17224
rect 21959 17221 21971 17255
rect 23658 17252 23664 17264
rect 23619 17224 23664 17252
rect 21913 17215 21971 17221
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 45462 17212 45468 17264
rect 45520 17224 45554 17264
rect 46768 17261 46796 17292
rect 46753 17255 46811 17261
rect 45520 17212 45526 17224
rect 46753 17221 46765 17255
rect 46799 17221 46811 17255
rect 46753 17215 46811 17221
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17678 17184 17684 17196
rect 17639 17156 17684 17184
rect 17129 17147 17187 17153
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 24762 17184 24768 17196
rect 24504 17156 24768 17184
rect 2406 17076 2412 17128
rect 2464 17116 2470 17128
rect 2464 17088 2774 17116
rect 2464 17076 2470 17088
rect 2746 17048 2774 17088
rect 3970 17076 3976 17128
rect 4028 17116 4034 17128
rect 6914 17116 6920 17128
rect 4028 17088 6920 17116
rect 4028 17076 4034 17088
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 19518 17116 19524 17128
rect 19479 17088 19524 17116
rect 19518 17076 19524 17088
rect 19576 17076 19582 17128
rect 23569 17119 23627 17125
rect 23569 17116 23581 17119
rect 22066 17088 23581 17116
rect 22066 17048 22094 17088
rect 23569 17085 23581 17088
rect 23615 17116 23627 17119
rect 23658 17116 23664 17128
rect 23615 17088 23664 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 23658 17076 23664 17088
rect 23716 17116 23722 17128
rect 24504 17116 24532 17156
rect 24762 17144 24768 17156
rect 24820 17144 24826 17196
rect 25222 17144 25228 17196
rect 25280 17184 25286 17196
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 25280 17156 25421 17184
rect 25280 17144 25286 17156
rect 25409 17153 25421 17156
rect 25455 17153 25467 17187
rect 25682 17184 25688 17196
rect 25643 17156 25688 17184
rect 25409 17147 25467 17153
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 26418 17144 26424 17196
rect 26476 17184 26482 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26476 17156 26985 17184
rect 26476 17144 26482 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 27154 17184 27160 17196
rect 27115 17156 27160 17184
rect 26973 17147 27031 17153
rect 27154 17144 27160 17156
rect 27212 17144 27218 17196
rect 45738 17144 45744 17196
rect 45796 17184 45802 17196
rect 47578 17184 47584 17196
rect 45796 17156 46138 17184
rect 47539 17156 47584 17184
rect 45796 17144 45802 17156
rect 47578 17144 47584 17156
rect 47636 17184 47642 17196
rect 47854 17184 47860 17196
rect 47636 17156 47860 17184
rect 47636 17144 47642 17156
rect 47854 17144 47860 17156
rect 47912 17144 47918 17196
rect 23716 17088 24532 17116
rect 24581 17119 24639 17125
rect 23716 17076 23722 17088
rect 24581 17085 24593 17119
rect 24627 17116 24639 17119
rect 24627 17088 25452 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 2746 17020 18092 17048
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1452 16952 2053 16980
rect 1452 16940 1458 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16724 16952 16957 16980
rect 16724 16940 16730 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17773 16983 17831 16989
rect 17773 16949 17785 16983
rect 17819 16980 17831 16983
rect 17954 16980 17960 16992
rect 17819 16952 17960 16980
rect 17819 16949 17831 16952
rect 17773 16943 17831 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18064 16980 18092 17020
rect 20805 17020 22094 17048
rect 20805 16980 20833 17020
rect 25424 16992 25452 17088
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25556 17088 25789 17116
rect 25556 17076 25562 17088
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 46198 17076 46204 17128
rect 46256 17116 46262 17128
rect 46256 17088 46301 17116
rect 46256 17076 46262 17088
rect 18064 16952 20833 16980
rect 25406 16940 25412 16992
rect 25464 16980 25470 16992
rect 25501 16983 25559 16989
rect 25501 16980 25513 16983
rect 25464 16952 25513 16980
rect 25464 16940 25470 16952
rect 25501 16949 25513 16952
rect 25547 16949 25559 16983
rect 25501 16943 25559 16949
rect 25869 16983 25927 16989
rect 25869 16949 25881 16983
rect 25915 16980 25927 16983
rect 26142 16980 26148 16992
rect 25915 16952 26148 16980
rect 25915 16949 25927 16952
rect 25869 16943 25927 16949
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 47670 16980 47676 16992
rect 47631 16952 47676 16980
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 19334 16776 19340 16788
rect 14384 16748 19340 16776
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 14384 16581 14412 16748
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 19889 16779 19947 16785
rect 19889 16776 19901 16779
rect 19576 16748 19901 16776
rect 19576 16736 19582 16748
rect 19889 16745 19901 16748
rect 19935 16745 19947 16779
rect 46566 16776 46572 16788
rect 19889 16739 19947 16745
rect 23400 16748 46572 16776
rect 16666 16640 16672 16652
rect 16627 16612 16672 16640
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 23400 16584 23428 16748
rect 46566 16736 46572 16748
rect 46624 16736 46630 16788
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 26016 16680 26924 16708
rect 26016 16668 26022 16680
rect 25501 16643 25559 16649
rect 25501 16609 25513 16643
rect 25547 16640 25559 16643
rect 26896 16640 26924 16680
rect 25547 16612 26832 16640
rect 26896 16612 27016 16640
rect 25547 16609 25559 16612
rect 25501 16603 25559 16609
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 19150 16532 19156 16584
rect 19208 16572 19214 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 19208 16544 19901 16572
rect 19208 16532 19214 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 23382 16572 23388 16584
rect 23295 16544 23388 16572
rect 19889 16535 19947 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 25958 16572 25964 16584
rect 25056 16544 25452 16572
rect 25919 16544 25964 16572
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2130 16504 2136 16516
rect 1627 16476 2136 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16504 14611 16507
rect 15010 16504 15016 16516
rect 14599 16476 15016 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16473 16267 16507
rect 16942 16504 16948 16516
rect 16903 16476 16948 16504
rect 16209 16467 16267 16473
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 16224 16436 16252 16467
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 18690 16504 18696 16516
rect 18603 16476 18696 16504
rect 18690 16464 18696 16476
rect 18748 16504 18754 16516
rect 25056 16504 25084 16544
rect 18748 16476 25084 16504
rect 25133 16507 25191 16513
rect 18748 16464 18754 16476
rect 25133 16473 25145 16507
rect 25179 16473 25191 16507
rect 25133 16467 25191 16473
rect 23474 16436 23480 16448
rect 3476 16408 16252 16436
rect 23435 16408 23480 16436
rect 3476 16396 3482 16408
rect 23474 16396 23480 16408
rect 23532 16396 23538 16448
rect 25148 16436 25176 16467
rect 25222 16464 25228 16516
rect 25280 16504 25286 16516
rect 25317 16507 25375 16513
rect 25317 16504 25329 16507
rect 25280 16476 25329 16504
rect 25280 16464 25286 16476
rect 25317 16473 25329 16476
rect 25363 16473 25375 16507
rect 25424 16504 25452 16544
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 26142 16572 26148 16584
rect 26103 16544 26148 16572
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26804 16581 26832 16612
rect 26988 16581 27016 16612
rect 27062 16600 27068 16652
rect 27120 16640 27126 16652
rect 27157 16643 27215 16649
rect 27157 16640 27169 16643
rect 27120 16612 27169 16640
rect 27120 16600 27126 16612
rect 27157 16609 27169 16612
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47026 16640 47032 16652
rect 46339 16612 47032 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47026 16600 47032 16612
rect 47084 16600 47090 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 26789 16575 26847 16581
rect 26789 16541 26801 16575
rect 26835 16541 26847 16575
rect 26789 16535 26847 16541
rect 26973 16575 27031 16581
rect 26973 16541 26985 16575
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 40034 16504 40040 16516
rect 25424 16476 26924 16504
rect 25317 16467 25375 16473
rect 25406 16436 25412 16448
rect 25148 16408 25412 16436
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 26326 16436 26332 16448
rect 26287 16408 26332 16436
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 26896 16436 26924 16476
rect 31726 16476 40040 16504
rect 31726 16436 31754 16476
rect 40034 16464 40040 16476
rect 40092 16464 40098 16516
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 26896 16408 31754 16436
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 15010 16232 15016 16244
rect 14971 16204 15016 16232
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17000 16204 17509 16232
rect 17000 16192 17006 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18564 16204 22094 16232
rect 18564 16192 18570 16204
rect 19150 16124 19156 16176
rect 19208 16164 19214 16176
rect 19208 16136 20944 16164
rect 19208 16124 19214 16136
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 14921 16099 14979 16105
rect 2087 16068 2774 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2746 15892 2774 16068
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15102 16096 15108 16108
rect 14967 16068 15108 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 18690 16096 18696 16108
rect 17175 16068 18696 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 19978 16096 19984 16108
rect 19659 16068 19984 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17310 16028 17316 16040
rect 17267 16000 17316 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 19444 16028 19472 16059
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20916 16105 20944 16136
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16065 20959 16099
rect 22066 16096 22094 16204
rect 25498 16192 25504 16244
rect 25556 16232 25562 16244
rect 25958 16232 25964 16244
rect 25556 16204 25964 16232
rect 25556 16192 25562 16204
rect 25958 16192 25964 16204
rect 26016 16232 26022 16244
rect 26145 16235 26203 16241
rect 26145 16232 26157 16235
rect 26016 16204 26157 16232
rect 26016 16192 26022 16204
rect 26145 16201 26157 16204
rect 26191 16201 26203 16235
rect 26145 16195 26203 16201
rect 26234 16192 26240 16244
rect 26292 16232 26298 16244
rect 26292 16204 26337 16232
rect 26292 16192 26298 16204
rect 26510 16192 26516 16244
rect 26568 16232 26574 16244
rect 26568 16204 28028 16232
rect 26568 16192 26574 16204
rect 23474 16164 23480 16176
rect 23435 16136 23480 16164
rect 23474 16124 23480 16136
rect 23532 16124 23538 16176
rect 26421 16167 26479 16173
rect 26421 16133 26433 16167
rect 26467 16164 26479 16167
rect 27893 16167 27951 16173
rect 27893 16164 27905 16167
rect 26467 16136 27905 16164
rect 26467 16133 26479 16136
rect 26421 16127 26479 16133
rect 23293 16099 23351 16105
rect 23293 16096 23305 16099
rect 22066 16068 23305 16096
rect 20901 16059 20959 16065
rect 23293 16065 23305 16068
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26142 16096 26148 16108
rect 26099 16068 26148 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 27062 16096 27068 16108
rect 27023 16068 27068 16096
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 27264 16105 27292 16136
rect 27893 16133 27905 16136
rect 27939 16133 27951 16167
rect 27893 16127 27951 16133
rect 27249 16099 27307 16105
rect 27249 16065 27261 16099
rect 27295 16065 27307 16099
rect 27798 16096 27804 16108
rect 27759 16068 27804 16096
rect 27249 16059 27307 16065
rect 27798 16056 27804 16068
rect 27856 16056 27862 16108
rect 28000 16105 28028 16204
rect 45462 16164 45468 16176
rect 43916 16136 45468 16164
rect 27985 16099 28043 16105
rect 27985 16065 27997 16099
rect 28031 16065 28043 16099
rect 40034 16096 40040 16108
rect 39995 16068 40040 16096
rect 27985 16059 28043 16065
rect 40034 16056 40040 16068
rect 40092 16056 40098 16108
rect 43916 16105 43944 16136
rect 45462 16124 45468 16136
rect 45520 16124 45526 16176
rect 46382 16164 46388 16176
rect 46295 16136 46388 16164
rect 46382 16124 46388 16136
rect 46440 16164 46446 16176
rect 47949 16167 48007 16173
rect 47949 16164 47961 16167
rect 46440 16136 47961 16164
rect 46440 16124 46446 16136
rect 47949 16133 47961 16136
rect 47995 16133 48007 16167
rect 47949 16127 48007 16133
rect 43901 16099 43959 16105
rect 43901 16065 43913 16099
rect 43947 16065 43959 16099
rect 43901 16059 43959 16065
rect 46753 16099 46811 16105
rect 46753 16065 46765 16099
rect 46799 16096 46811 16099
rect 47118 16096 47124 16108
rect 46799 16068 47124 16096
rect 46799 16065 46811 16068
rect 46753 16059 46811 16065
rect 47118 16056 47124 16068
rect 47176 16056 47182 16108
rect 47581 16099 47639 16105
rect 47581 16065 47593 16099
rect 47627 16096 47639 16099
rect 47670 16096 47676 16108
rect 47627 16068 47676 16096
rect 47627 16065 47639 16068
rect 47581 16059 47639 16065
rect 47670 16056 47676 16068
rect 47728 16056 47734 16108
rect 47765 16099 47823 16105
rect 47765 16065 47777 16099
rect 47811 16065 47823 16099
rect 47765 16059 47823 16065
rect 20438 16028 20444 16040
rect 19444 16000 20444 16028
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 25133 16031 25191 16037
rect 25133 15997 25145 16031
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 25869 16031 25927 16037
rect 25869 15997 25881 16031
rect 25915 16028 25927 16031
rect 40221 16031 40279 16037
rect 25915 16000 35894 16028
rect 25915 15997 25927 16000
rect 25869 15991 25927 15997
rect 2866 15892 2872 15904
rect 2746 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15892 2930 15904
rect 18598 15892 18604 15904
rect 2924 15864 18604 15892
rect 2924 15852 2930 15864
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 25148 15892 25176 15991
rect 27154 15920 27160 15972
rect 27212 15960 27218 15972
rect 27249 15963 27307 15969
rect 27249 15960 27261 15963
rect 27212 15932 27261 15960
rect 27212 15920 27218 15932
rect 27249 15929 27261 15932
rect 27295 15929 27307 15963
rect 35866 15960 35894 16000
rect 40221 15997 40233 16031
rect 40267 16028 40279 16031
rect 40494 16028 40500 16040
rect 40267 16000 40500 16028
rect 40267 15997 40279 16000
rect 40221 15991 40279 15997
rect 40494 15988 40500 16000
rect 40552 15988 40558 16040
rect 41874 16028 41880 16040
rect 41835 16000 41880 16028
rect 41874 15988 41880 16000
rect 41932 15988 41938 16040
rect 44082 16028 44088 16040
rect 44043 16000 44088 16028
rect 44082 15988 44088 16000
rect 44140 15988 44146 16040
rect 45462 16028 45468 16040
rect 45423 16000 45468 16028
rect 45462 15988 45468 16000
rect 45520 15988 45526 16040
rect 46198 16028 46204 16040
rect 46111 16000 46204 16028
rect 46198 15988 46204 16000
rect 46256 16028 46262 16040
rect 46845 16031 46903 16037
rect 46845 16028 46857 16031
rect 46256 16000 46857 16028
rect 46256 15988 46262 16000
rect 46845 15997 46857 16000
rect 46891 15997 46903 16031
rect 46845 15991 46903 15997
rect 46934 15988 46940 16040
rect 46992 16028 46998 16040
rect 47780 16028 47808 16059
rect 48038 16028 48044 16040
rect 46992 16000 48044 16028
rect 46992 15988 46998 16000
rect 48038 15988 48044 16000
rect 48096 15988 48102 16040
rect 46216 15960 46244 15988
rect 35866 15932 46244 15960
rect 27249 15923 27307 15929
rect 46658 15920 46664 15972
rect 46716 15960 46722 15972
rect 47029 15963 47087 15969
rect 47029 15960 47041 15963
rect 46716 15932 47041 15960
rect 46716 15920 46722 15932
rect 47029 15929 47041 15932
rect 47075 15929 47087 15963
rect 47029 15923 47087 15929
rect 46842 15892 46848 15904
rect 25148 15864 46848 15892
rect 46842 15852 46848 15864
rect 46900 15852 46906 15904
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 19797 15691 19855 15697
rect 19797 15657 19809 15691
rect 19843 15657 19855 15691
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 19797 15651 19855 15657
rect 19150 15552 19156 15564
rect 17144 15524 19156 15552
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1820 15456 2053 15484
rect 1820 15444 1826 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 2041 15447 2099 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 17144 15493 17172 15524
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15453 17187 15487
rect 17678 15484 17684 15496
rect 17639 15456 17684 15484
rect 17129 15447 17187 15453
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 19812 15484 19840 15651
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 25498 15688 25504 15700
rect 25459 15660 25504 15688
rect 25498 15648 25504 15660
rect 25556 15648 25562 15700
rect 27706 15648 27712 15700
rect 27764 15688 27770 15700
rect 27801 15691 27859 15697
rect 27801 15688 27813 15691
rect 27764 15660 27813 15688
rect 27764 15648 27770 15660
rect 27801 15657 27813 15660
rect 27847 15657 27859 15691
rect 40494 15688 40500 15700
rect 40455 15660 40500 15688
rect 27801 15651 27859 15657
rect 40494 15648 40500 15660
rect 40552 15648 40558 15700
rect 43993 15691 44051 15697
rect 43993 15657 44005 15691
rect 44039 15688 44051 15691
rect 44082 15688 44088 15700
rect 44039 15660 44088 15688
rect 44039 15657 44051 15660
rect 43993 15651 44051 15657
rect 44082 15648 44088 15660
rect 44140 15648 44146 15700
rect 45738 15688 45744 15700
rect 45699 15660 45744 15688
rect 45738 15648 45744 15660
rect 45796 15648 45802 15700
rect 47118 15648 47124 15700
rect 47176 15688 47182 15700
rect 47949 15691 48007 15697
rect 47949 15688 47961 15691
rect 47176 15660 47961 15688
rect 47176 15648 47182 15660
rect 47949 15657 47961 15660
rect 47995 15657 48007 15691
rect 47949 15651 48007 15657
rect 19978 15620 19984 15632
rect 19939 15592 19984 15620
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 46382 15552 46388 15564
rect 20588 15524 20760 15552
rect 20588 15512 20594 15524
rect 20254 15484 20260 15496
rect 19812 15456 20260 15484
rect 20254 15444 20260 15456
rect 20312 15484 20318 15496
rect 20732 15493 20760 15524
rect 45664 15524 46388 15552
rect 20625 15487 20683 15493
rect 20625 15484 20637 15487
rect 20312 15456 20637 15484
rect 20312 15444 20318 15456
rect 20625 15453 20637 15456
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15453 20775 15487
rect 20717 15447 20775 15453
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 19392 15388 19625 15416
rect 19392 15376 19398 15388
rect 19613 15385 19625 15388
rect 19659 15416 19671 15419
rect 20441 15419 20499 15425
rect 20441 15416 20453 15419
rect 19659 15388 20453 15416
rect 19659 15385 19671 15388
rect 19613 15379 19671 15385
rect 20441 15385 20453 15388
rect 20487 15416 20499 15419
rect 20530 15416 20536 15428
rect 20487 15388 20536 15416
rect 20487 15385 20499 15388
rect 20441 15379 20499 15385
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 15194 15348 15200 15360
rect 15155 15320 15200 15348
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 17129 15351 17187 15357
rect 17129 15348 17141 15351
rect 16724 15320 17141 15348
rect 16724 15308 16730 15320
rect 17129 15317 17141 15320
rect 17175 15317 17187 15351
rect 17129 15311 17187 15317
rect 17773 15351 17831 15357
rect 17773 15317 17785 15351
rect 17819 15348 17831 15351
rect 17954 15348 17960 15360
rect 17819 15320 17960 15348
rect 17819 15317 17831 15320
rect 17773 15311 17831 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 19823 15351 19881 15357
rect 19823 15317 19835 15351
rect 19869 15348 19881 15351
rect 20732 15348 20760 15447
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 21177 15487 21235 15493
rect 21177 15484 21189 15487
rect 20956 15456 21189 15484
rect 20956 15444 20962 15456
rect 21177 15453 21189 15456
rect 21223 15453 21235 15487
rect 21358 15484 21364 15496
rect 21319 15456 21364 15484
rect 21177 15447 21235 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 21591 15456 22201 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 22189 15447 22247 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15453 25651 15487
rect 25593 15447 25651 15453
rect 25222 15376 25228 15428
rect 25280 15416 25286 15428
rect 25608 15416 25636 15447
rect 26326 15444 26332 15496
rect 26384 15484 26390 15496
rect 26513 15487 26571 15493
rect 26513 15484 26525 15487
rect 26384 15456 26525 15484
rect 26384 15444 26390 15456
rect 26513 15453 26525 15456
rect 26559 15453 26571 15487
rect 27154 15484 27160 15496
rect 27115 15456 27160 15484
rect 26513 15447 26571 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 31205 15487 31263 15493
rect 31205 15453 31217 15487
rect 31251 15484 31263 15487
rect 40310 15484 40316 15496
rect 31251 15456 40316 15484
rect 31251 15453 31263 15456
rect 31205 15447 31263 15453
rect 40310 15444 40316 15456
rect 40368 15484 40374 15496
rect 40405 15487 40463 15493
rect 40405 15484 40417 15487
rect 40368 15456 40417 15484
rect 40368 15444 40374 15456
rect 40405 15453 40417 15456
rect 40451 15453 40463 15487
rect 40405 15447 40463 15453
rect 43530 15444 43536 15496
rect 43588 15484 43594 15496
rect 43898 15484 43904 15496
rect 43588 15456 43904 15484
rect 43588 15444 43594 15456
rect 43898 15444 43904 15456
rect 43956 15444 43962 15496
rect 45664 15493 45692 15524
rect 46382 15512 46388 15524
rect 46440 15512 46446 15564
rect 47136 15552 47164 15648
rect 46492 15524 47164 15552
rect 45649 15487 45707 15493
rect 45649 15453 45661 15487
rect 45695 15453 45707 15487
rect 45649 15447 45707 15453
rect 45833 15487 45891 15493
rect 45833 15453 45845 15487
rect 45879 15484 45891 15487
rect 46492 15484 46520 15524
rect 46658 15484 46664 15496
rect 45879 15456 46520 15484
rect 46619 15456 46664 15484
rect 45879 15453 45891 15456
rect 45833 15447 45891 15453
rect 46658 15444 46664 15456
rect 46716 15444 46722 15496
rect 47026 15484 47032 15496
rect 46987 15456 47032 15484
rect 47026 15444 47032 15456
rect 47084 15444 47090 15496
rect 47670 15444 47676 15496
rect 47728 15484 47734 15496
rect 47857 15487 47915 15493
rect 47857 15484 47869 15487
rect 47728 15456 47869 15484
rect 47728 15444 47734 15456
rect 47857 15453 47869 15456
rect 47903 15453 47915 15487
rect 48038 15484 48044 15496
rect 47999 15456 48044 15484
rect 47857 15447 47915 15453
rect 25280 15388 25636 15416
rect 25280 15376 25286 15388
rect 46290 15376 46296 15428
rect 46348 15416 46354 15428
rect 47397 15419 47455 15425
rect 47397 15416 47409 15419
rect 46348 15388 47409 15416
rect 46348 15376 46354 15388
rect 47397 15385 47409 15388
rect 47443 15385 47455 15419
rect 47872 15416 47900 15447
rect 48038 15444 48044 15456
rect 48096 15444 48102 15496
rect 47872 15388 48084 15416
rect 47397 15379 47455 15385
rect 48056 15360 48084 15388
rect 20806 15348 20812 15360
rect 19869 15320 20812 15348
rect 19869 15317 19881 15320
rect 19823 15311 19881 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 22005 15351 22063 15357
rect 22005 15317 22017 15351
rect 22051 15348 22063 15351
rect 22094 15348 22100 15360
rect 22051 15320 22100 15348
rect 22051 15317 22063 15320
rect 22005 15311 22063 15317
rect 22094 15308 22100 15320
rect 22152 15308 22158 15360
rect 30558 15308 30564 15360
rect 30616 15348 30622 15360
rect 31297 15351 31355 15357
rect 31297 15348 31309 15351
rect 30616 15320 31309 15348
rect 30616 15308 30622 15320
rect 31297 15317 31309 15320
rect 31343 15317 31355 15351
rect 31297 15311 31355 15317
rect 48038 15308 48044 15360
rect 48096 15308 48102 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 3234 15104 3240 15156
rect 3292 15144 3298 15156
rect 26145 15147 26203 15153
rect 3292 15116 26004 15144
rect 3292 15104 3298 15116
rect 17954 15036 17960 15088
rect 18012 15036 18018 15088
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 19521 15079 19579 15085
rect 19521 15076 19533 15079
rect 19484 15048 19533 15076
rect 19484 15036 19490 15048
rect 19521 15045 19533 15048
rect 19567 15045 19579 15079
rect 21726 15076 21732 15088
rect 20746 15048 21732 15076
rect 19521 15039 19579 15045
rect 21726 15036 21732 15048
rect 21784 15036 21790 15088
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 22152 15048 22197 15076
rect 22152 15036 22158 15048
rect 22830 15036 22836 15088
rect 22888 15036 22894 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 25976 15017 26004 15116
rect 26145 15113 26157 15147
rect 26191 15144 26203 15147
rect 26234 15144 26240 15156
rect 26191 15116 26240 15144
rect 26191 15113 26203 15116
rect 26145 15107 26203 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 27062 15144 27068 15156
rect 27023 15116 27068 15144
rect 27062 15104 27068 15116
rect 27120 15104 27126 15156
rect 47026 15104 47032 15156
rect 47084 15144 47090 15156
rect 47673 15147 47731 15153
rect 47673 15144 47685 15147
rect 47084 15116 47685 15144
rect 47084 15104 47090 15116
rect 47673 15113 47685 15116
rect 47719 15113 47731 15147
rect 47673 15107 47731 15113
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21048 14980 21833 15008
rect 21048 14968 21054 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26252 15008 26280 15104
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26252 14980 26985 15008
rect 26145 14971 26203 14977
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 46293 15011 46351 15017
rect 46293 14977 46305 15011
rect 46339 15008 46351 15011
rect 46382 15008 46388 15020
rect 46339 14980 46388 15008
rect 46339 14977 46351 14980
rect 46293 14971 46351 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 16945 14943 17003 14949
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17586 14940 17592 14952
rect 16991 14912 17592 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 19242 14940 19248 14952
rect 19203 14912 19248 14940
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 20530 14832 20536 14884
rect 20588 14872 20594 14884
rect 20993 14875 21051 14881
rect 20993 14872 21005 14875
rect 20588 14844 21005 14872
rect 20588 14832 20594 14844
rect 20993 14841 21005 14844
rect 21039 14841 21051 14875
rect 25976 14872 26004 14971
rect 26160 14940 26188 14971
rect 46382 14968 46388 14980
rect 46440 14968 46446 15020
rect 46477 15011 46535 15017
rect 46477 14977 46489 15011
rect 46523 14977 46535 15011
rect 46477 14971 46535 14977
rect 26510 14940 26516 14952
rect 26160 14912 26516 14940
rect 26510 14900 26516 14912
rect 26568 14940 26574 14952
rect 26786 14940 26792 14952
rect 26568 14912 26792 14940
rect 26568 14900 26574 14912
rect 26786 14900 26792 14912
rect 26844 14900 26850 14952
rect 27706 14900 27712 14952
rect 27764 14940 27770 14952
rect 43533 14943 43591 14949
rect 43533 14940 43545 14943
rect 27764 14912 43545 14940
rect 27764 14900 27770 14912
rect 43533 14909 43545 14912
rect 43579 14909 43591 14943
rect 43714 14940 43720 14952
rect 43675 14912 43720 14940
rect 43533 14903 43591 14909
rect 43714 14900 43720 14912
rect 43772 14900 43778 14952
rect 45094 14940 45100 14952
rect 45055 14912 45100 14940
rect 45094 14900 45100 14912
rect 45152 14900 45158 14952
rect 46492 14940 46520 14971
rect 46750 14968 46756 15020
rect 46808 15008 46814 15020
rect 47581 15011 47639 15017
rect 47581 15008 47593 15011
rect 46808 14980 47593 15008
rect 46808 14968 46814 14980
rect 47581 14977 47593 14980
rect 47627 14977 47639 15011
rect 47762 15008 47768 15020
rect 47723 14980 47768 15008
rect 47581 14971 47639 14977
rect 47762 14968 47768 14980
rect 47820 14968 47826 15020
rect 46842 14940 46848 14952
rect 46492 14912 46848 14940
rect 46842 14900 46848 14912
rect 46900 14900 46906 14952
rect 27798 14872 27804 14884
rect 25976 14844 27804 14872
rect 20993 14835 21051 14841
rect 27798 14832 27804 14844
rect 27856 14832 27862 14884
rect 18414 14804 18420 14816
rect 18375 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 23566 14804 23572 14816
rect 20312 14776 23572 14804
rect 20312 14764 20318 14776
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 46385 14807 46443 14813
rect 46385 14773 46397 14807
rect 46431 14804 46443 14807
rect 46474 14804 46480 14816
rect 46431 14776 46480 14804
rect 46431 14773 46443 14776
rect 46385 14767 46443 14773
rect 46474 14764 46480 14776
rect 46532 14764 46538 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 17586 14600 17592 14612
rect 17547 14572 17592 14600
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19484 14572 19625 14600
rect 19484 14560 19490 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 20070 14600 20076 14612
rect 19843 14572 20076 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 21177 14603 21235 14609
rect 21177 14569 21189 14603
rect 21223 14600 21235 14603
rect 21358 14600 21364 14612
rect 21223 14572 21364 14600
rect 21223 14569 21235 14572
rect 21177 14563 21235 14569
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 21726 14600 21732 14612
rect 21687 14572 21732 14600
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 22830 14560 22836 14612
rect 22888 14600 22894 14612
rect 22925 14603 22983 14609
rect 22925 14600 22937 14603
rect 22888 14572 22937 14600
rect 22888 14560 22894 14572
rect 22925 14569 22937 14572
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 43625 14603 43683 14609
rect 43625 14569 43637 14603
rect 43671 14600 43683 14603
rect 43714 14600 43720 14612
rect 43671 14572 43720 14600
rect 43671 14569 43683 14572
rect 43625 14563 43683 14569
rect 43714 14560 43720 14572
rect 43772 14560 43778 14612
rect 47397 14603 47455 14609
rect 47397 14569 47409 14603
rect 47443 14600 47455 14603
rect 47762 14600 47768 14612
rect 47443 14572 47768 14600
rect 47443 14569 47455 14572
rect 47397 14563 47455 14569
rect 47762 14560 47768 14572
rect 47820 14560 47826 14612
rect 3510 14492 3516 14544
rect 3568 14532 3574 14544
rect 17957 14535 18015 14541
rect 3568 14504 15516 14532
rect 3568 14492 3574 14504
rect 15194 14464 15200 14476
rect 15155 14436 15200 14464
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15488 14473 15516 14504
rect 17957 14501 17969 14535
rect 18003 14532 18015 14535
rect 19978 14532 19984 14544
rect 18003 14504 19984 14532
rect 18003 14501 18015 14504
rect 17957 14495 18015 14501
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 30377 14467 30435 14473
rect 30377 14464 30389 14467
rect 23624 14436 30389 14464
rect 23624 14424 23630 14436
rect 30377 14433 30389 14436
rect 30423 14433 30435 14467
rect 30558 14464 30564 14476
rect 30519 14436 30564 14464
rect 30377 14427 30435 14433
rect 30558 14424 30564 14436
rect 30616 14424 30622 14476
rect 46750 14464 46756 14476
rect 46308 14436 46756 14464
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15028 14328 15056 14359
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17368 14368 17785 14396
rect 17368 14356 17374 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18414 14396 18420 14408
rect 18095 14368 18420 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18064 14328 18092 14359
rect 18414 14356 18420 14368
rect 18472 14396 18478 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 18472 14368 19472 14396
rect 18472 14356 18478 14368
rect 19444 14337 19472 14368
rect 20272 14368 21005 14396
rect 20272 14340 20300 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 21818 14396 21824 14408
rect 21683 14368 21824 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 21818 14356 21824 14368
rect 21876 14396 21882 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 21876 14368 22845 14396
rect 21876 14356 21882 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 43530 14396 43536 14408
rect 43491 14368 43536 14396
rect 22833 14359 22891 14365
rect 43530 14356 43536 14368
rect 43588 14356 43594 14408
rect 46308 14405 46336 14436
rect 46750 14424 46756 14436
rect 46808 14424 46814 14476
rect 46293 14399 46351 14405
rect 46293 14365 46305 14399
rect 46339 14365 46351 14399
rect 46474 14396 46480 14408
rect 46435 14368 46480 14396
rect 46293 14359 46351 14365
rect 46474 14356 46480 14368
rect 46532 14356 46538 14408
rect 46569 14399 46627 14405
rect 46569 14365 46581 14399
rect 46615 14396 46627 14399
rect 46658 14396 46664 14408
rect 46615 14368 46664 14396
rect 46615 14365 46627 14368
rect 46569 14359 46627 14365
rect 46658 14356 46664 14368
rect 46716 14356 46722 14408
rect 46842 14356 46848 14408
rect 46900 14396 46906 14408
rect 47029 14399 47087 14405
rect 47029 14396 47041 14399
rect 46900 14368 47041 14396
rect 46900 14356 46906 14368
rect 47029 14365 47041 14368
rect 47075 14365 47087 14399
rect 47029 14359 47087 14365
rect 47213 14399 47271 14405
rect 47213 14365 47225 14399
rect 47259 14365 47271 14399
rect 47213 14359 47271 14365
rect 15028 14300 18092 14328
rect 19429 14331 19487 14337
rect 19429 14297 19441 14331
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 19645 14331 19703 14337
rect 19645 14297 19657 14331
rect 19691 14328 19703 14331
rect 20254 14328 20260 14340
rect 19691 14300 20260 14328
rect 19691 14297 19703 14300
rect 19645 14291 19703 14297
rect 20254 14288 20260 14300
rect 20312 14288 20318 14340
rect 20806 14328 20812 14340
rect 20767 14300 20812 14328
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 32214 14328 32220 14340
rect 32175 14300 32220 14328
rect 32214 14288 32220 14300
rect 32272 14288 32278 14340
rect 46382 14288 46388 14340
rect 46440 14328 46446 14340
rect 47228 14328 47256 14359
rect 46440 14300 47256 14328
rect 46440 14288 46446 14300
rect 46106 14260 46112 14272
rect 46067 14232 46112 14260
rect 46106 14220 46112 14232
rect 46164 14220 46170 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 41046 14056 41052 14068
rect 2188 14028 41052 14056
rect 2188 14016 2194 14028
rect 41046 14016 41052 14028
rect 41104 14016 41110 14068
rect 46661 14059 46719 14065
rect 46661 14025 46673 14059
rect 46707 14056 46719 14059
rect 46750 14056 46756 14068
rect 46707 14028 46756 14056
rect 46707 14025 46719 14028
rect 46661 14019 46719 14025
rect 46750 14016 46756 14028
rect 46808 14016 46814 14068
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19300 13960 19441 13988
rect 19300 13948 19306 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 20898 13988 20904 14000
rect 20859 13960 20904 13988
rect 19429 13951 19487 13957
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 45526 13960 47624 13988
rect 19150 13920 19156 13932
rect 19111 13892 19156 13920
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 20806 13920 20812 13932
rect 20767 13892 20812 13920
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13889 21051 13923
rect 20993 13883 21051 13889
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 21008 13852 21036 13883
rect 20312 13824 21036 13852
rect 20312 13812 20318 13824
rect 43530 13812 43536 13864
rect 43588 13852 43594 13864
rect 45526 13852 45554 13960
rect 45649 13923 45707 13929
rect 45649 13889 45661 13923
rect 45695 13920 45707 13923
rect 45738 13920 45744 13932
rect 45695 13892 45744 13920
rect 45695 13889 45707 13892
rect 45649 13883 45707 13889
rect 45738 13880 45744 13892
rect 45796 13880 45802 13932
rect 46014 13920 46020 13932
rect 45833 13889 45891 13895
rect 45975 13892 46020 13920
rect 45833 13864 45845 13889
rect 45879 13864 45891 13889
rect 46014 13880 46020 13892
rect 46072 13880 46078 13932
rect 46106 13880 46112 13932
rect 46164 13920 46170 13932
rect 46164 13892 46209 13920
rect 46164 13880 46170 13892
rect 46382 13880 46388 13932
rect 46440 13920 46446 13932
rect 46569 13923 46627 13929
rect 46569 13920 46581 13923
rect 46440 13892 46581 13920
rect 46440 13880 46446 13892
rect 46569 13889 46581 13892
rect 46615 13889 46627 13923
rect 46750 13920 46756 13932
rect 46711 13892 46756 13920
rect 46569 13883 46627 13889
rect 46750 13880 46756 13892
rect 46808 13880 46814 13932
rect 47596 13929 47624 13960
rect 47581 13923 47639 13929
rect 47581 13889 47593 13923
rect 47627 13889 47639 13923
rect 47581 13883 47639 13889
rect 43588 13824 45554 13852
rect 43588 13812 43594 13824
rect 45830 13812 45836 13864
rect 45888 13812 45894 13864
rect 46474 13812 46480 13864
rect 46532 13852 46538 13864
rect 47673 13855 47731 13861
rect 47673 13852 47685 13855
rect 46532 13824 47685 13852
rect 46532 13812 46538 13824
rect 47673 13821 47685 13824
rect 47719 13821 47731 13855
rect 47673 13815 47731 13821
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 5442 13716 5448 13728
rect 4028 13688 5448 13716
rect 4028 13676 4034 13688
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13308 20223 13311
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 20211 13280 20821 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20809 13277 20821 13280
rect 20855 13308 20867 13311
rect 23382 13308 23388 13320
rect 20855 13280 23388 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 46106 13308 46112 13320
rect 46067 13280 46112 13308
rect 46106 13268 46112 13280
rect 46164 13268 46170 13320
rect 46658 13308 46664 13320
rect 46619 13280 46664 13308
rect 46658 13268 46664 13280
rect 46716 13268 46722 13320
rect 46934 13268 46940 13320
rect 46992 13308 46998 13320
rect 48133 13311 48191 13317
rect 48133 13308 48145 13311
rect 46992 13280 48145 13308
rect 46992 13268 46998 13280
rect 48133 13277 48145 13280
rect 48179 13277 48191 13311
rect 48133 13271 48191 13277
rect 47486 13240 47492 13252
rect 47447 13212 47492 13240
rect 47486 13200 47492 13212
rect 47544 13200 47550 13252
rect 20254 13172 20260 13184
rect 20215 13144 20260 13172
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20898 13172 20904 13184
rect 20859 13144 20904 13172
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 46658 12968 46664 12980
rect 46619 12940 46664 12968
rect 46658 12928 46664 12940
rect 46716 12928 46722 12980
rect 19613 12903 19671 12909
rect 19613 12869 19625 12903
rect 19659 12900 19671 12903
rect 20254 12900 20260 12912
rect 19659 12872 20260 12900
rect 19659 12869 19671 12872
rect 19613 12863 19671 12869
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 45005 12903 45063 12909
rect 45005 12869 45017 12903
rect 45051 12900 45063 12903
rect 45830 12900 45836 12912
rect 45051 12872 45836 12900
rect 45051 12869 45063 12872
rect 45005 12863 45063 12869
rect 45830 12860 45836 12872
rect 45888 12900 45894 12912
rect 45888 12872 46612 12900
rect 45888 12860 45894 12872
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 46584 12841 46612 12872
rect 44913 12835 44971 12841
rect 44913 12801 44925 12835
rect 44959 12801 44971 12835
rect 44913 12795 44971 12801
rect 45097 12835 45155 12841
rect 45097 12801 45109 12835
rect 45143 12832 45155 12835
rect 45741 12835 45799 12841
rect 45143 12804 45600 12832
rect 45143 12801 45155 12804
rect 45097 12795 45155 12801
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 20622 12764 20628 12776
rect 19475 12736 20628 12764
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 21266 12764 21272 12776
rect 21227 12736 21272 12764
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 44928 12696 44956 12795
rect 45572 12773 45600 12804
rect 45741 12801 45753 12835
rect 45787 12832 45799 12835
rect 45925 12835 45983 12841
rect 45787 12804 45876 12832
rect 45787 12801 45799 12804
rect 45741 12795 45799 12801
rect 45848 12776 45876 12804
rect 45925 12801 45937 12835
rect 45971 12832 45983 12835
rect 46385 12835 46443 12841
rect 46385 12832 46397 12835
rect 45971 12804 46397 12832
rect 45971 12801 45983 12804
rect 45925 12795 45983 12801
rect 46385 12801 46397 12804
rect 46431 12801 46443 12835
rect 46385 12795 46443 12801
rect 46569 12835 46627 12841
rect 46569 12801 46581 12835
rect 46615 12801 46627 12835
rect 46569 12795 46627 12801
rect 45557 12767 45615 12773
rect 45557 12733 45569 12767
rect 45603 12764 45615 12767
rect 45603 12736 45784 12764
rect 45603 12733 45615 12736
rect 45557 12727 45615 12733
rect 45756 12708 45784 12736
rect 45830 12724 45836 12776
rect 45888 12724 45894 12776
rect 44928 12668 45554 12696
rect 45526 12640 45554 12668
rect 45738 12656 45744 12708
rect 45796 12656 45802 12708
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 34790 12628 34796 12640
rect 1627 12600 34796 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 34790 12588 34796 12600
rect 34848 12588 34854 12640
rect 45526 12600 45560 12640
rect 45554 12588 45560 12600
rect 45612 12628 45618 12640
rect 45848 12628 45876 12724
rect 45612 12600 45876 12628
rect 45612 12588 45618 12600
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 45741 12427 45799 12433
rect 45741 12393 45753 12427
rect 45787 12424 45799 12427
rect 46014 12424 46020 12436
rect 45787 12396 46020 12424
rect 45787 12393 45799 12396
rect 45741 12387 45799 12393
rect 46014 12384 46020 12396
rect 46072 12384 46078 12436
rect 46934 12356 46940 12368
rect 46308 12328 46940 12356
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19521 12291 19579 12297
rect 19521 12288 19533 12291
rect 19484 12260 19533 12288
rect 19484 12248 19490 12260
rect 19521 12257 19533 12260
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12288 19763 12291
rect 20898 12288 20904 12300
rect 19751 12260 20904 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 46308 12297 46336 12328
rect 46934 12316 46940 12328
rect 46992 12316 46998 12368
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12257 46351 12291
rect 46474 12288 46480 12300
rect 46435 12260 46480 12288
rect 46293 12251 46351 12257
rect 46474 12248 46480 12260
rect 46532 12248 46538 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 45554 12180 45560 12232
rect 45612 12220 45618 12232
rect 45649 12223 45707 12229
rect 45649 12220 45661 12223
rect 45612 12192 45661 12220
rect 45612 12180 45618 12192
rect 45649 12189 45661 12192
rect 45695 12189 45707 12223
rect 45649 12183 45707 12189
rect 14826 12112 14832 12164
rect 14884 12152 14890 12164
rect 21361 12155 21419 12161
rect 21361 12152 21373 12155
rect 14884 12124 21373 12152
rect 14884 12112 14890 12124
rect 21361 12121 21373 12124
rect 21407 12121 21419 12155
rect 45664 12152 45692 12183
rect 45738 12180 45744 12232
rect 45796 12220 45802 12232
rect 45833 12223 45891 12229
rect 45833 12220 45845 12223
rect 45796 12192 45845 12220
rect 45796 12180 45802 12192
rect 45833 12189 45845 12192
rect 45879 12189 45891 12223
rect 45833 12183 45891 12189
rect 46290 12152 46296 12164
rect 45664 12124 46296 12152
rect 21361 12115 21419 12121
rect 46290 12112 46296 12124
rect 46348 12112 46354 12164
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 46106 11812 46112 11824
rect 46067 11784 46112 11812
rect 46106 11772 46112 11784
rect 46164 11772 46170 11824
rect 46014 11676 46020 11688
rect 45975 11648 46020 11676
rect 46014 11636 46020 11648
rect 46072 11636 46078 11688
rect 46290 11676 46296 11688
rect 46251 11648 46296 11676
rect 46290 11636 46296 11648
rect 46348 11636 46354 11688
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 47670 11064 47676 11076
rect 46523 11036 47676 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 47670 11024 47676 11036
rect 47728 11024 47734 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 47670 10792 47676 10804
rect 47631 10764 47676 10792
rect 47670 10752 47676 10764
rect 47728 10752 47734 10804
rect 41046 10616 41052 10668
rect 41104 10656 41110 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 41104 10628 47593 10656
rect 41104 10616 41110 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 4798 10452 4804 10464
rect 2832 10424 4804 10452
rect 2832 10412 2838 10424
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 46290 10412 46296 10464
rect 46348 10452 46354 10464
rect 47029 10455 47087 10461
rect 47029 10452 47041 10455
rect 46348 10424 47041 10452
rect 46348 10412 46354 10424
rect 47029 10421 47041 10424
rect 47075 10421 47087 10455
rect 47029 10415 47087 10421
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 19116 10084 19257 10112
rect 19116 10072 19122 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 19245 10075 19303 10081
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 19426 9976 19432 9988
rect 19387 9948 19432 9976
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 20990 9936 20996 9988
rect 21048 9976 21054 9988
rect 21085 9979 21143 9985
rect 21085 9976 21097 9979
rect 21048 9948 21097 9976
rect 21048 9936 21054 9948
rect 21085 9945 21097 9948
rect 21131 9945 21143 9979
rect 21085 9939 21143 9945
rect 46477 9979 46535 9985
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 19426 9636 19432 9648
rect 19291 9608 19432 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 47670 9636 47676 9648
rect 47631 9608 47676 9636
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 19153 9571 19211 9577
rect 19153 9568 19165 9571
rect 18288 9540 19165 9568
rect 18288 9528 18294 9540
rect 19153 9537 19165 9540
rect 19199 9568 19211 9571
rect 42702 9568 42708 9580
rect 19199 9540 42708 9568
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 42702 9528 42708 9540
rect 42760 9528 42766 9580
rect 46842 9528 46848 9580
rect 46900 9568 46906 9580
rect 47029 9571 47087 9577
rect 47029 9568 47041 9571
rect 46900 9540 47041 9568
rect 46900 9528 46906 9540
rect 47029 9537 47041 9540
rect 47075 9537 47087 9571
rect 47029 9531 47087 9537
rect 47581 9571 47639 9577
rect 47581 9537 47593 9571
rect 47627 9568 47639 9571
rect 47854 9568 47860 9580
rect 47627 9540 47860 9568
rect 47627 9537 47639 9540
rect 47581 9531 47639 9537
rect 45370 9460 45376 9512
rect 45428 9500 45434 9512
rect 47596 9500 47624 9531
rect 47854 9528 47860 9540
rect 47912 9528 47918 9580
rect 45428 9472 47624 9500
rect 45428 9460 45434 9472
rect 46106 9392 46112 9444
rect 46164 9432 46170 9444
rect 46845 9435 46903 9441
rect 46845 9432 46857 9435
rect 46164 9404 46857 9432
rect 46164 9392 46170 9404
rect 46845 9401 46857 9404
rect 46891 9401 46903 9435
rect 46845 9395 46903 9401
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 47302 8956 47308 8968
rect 47263 8928 47308 8956
rect 47302 8916 47308 8928
rect 47360 8916 47366 8968
rect 47394 8916 47400 8968
rect 47452 8956 47458 8968
rect 47581 8959 47639 8965
rect 47581 8956 47593 8959
rect 47452 8928 47593 8956
rect 47452 8916 47458 8928
rect 47581 8925 47593 8928
rect 47627 8925 47639 8959
rect 47581 8919 47639 8925
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 47762 8548 47768 8560
rect 47723 8520 47768 8548
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 38010 8304 38016 8356
rect 38068 8344 38074 8356
rect 47949 8347 48007 8353
rect 47949 8344 47961 8347
rect 38068 8316 47961 8344
rect 38068 8304 38074 8316
rect 47949 8313 47961 8316
rect 47995 8313 48007 8347
rect 47949 8307 48007 8313
rect 41874 8236 41880 8288
rect 41932 8276 41938 8288
rect 45554 8276 45560 8288
rect 41932 8248 45560 8276
rect 41932 8236 41938 8248
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 46198 7896 46204 7948
rect 46256 7936 46262 7948
rect 46293 7939 46351 7945
rect 46293 7936 46305 7939
rect 46256 7908 46305 7936
rect 46256 7896 46262 7908
rect 46293 7905 46305 7908
rect 46339 7905 46351 7939
rect 46293 7899 46351 7905
rect 46477 7939 46535 7945
rect 46477 7905 46489 7939
rect 46523 7936 46535 7939
rect 47394 7936 47400 7948
rect 46523 7908 47400 7936
rect 46523 7905 46535 7908
rect 46477 7899 46535 7905
rect 47394 7896 47400 7908
rect 47452 7896 47458 7948
rect 47946 7936 47952 7948
rect 47907 7908 47952 7936
rect 47946 7896 47952 7908
rect 48004 7896 48010 7948
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 48130 7392 48136 7404
rect 48091 7364 48136 7392
rect 48130 7352 48136 7364
rect 48188 7352 48194 7404
rect 47118 7148 47124 7200
rect 47176 7188 47182 7200
rect 47949 7191 48007 7197
rect 47949 7188 47961 7191
rect 47176 7160 47961 7188
rect 47176 7148 47182 7160
rect 47949 7157 47961 7160
rect 47995 7157 48007 7191
rect 47949 7151 48007 7157
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 47118 6848 47124 6860
rect 47079 6820 47124 6848
rect 47118 6808 47124 6820
rect 47176 6808 47182 6860
rect 48038 6848 48044 6860
rect 47999 6820 48044 6848
rect 48038 6808 48044 6820
rect 48096 6808 48102 6860
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 47213 6715 47271 6721
rect 47213 6712 47225 6715
rect 1912 6684 26234 6712
rect 1912 6672 1918 6684
rect 26206 6644 26234 6684
rect 41386 6684 47225 6712
rect 41386 6644 41414 6684
rect 47213 6681 47225 6684
rect 47259 6681 47271 6715
rect 47213 6675 47271 6681
rect 26206 6616 41414 6644
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 46477 6307 46535 6313
rect 46477 6273 46489 6307
rect 46523 6304 46535 6307
rect 46750 6304 46756 6316
rect 46523 6276 46756 6304
rect 46523 6273 46535 6276
rect 46477 6267 46535 6273
rect 46750 6264 46756 6276
rect 46808 6264 46814 6316
rect 48130 6304 48136 6316
rect 48091 6276 48136 6304
rect 48130 6264 48136 6276
rect 48188 6264 48194 6316
rect 46198 6236 46204 6248
rect 46159 6208 46204 6236
rect 46198 6196 46204 6208
rect 46256 6196 46262 6248
rect 47946 6100 47952 6112
rect 47907 6072 47952 6100
rect 47946 6060 47952 6072
rect 48004 6060 48010 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 41230 5720 41236 5772
rect 41288 5760 41294 5772
rect 46293 5763 46351 5769
rect 46293 5760 46305 5763
rect 41288 5732 46305 5760
rect 41288 5720 41294 5732
rect 46293 5729 46305 5732
rect 46339 5729 46351 5763
rect 47854 5760 47860 5772
rect 47815 5732 47860 5760
rect 46293 5723 46351 5729
rect 47854 5720 47860 5732
rect 47912 5720 47918 5772
rect 46198 5584 46204 5636
rect 46256 5624 46262 5636
rect 46477 5627 46535 5633
rect 46477 5624 46489 5627
rect 46256 5596 46489 5624
rect 46256 5584 46262 5596
rect 46477 5593 46489 5596
rect 46523 5593 46535 5627
rect 46477 5587 46535 5593
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 45646 5352 45652 5364
rect 31726 5324 45652 5352
rect 19613 5287 19671 5293
rect 19613 5284 19625 5287
rect 18248 5256 19625 5284
rect 18248 5225 18276 5256
rect 19613 5253 19625 5256
rect 19659 5253 19671 5287
rect 23474 5284 23480 5296
rect 19613 5247 19671 5253
rect 22480 5256 23480 5284
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18322 5176 18328 5228
rect 18380 5216 18386 5228
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18380 5188 18889 5216
rect 18380 5176 18386 5188
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 19521 5219 19579 5225
rect 19521 5216 19533 5219
rect 19024 5188 19533 5216
rect 19024 5176 19030 5188
rect 19521 5185 19533 5188
rect 19567 5185 19579 5219
rect 20254 5216 20260 5228
rect 20215 5188 20260 5216
rect 19521 5179 19579 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20901 5219 20959 5225
rect 20901 5185 20913 5219
rect 20947 5216 20959 5219
rect 21726 5216 21732 5228
rect 20947 5188 21732 5216
rect 20947 5185 20959 5188
rect 20901 5179 20959 5185
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5216 21879 5219
rect 21910 5216 21916 5228
rect 21867 5188 21916 5216
rect 21867 5185 21879 5188
rect 21821 5179 21879 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 22480 5225 22508 5256
rect 23474 5244 23480 5256
rect 23532 5244 23538 5296
rect 31205 5287 31263 5293
rect 31205 5253 31217 5287
rect 31251 5284 31263 5287
rect 31726 5284 31754 5324
rect 45646 5312 45652 5324
rect 45704 5312 45710 5364
rect 46014 5284 46020 5296
rect 31251 5256 31754 5284
rect 45975 5256 46020 5284
rect 31251 5253 31263 5256
rect 31205 5247 31263 5253
rect 46014 5244 46020 5256
rect 46072 5244 46078 5296
rect 46109 5287 46167 5293
rect 46109 5253 46121 5287
rect 46155 5284 46167 5287
rect 47946 5284 47952 5296
rect 46155 5256 47952 5284
rect 46155 5253 46167 5256
rect 46109 5247 46167 5253
rect 47946 5244 47952 5256
rect 48004 5244 48010 5296
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 23109 5219 23167 5225
rect 23109 5185 23121 5219
rect 23155 5216 23167 5219
rect 23842 5216 23848 5228
rect 23155 5188 23848 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 43254 5176 43260 5228
rect 43312 5216 43318 5228
rect 45281 5219 45339 5225
rect 45281 5216 45293 5219
rect 43312 5188 45293 5216
rect 43312 5176 43318 5188
rect 45281 5185 45293 5188
rect 45327 5185 45339 5219
rect 47854 5216 47860 5228
rect 47815 5188 47860 5216
rect 45281 5179 45339 5185
rect 47854 5176 47860 5188
rect 47912 5176 47918 5228
rect 48038 5176 48044 5228
rect 48096 5176 48102 5228
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 29365 5151 29423 5157
rect 29365 5148 29377 5151
rect 4120 5120 29377 5148
rect 4120 5108 4126 5120
rect 29365 5117 29377 5120
rect 29411 5117 29423 5151
rect 29365 5111 29423 5117
rect 29549 5151 29607 5157
rect 29549 5117 29561 5151
rect 29595 5148 29607 5151
rect 30006 5148 30012 5160
rect 29595 5120 30012 5148
rect 29595 5117 29607 5120
rect 29549 5111 29607 5117
rect 30006 5108 30012 5120
rect 30064 5108 30070 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48056 5148 48084 5176
rect 46891 5120 48084 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18969 5083 19027 5089
rect 18969 5080 18981 5083
rect 18012 5052 18981 5080
rect 18012 5040 18018 5052
rect 18969 5049 18981 5052
rect 19015 5049 19027 5083
rect 18969 5043 19027 5049
rect 28718 5040 28724 5092
rect 28776 5080 28782 5092
rect 48041 5083 48099 5089
rect 48041 5080 48053 5083
rect 28776 5052 48053 5080
rect 28776 5040 28782 5052
rect 48041 5049 48053 5052
rect 48087 5049 48099 5083
rect 48041 5043 48099 5049
rect 18325 5015 18383 5021
rect 18325 4981 18337 5015
rect 18371 5012 18383 5015
rect 18874 5012 18880 5024
rect 18371 4984 18880 5012
rect 18371 4981 18383 4984
rect 18325 4975 18383 4981
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20993 5015 21051 5021
rect 20993 4981 21005 5015
rect 21039 5012 21051 5015
rect 21818 5012 21824 5024
rect 21039 4984 21824 5012
rect 21039 4981 21051 4984
rect 20993 4975 21051 4981
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22370 5012 22376 5024
rect 21959 4984 22376 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 23106 5012 23112 5024
rect 22603 4984 23112 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 23198 4972 23204 5024
rect 23256 5012 23262 5024
rect 45373 5015 45431 5021
rect 23256 4984 23301 5012
rect 23256 4972 23262 4984
rect 45373 4981 45385 5015
rect 45419 5012 45431 5015
rect 45922 5012 45928 5024
rect 45419 4984 45928 5012
rect 45419 4981 45431 4984
rect 45373 4975 45431 4981
rect 45922 4972 45928 4984
rect 45980 4972 45986 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 18322 4808 18328 4820
rect 18283 4780 18328 4808
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 20312 4780 21281 4808
rect 20312 4768 20318 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21784 4780 21925 4808
rect 21784 4768 21790 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 21913 4771 21971 4777
rect 47486 4740 47492 4752
rect 45756 4712 47492 4740
rect 20346 4632 20352 4684
rect 20404 4672 20410 4684
rect 45756 4681 45784 4712
rect 47486 4700 47492 4712
rect 47544 4700 47550 4752
rect 45741 4675 45799 4681
rect 20404 4644 21864 4672
rect 20404 4632 20410 4644
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4604 19303 4607
rect 19426 4604 19432 4616
rect 19291 4576 19432 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 18248 4536 18276 4567
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 19978 4604 19984 4616
rect 19935 4576 19984 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20530 4604 20536 4616
rect 20491 4576 20536 4604
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 21836 4613 21864 4644
rect 45741 4641 45753 4675
rect 45787 4641 45799 4675
rect 45922 4672 45928 4684
rect 45883 4644 45928 4672
rect 45741 4635 45799 4641
rect 45922 4632 45928 4644
rect 45980 4632 45986 4684
rect 46934 4672 46940 4684
rect 46895 4644 46940 4672
rect 46934 4632 46940 4644
rect 46992 4632 46998 4684
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 21177 4607 21235 4613
rect 21177 4604 21189 4607
rect 20671 4576 21189 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 21177 4573 21189 4576
rect 21223 4573 21235 4607
rect 21177 4567 21235 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4573 21879 4607
rect 22462 4604 22468 4616
rect 22423 4576 22468 4604
rect 21821 4567 21879 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 23106 4604 23112 4616
rect 23067 4576 23112 4604
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 42426 4564 42432 4616
rect 42484 4604 42490 4616
rect 42521 4607 42579 4613
rect 42521 4604 42533 4607
rect 42484 4576 42533 4604
rect 42484 4564 42490 4576
rect 42521 4573 42533 4576
rect 42567 4573 42579 4607
rect 42521 4567 42579 4573
rect 43806 4564 43812 4616
rect 43864 4604 43870 4616
rect 44085 4607 44143 4613
rect 44085 4604 44097 4607
rect 43864 4576 44097 4604
rect 43864 4564 43870 4576
rect 44085 4573 44097 4576
rect 44131 4573 44143 4607
rect 44085 4567 44143 4573
rect 45186 4564 45192 4616
rect 45244 4604 45250 4616
rect 45281 4607 45339 4613
rect 45281 4604 45293 4607
rect 45244 4576 45293 4604
rect 45244 4564 45250 4576
rect 45281 4573 45293 4576
rect 45327 4573 45339 4607
rect 45281 4567 45339 4573
rect 20070 4536 20076 4548
rect 18248 4508 20076 4536
rect 20070 4496 20076 4508
rect 20128 4496 20134 4548
rect 19334 4468 19340 4480
rect 19295 4440 19340 4468
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19981 4471 20039 4477
rect 19981 4437 19993 4471
rect 20027 4468 20039 4471
rect 20530 4468 20536 4480
rect 20027 4440 20536 4468
rect 20027 4437 20039 4440
rect 19981 4431 20039 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 22557 4471 22615 4477
rect 22557 4437 22569 4471
rect 22603 4468 22615 4471
rect 23106 4468 23112 4480
rect 22603 4440 23112 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 23201 4471 23259 4477
rect 23201 4437 23213 4471
rect 23247 4468 23259 4471
rect 23750 4468 23756 4480
rect 23247 4440 23756 4468
rect 23247 4437 23259 4440
rect 23201 4431 23259 4437
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 43070 4428 43076 4480
rect 43128 4468 43134 4480
rect 43901 4471 43959 4477
rect 43901 4468 43913 4471
rect 43128 4440 43913 4468
rect 43128 4428 43134 4440
rect 43901 4437 43913 4440
rect 43947 4437 43959 4471
rect 43901 4431 43959 4437
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19426 4264 19432 4276
rect 19383 4236 19432 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 19978 4264 19984 4276
rect 19939 4236 19984 4264
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20622 4264 20628 4276
rect 20583 4236 20628 4264
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 21910 4264 21916 4276
rect 21871 4236 21916 4264
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22557 4267 22615 4273
rect 22557 4264 22569 4267
rect 22520 4236 22569 4264
rect 22520 4224 22526 4236
rect 22557 4233 22569 4236
rect 22603 4233 22615 4267
rect 22557 4227 22615 4233
rect 22664 4236 24900 4264
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 21266 4196 21272 4208
rect 18104 4168 18276 4196
rect 18104 4156 18110 4168
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2774 4128 2780 4140
rect 2735 4100 2780 4128
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 6546 4088 6552 4100
rect 6604 4128 6610 4140
rect 7098 4128 7104 4140
rect 6604 4100 7104 4128
rect 6604 4088 6610 4100
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7374 4128 7380 4140
rect 7248 4100 7380 4128
rect 7248 4088 7254 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 7837 4091 7895 4097
rect 7852 4060 7880 4091
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17954 4128 17960 4140
rect 17543 4100 17960 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18248 4128 18276 4168
rect 18800 4168 21272 4196
rect 18800 4128 18828 4168
rect 21266 4156 21272 4168
rect 21324 4156 21330 4208
rect 22664 4196 22692 4236
rect 21652 4168 21956 4196
rect 18248 4100 18828 4128
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 19245 4131 19303 4137
rect 19245 4128 19257 4131
rect 18932 4100 19257 4128
rect 18932 4088 18938 4100
rect 19245 4097 19257 4100
rect 19291 4097 19303 4131
rect 19245 4091 19303 4097
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19392 4100 19901 4128
rect 19392 4088 19398 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 19889 4091 19947 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21652 4128 21680 4168
rect 21818 4128 21824 4140
rect 21232 4100 21680 4128
rect 21779 4100 21824 4128
rect 21232 4088 21238 4100
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 21928 4128 21956 4168
rect 22296 4168 22692 4196
rect 23584 4168 24716 4196
rect 22296 4128 22324 4168
rect 21928 4100 22324 4128
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 22428 4100 22477 4128
rect 22428 4088 22434 4100
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 23106 4128 23112 4140
rect 23067 4100 23112 4128
rect 22465 4091 22523 4097
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23584 4128 23612 4168
rect 23750 4128 23756 4140
rect 23216 4100 23612 4128
rect 23711 4100 23756 4128
rect 7852 4032 20208 4060
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7929 3995 7987 4001
rect 7929 3992 7941 3995
rect 6972 3964 7941 3992
rect 6972 3952 6978 3964
rect 7929 3961 7941 3964
rect 7975 3961 7987 3995
rect 7929 3955 7987 3961
rect 10870 3952 10876 4004
rect 10928 3992 10934 4004
rect 17589 3995 17647 4001
rect 10928 3964 12434 3992
rect 10928 3952 10934 3964
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2004 3896 2237 3924
rect 2004 3884 2010 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2832 3896 2881 3924
rect 2832 3884 2838 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 6638 3924 6644 3936
rect 6599 3896 6644 3924
rect 2869 3887 2927 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7282 3924 7288 3936
rect 7243 3896 7288 3924
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 9490 3924 9496 3936
rect 9451 3896 9496 3924
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 11296 3896 11989 3924
rect 11296 3884 11302 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 12406 3924 12434 3964
rect 17589 3961 17601 3995
rect 17635 3992 17647 3995
rect 18966 3992 18972 4004
rect 17635 3964 18972 3992
rect 17635 3961 17647 3964
rect 17589 3955 17647 3961
rect 18966 3952 18972 3964
rect 19024 3952 19030 4004
rect 19058 3952 19064 4004
rect 19116 3992 19122 4004
rect 20180 3992 20208 4032
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 23216 4060 23244 4100
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24581 4131 24639 4137
rect 23900 4100 23945 4128
rect 23900 4088 23906 4100
rect 24581 4097 24593 4131
rect 24627 4097 24639 4131
rect 24688 4128 24716 4168
rect 24872 4128 24900 4236
rect 39482 4224 39488 4276
rect 39540 4264 39546 4276
rect 39945 4267 40003 4273
rect 39945 4264 39957 4267
rect 39540 4236 39957 4264
rect 39540 4224 39546 4236
rect 39945 4233 39957 4236
rect 39991 4233 40003 4267
rect 39945 4227 40003 4233
rect 40972 4236 45232 4264
rect 40972 4196 41000 4236
rect 38626 4168 41000 4196
rect 38626 4140 38654 4168
rect 24688 4100 24808 4128
rect 24872 4100 36584 4128
rect 24581 4091 24639 4097
rect 22336 4032 23244 4060
rect 22336 4020 22342 4032
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 24596 4060 24624 4091
rect 23348 4032 24624 4060
rect 23348 4020 23354 4032
rect 24670 3992 24676 4004
rect 19116 3964 19380 3992
rect 20180 3964 24676 3992
rect 19116 3952 19122 3964
rect 18046 3924 18052 3936
rect 12406 3896 18052 3924
rect 11977 3887 12035 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 19242 3924 19248 3936
rect 18279 3896 19248 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 19352 3924 19380 3964
rect 24670 3952 24676 3964
rect 24728 3952 24734 4004
rect 22002 3924 22008 3936
rect 19352 3896 22008 3924
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 22796 3896 23213 3924
rect 22796 3884 22802 3896
rect 23201 3893 23213 3896
rect 23247 3893 23259 3927
rect 23201 3887 23259 3893
rect 24397 3927 24455 3933
rect 24397 3893 24409 3927
rect 24443 3924 24455 3927
rect 24486 3924 24492 3936
rect 24443 3896 24492 3924
rect 24443 3893 24455 3896
rect 24397 3887 24455 3893
rect 24486 3884 24492 3896
rect 24544 3884 24550 3936
rect 24780 3924 24808 4100
rect 29362 4020 29368 4072
rect 29420 4060 29426 4072
rect 36262 4060 36268 4072
rect 29420 4032 36268 4060
rect 29420 4020 29426 4032
rect 36262 4020 36268 4032
rect 36320 4020 36326 4072
rect 36556 4060 36584 4100
rect 38562 4088 38568 4140
rect 38620 4100 38654 4140
rect 38620 4088 38626 4100
rect 39206 4088 39212 4140
rect 39264 4128 39270 4140
rect 39850 4128 39856 4140
rect 39264 4100 39309 4128
rect 39811 4100 39856 4128
rect 39264 4088 39270 4100
rect 39850 4088 39856 4100
rect 39908 4088 39914 4140
rect 40972 4137 41000 4168
rect 41230 4156 41236 4208
rect 41288 4196 41294 4208
rect 41288 4168 41552 4196
rect 41288 4156 41294 4168
rect 40957 4131 41015 4137
rect 40957 4097 40969 4131
rect 41003 4097 41015 4131
rect 40957 4091 41015 4097
rect 41046 4088 41052 4140
rect 41104 4128 41110 4140
rect 41414 4128 41420 4140
rect 41104 4100 41420 4128
rect 41104 4088 41110 4100
rect 41414 4088 41420 4100
rect 41472 4088 41478 4140
rect 39390 4060 39396 4072
rect 36556 4032 39396 4060
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 41138 4060 41144 4072
rect 41099 4032 41144 4060
rect 41138 4020 41144 4032
rect 41196 4020 41202 4072
rect 41524 4060 41552 4168
rect 42904 4137 42932 4236
rect 43070 4196 43076 4208
rect 43031 4168 43076 4196
rect 43070 4156 43076 4168
rect 43128 4156 43134 4208
rect 45204 4196 45232 4236
rect 45646 4224 45652 4276
rect 45704 4264 45710 4276
rect 45922 4264 45928 4276
rect 45704 4236 45928 4264
rect 45704 4224 45710 4236
rect 45922 4224 45928 4236
rect 45980 4224 45986 4276
rect 46014 4196 46020 4208
rect 45204 4168 46020 4196
rect 42889 4131 42947 4137
rect 42889 4097 42901 4131
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 44729 4131 44787 4137
rect 44729 4097 44741 4131
rect 44775 4128 44787 4131
rect 45002 4128 45008 4140
rect 44775 4100 45008 4128
rect 44775 4097 44787 4100
rect 44729 4091 44787 4097
rect 44744 4060 44772 4091
rect 45002 4088 45008 4100
rect 45060 4088 45066 4140
rect 45204 4137 45232 4168
rect 46014 4156 46020 4168
rect 46072 4156 46078 4208
rect 45189 4131 45247 4137
rect 45189 4097 45201 4131
rect 45235 4097 45247 4131
rect 45189 4091 45247 4097
rect 47857 4131 47915 4137
rect 47857 4097 47869 4131
rect 47903 4128 47915 4131
rect 48314 4128 48320 4140
rect 47903 4100 48320 4128
rect 47903 4097 47915 4100
rect 47857 4091 47915 4097
rect 48314 4088 48320 4100
rect 48372 4088 48378 4140
rect 41524 4032 44772 4060
rect 45373 4063 45431 4069
rect 45373 4029 45385 4063
rect 45419 4060 45431 4063
rect 45830 4060 45836 4072
rect 45419 4032 45836 4060
rect 45419 4029 45431 4032
rect 45373 4023 45431 4029
rect 45830 4020 45836 4032
rect 45888 4020 45894 4072
rect 45922 4020 45928 4072
rect 45980 4060 45986 4072
rect 45980 4032 46025 4060
rect 45980 4020 45986 4032
rect 24854 3952 24860 4004
rect 24912 3992 24918 4004
rect 24912 3964 39988 3992
rect 24912 3952 24918 3964
rect 38378 3924 38384 3936
rect 24780 3896 38384 3924
rect 38378 3884 38384 3896
rect 38436 3884 38442 3936
rect 38470 3884 38476 3936
rect 38528 3924 38534 3936
rect 39301 3927 39359 3933
rect 39301 3924 39313 3927
rect 38528 3896 39313 3924
rect 38528 3884 38534 3896
rect 39301 3893 39313 3896
rect 39347 3893 39359 3927
rect 39960 3924 39988 3964
rect 40034 3952 40040 4004
rect 40092 3992 40098 4004
rect 48041 3995 48099 4001
rect 48041 3992 48053 3995
rect 40092 3964 48053 3992
rect 40092 3952 40098 3964
rect 48041 3961 48053 3964
rect 48087 3961 48099 3995
rect 48041 3955 48099 3961
rect 41046 3924 41052 3936
rect 39960 3896 41052 3924
rect 39301 3887 39359 3893
rect 41046 3884 41052 3896
rect 41104 3884 41110 3936
rect 41322 3924 41328 3936
rect 41283 3896 41328 3924
rect 41322 3884 41328 3896
rect 41380 3884 41386 3936
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 45462 3924 45468 3936
rect 41472 3896 45468 3924
rect 41472 3884 41478 3896
rect 45462 3884 45468 3896
rect 45520 3884 45526 3936
rect 45554 3884 45560 3936
rect 45612 3924 45618 3936
rect 47762 3924 47768 3936
rect 45612 3896 47768 3924
rect 45612 3884 45618 3896
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7156 3692 11836 3720
rect 7156 3680 7162 3692
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 10870 3652 10876 3664
rect 3476 3624 10876 3652
rect 3476 3612 3482 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 11020 3624 11560 3652
rect 11020 3612 11026 3624
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7190 3584 7196 3596
rect 7151 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11532 3593 11560 3624
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3553 11575 3587
rect 11808 3584 11836 3692
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 11940 3692 13860 3720
rect 11940 3680 11946 3692
rect 13832 3652 13860 3692
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 18690 3720 18696 3732
rect 13964 3692 18696 3720
rect 13964 3680 13970 3692
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 19978 3720 19984 3732
rect 19306 3692 19984 3720
rect 18598 3652 18604 3664
rect 13832 3624 18604 3652
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 17129 3587 17187 3593
rect 11808 3556 13860 3584
rect 11517 3547 11575 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2317 3519 2375 3525
rect 2317 3516 2329 3519
rect 1820 3488 2329 3516
rect 1820 3476 1826 3488
rect 2317 3485 2329 3488
rect 2363 3485 2375 3519
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2317 3479 2375 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 7852 3488 9137 3516
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7852 3448 7880 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9950 3516 9956 3528
rect 9911 3488 9956 3516
rect 9125 3479 9183 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13722 3516 13728 3528
rect 13587 3488 13728 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13832 3516 13860 3556
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 19306 3584 19334 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 32122 3720 32128 3732
rect 20220 3692 32128 3720
rect 20220 3680 20226 3692
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 38930 3720 38936 3732
rect 32824 3692 38936 3720
rect 32824 3680 32830 3692
rect 38930 3680 38936 3692
rect 38988 3680 38994 3732
rect 39206 3720 39212 3732
rect 39167 3692 39212 3720
rect 39206 3680 39212 3692
rect 39264 3680 39270 3732
rect 47026 3720 47032 3732
rect 39316 3692 47032 3720
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19484 3624 26280 3652
rect 19484 3612 19490 3624
rect 17175 3556 19334 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 19978 3544 19984 3596
rect 20036 3584 20042 3596
rect 20036 3556 24164 3584
rect 20036 3544 20042 3556
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13832 3488 14105 3516
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 14093 3479 14151 3485
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3516 18107 3519
rect 18414 3516 18420 3528
rect 18095 3488 18420 3516
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 15194 3448 15200 3460
rect 7156 3420 7880 3448
rect 9876 3420 15200 3448
rect 7156 3408 7162 3420
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 9876 3380 9904 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 15562 3448 15568 3460
rect 15519 3420 15568 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 19058 3448 19064 3460
rect 17552 3420 19064 3448
rect 17552 3408 17558 3420
rect 19058 3408 19064 3420
rect 19116 3408 19122 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 20272 3448 20300 3479
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20404 3488 20729 3516
rect 20404 3476 20410 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 21545 3519 21603 3525
rect 21545 3485 21557 3519
rect 21591 3516 21603 3519
rect 21818 3516 21824 3528
rect 21591 3488 21824 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 21818 3476 21824 3488
rect 21876 3476 21882 3528
rect 22738 3516 22744 3528
rect 22699 3488 22744 3516
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 22879 3488 23397 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23532 3488 23577 3516
rect 23532 3476 23538 3488
rect 19392 3420 20300 3448
rect 19392 3408 19398 3420
rect 21910 3408 21916 3460
rect 21968 3448 21974 3460
rect 22097 3451 22155 3457
rect 22097 3448 22109 3451
rect 21968 3420 22109 3448
rect 21968 3408 21974 3420
rect 22097 3417 22109 3420
rect 22143 3417 22155 3451
rect 24136 3448 24164 3556
rect 24578 3544 24584 3596
rect 24636 3584 24642 3596
rect 25501 3587 25559 3593
rect 25501 3584 25513 3587
rect 24636 3556 25513 3584
rect 24636 3544 24642 3556
rect 25501 3553 25513 3556
rect 25547 3553 25559 3587
rect 26252 3584 26280 3624
rect 26326 3612 26332 3664
rect 26384 3652 26390 3664
rect 39316 3652 39344 3692
rect 47026 3680 47032 3692
rect 47084 3680 47090 3732
rect 26384 3624 39344 3652
rect 26384 3612 26390 3624
rect 39390 3612 39396 3664
rect 39448 3652 39454 3664
rect 42518 3652 42524 3664
rect 39448 3624 42524 3652
rect 39448 3612 39454 3624
rect 42518 3612 42524 3624
rect 42576 3612 42582 3664
rect 45646 3612 45652 3664
rect 45704 3652 45710 3664
rect 47578 3652 47584 3664
rect 45704 3624 47584 3652
rect 45704 3612 45710 3624
rect 47578 3612 47584 3624
rect 47636 3612 47642 3664
rect 26786 3584 26792 3596
rect 26252 3556 26648 3584
rect 26747 3556 26792 3584
rect 25501 3547 25559 3553
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 24670 3476 24676 3488
rect 24728 3516 24734 3528
rect 26326 3516 26332 3528
rect 24728 3488 26332 3516
rect 24728 3476 24734 3488
rect 26326 3476 26332 3488
rect 26384 3476 26390 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 26476 3488 26525 3516
rect 26476 3476 26482 3488
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 26620 3516 26648 3556
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 32968 3556 37872 3584
rect 32968 3525 32996 3556
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 26620 3488 32965 3516
rect 26513 3479 26571 3485
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 33042 3476 33048 3528
rect 33100 3516 33106 3528
rect 33100 3488 33145 3516
rect 33100 3476 33106 3488
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 33781 3519 33839 3525
rect 33781 3516 33793 3519
rect 33284 3488 33793 3516
rect 33284 3476 33290 3488
rect 33781 3485 33793 3488
rect 33827 3485 33839 3519
rect 33781 3479 33839 3485
rect 35897 3519 35955 3525
rect 35897 3485 35909 3519
rect 35943 3485 35955 3519
rect 37844 3518 37872 3556
rect 38010 3544 38016 3596
rect 38068 3584 38074 3596
rect 38068 3556 39620 3584
rect 38068 3544 38074 3556
rect 37844 3490 37964 3518
rect 38470 3516 38476 3528
rect 35897 3479 35955 3485
rect 32766 3448 32772 3460
rect 24136 3420 32772 3448
rect 22097 3411 22155 3417
rect 32766 3408 32772 3420
rect 32824 3408 32830 3460
rect 10042 3380 10048 3392
rect 1627 3352 9904 3380
rect 10003 3352 10048 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 13814 3380 13820 3392
rect 11664 3352 13820 3380
rect 11664 3340 11670 3352
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13964 3352 14197 3380
rect 13964 3340 13970 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3380 18199 3383
rect 18506 3380 18512 3392
rect 18187 3352 18512 3380
rect 18187 3349 18199 3352
rect 18141 3343 18199 3349
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19484 3352 19533 3380
rect 19484 3340 19490 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19521 3343 19579 3349
rect 20809 3383 20867 3389
rect 20809 3349 20821 3383
rect 20855 3380 20867 3383
rect 22002 3380 22008 3392
rect 20855 3352 22008 3380
rect 20855 3349 20867 3352
rect 20809 3343 20867 3349
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 22186 3380 22192 3392
rect 22147 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 27522 3380 27528 3392
rect 24912 3352 27528 3380
rect 24912 3340 24918 3352
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 30926 3340 30932 3392
rect 30984 3380 30990 3392
rect 32214 3380 32220 3392
rect 30984 3352 32220 3380
rect 30984 3340 30990 3352
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 35912 3380 35940 3479
rect 36081 3451 36139 3457
rect 36081 3417 36093 3451
rect 36127 3448 36139 3451
rect 36170 3448 36176 3460
rect 36127 3420 36176 3448
rect 36127 3417 36139 3420
rect 36081 3411 36139 3417
rect 36170 3408 36176 3420
rect 36228 3408 36234 3460
rect 36262 3408 36268 3460
rect 36320 3448 36326 3460
rect 37737 3451 37795 3457
rect 37737 3448 37749 3451
rect 36320 3420 37749 3448
rect 36320 3408 36326 3420
rect 37737 3417 37749 3420
rect 37783 3448 37795 3451
rect 37826 3448 37832 3460
rect 37783 3420 37832 3448
rect 37783 3417 37795 3420
rect 37737 3411 37795 3417
rect 37826 3408 37832 3420
rect 37884 3408 37890 3460
rect 37936 3448 37964 3490
rect 38431 3488 38476 3516
rect 38470 3476 38476 3488
rect 38528 3476 38534 3528
rect 39117 3519 39175 3525
rect 39117 3485 39129 3519
rect 39163 3516 39175 3519
rect 39482 3516 39488 3528
rect 39163 3488 39488 3516
rect 39163 3485 39175 3488
rect 39117 3479 39175 3485
rect 39482 3476 39488 3488
rect 39540 3476 39546 3528
rect 39592 3510 39620 3556
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 40037 3587 40095 3593
rect 40037 3584 40049 3587
rect 39816 3556 40049 3584
rect 39816 3544 39822 3556
rect 40037 3553 40049 3556
rect 40083 3553 40095 3587
rect 41322 3584 41328 3596
rect 41283 3556 41328 3584
rect 40037 3547 40095 3553
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 44453 3587 44511 3593
rect 44453 3553 44465 3587
rect 44499 3584 44511 3587
rect 45462 3584 45468 3596
rect 44499 3556 45468 3584
rect 44499 3553 44511 3556
rect 44453 3547 44511 3553
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 39942 3516 39948 3528
rect 39684 3510 39948 3516
rect 39592 3488 39948 3510
rect 39592 3482 39712 3488
rect 39942 3476 39948 3488
rect 40000 3476 40006 3528
rect 40310 3516 40316 3528
rect 40271 3488 40316 3516
rect 40310 3476 40316 3488
rect 40368 3476 40374 3528
rect 43625 3519 43683 3525
rect 43625 3516 43637 3519
rect 42720 3488 43637 3516
rect 37936 3420 39620 3448
rect 39592 3419 39620 3420
rect 38470 3380 38476 3392
rect 32732 3352 38476 3380
rect 32732 3340 32738 3352
rect 38470 3340 38476 3352
rect 38528 3340 38534 3392
rect 38565 3383 38623 3389
rect 38565 3349 38577 3383
rect 38611 3380 38623 3383
rect 39482 3380 39488 3392
rect 38611 3352 39488 3380
rect 38611 3349 38623 3352
rect 38565 3343 38623 3349
rect 39482 3340 39488 3352
rect 39540 3340 39546 3392
rect 39592 3391 39712 3419
rect 41138 3408 41144 3460
rect 41196 3448 41202 3460
rect 41322 3448 41328 3460
rect 41196 3420 41328 3448
rect 41196 3408 41202 3420
rect 41322 3408 41328 3420
rect 41380 3448 41386 3460
rect 41509 3451 41567 3457
rect 41509 3448 41521 3451
rect 41380 3420 41521 3448
rect 41380 3408 41386 3420
rect 41509 3417 41521 3420
rect 41555 3417 41567 3451
rect 42720 3448 42748 3488
rect 43625 3485 43637 3488
rect 43671 3485 43683 3519
rect 43625 3479 43683 3485
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3516 45063 3519
rect 45370 3516 45376 3528
rect 45051 3488 45376 3516
rect 45051 3485 45063 3488
rect 45005 3479 45063 3485
rect 45370 3476 45376 3488
rect 45428 3476 45434 3528
rect 45646 3476 45652 3528
rect 45704 3516 45710 3528
rect 46290 3516 46296 3528
rect 45704 3488 45747 3516
rect 46251 3488 46296 3516
rect 45704 3476 45710 3488
rect 46290 3476 46296 3488
rect 46348 3476 46354 3528
rect 41509 3411 41567 3417
rect 42352 3420 42748 3448
rect 42352 3392 42380 3420
rect 42978 3408 42984 3460
rect 43036 3448 43042 3460
rect 43165 3451 43223 3457
rect 43165 3448 43177 3451
rect 43036 3420 43177 3448
rect 43036 3408 43042 3420
rect 43165 3417 43177 3420
rect 43211 3448 43223 3451
rect 45554 3448 45560 3460
rect 43211 3420 45560 3448
rect 43211 3417 43223 3420
rect 43165 3411 43223 3417
rect 45554 3408 45560 3420
rect 45612 3408 45618 3460
rect 45741 3451 45799 3457
rect 45741 3417 45753 3451
rect 45787 3448 45799 3451
rect 46477 3451 46535 3457
rect 46477 3448 46489 3451
rect 45787 3420 46489 3448
rect 45787 3417 45799 3420
rect 45741 3411 45799 3417
rect 46477 3417 46489 3420
rect 46523 3417 46535 3451
rect 46477 3411 46535 3417
rect 48133 3451 48191 3457
rect 48133 3417 48145 3451
rect 48179 3448 48191 3451
rect 48958 3448 48964 3460
rect 48179 3420 48964 3448
rect 48179 3417 48191 3420
rect 48133 3411 48191 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 39684 3380 39712 3391
rect 42334 3380 42340 3392
rect 39684 3352 42340 3380
rect 42334 3340 42340 3352
rect 42392 3340 42398 3392
rect 42610 3340 42616 3392
rect 42668 3380 42674 3392
rect 43717 3383 43775 3389
rect 43717 3380 43729 3383
rect 42668 3352 43729 3380
rect 42668 3340 42674 3352
rect 43717 3349 43729 3352
rect 43763 3349 43775 3383
rect 43717 3343 43775 3349
rect 45097 3383 45155 3389
rect 45097 3349 45109 3383
rect 45143 3380 45155 3383
rect 45370 3380 45376 3392
rect 45143 3352 45376 3380
rect 45143 3349 45155 3352
rect 45097 3343 45155 3349
rect 45370 3340 45376 3352
rect 45428 3340 45434 3392
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 46290 3380 46296 3392
rect 45520 3352 46296 3380
rect 45520 3340 45526 3352
rect 46290 3340 46296 3352
rect 46348 3340 46354 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 17218 3176 17224 3188
rect 9692 3148 17224 3176
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 7282 3108 7288 3120
rect 7243 3080 7288 3108
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 9692 3117 9720 3148
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 18230 3176 18236 3188
rect 17368 3148 18236 3176
rect 17368 3136 17374 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 32766 3176 32772 3188
rect 18656 3148 24900 3176
rect 18656 3136 18662 3148
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3077 9735 3111
rect 13906 3108 13912 3120
rect 13867 3080 13912 3108
rect 9677 3071 9735 3077
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 24762 3108 24768 3120
rect 15252 3080 23244 3108
rect 24723 3080 24768 3108
rect 15252 3068 15258 3080
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6512 3012 6653 3040
rect 6512 3000 6518 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 7098 3040 7104 3052
rect 7059 3012 7104 3040
rect 6641 3003 6699 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 8536 3012 9505 3040
rect 8536 3000 8542 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11112 3012 11713 3040
rect 11112 3000 11118 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 13722 3040 13728 3052
rect 13683 3012 13728 3040
rect 11701 3003 11759 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17497 3003 17555 3009
rect 17880 3012 18337 3040
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 716 2944 2237 2972
rect 716 2932 722 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 2225 2935 2283 2941
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 15252 2944 17417 2972
rect 15252 2932 15258 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 15286 2904 15292 2916
rect 7064 2876 15292 2904
rect 7064 2864 7070 2876
rect 15286 2864 15292 2876
rect 15344 2864 15350 2916
rect 17310 2904 17316 2916
rect 17144 2876 17316 2904
rect 7374 2796 7380 2848
rect 7432 2836 7438 2848
rect 17144 2836 17172 2876
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 17512 2904 17540 3003
rect 17880 2981 17908 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 18325 3003 18383 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 21818 3040 21824 3052
rect 21779 3012 21824 3040
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2941 17923 2975
rect 19518 2972 19524 2984
rect 19479 2944 19524 2972
rect 17865 2935 17923 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 22002 2972 22008 2984
rect 21963 2944 22008 2972
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 23216 2972 23244 3080
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 24872 3108 24900 3148
rect 28276 3148 32772 3176
rect 28276 3117 28304 3148
rect 32766 3136 32772 3148
rect 32824 3136 32830 3188
rect 36170 3176 36176 3188
rect 32876 3148 36032 3176
rect 36131 3148 36176 3176
rect 28261 3111 28319 3117
rect 24872 3080 26234 3108
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 25130 2972 25136 2984
rect 23216 2944 24992 2972
rect 25091 2944 25136 2972
rect 24854 2904 24860 2916
rect 17512 2876 24860 2904
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 24964 2904 24992 2944
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 25222 2904 25228 2916
rect 24964 2876 25228 2904
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 26206 2904 26234 3080
rect 28261 3077 28273 3111
rect 28307 3077 28319 3111
rect 32876 3108 32904 3148
rect 33042 3108 33048 3120
rect 28261 3071 28319 3077
rect 31726 3080 32904 3108
rect 33003 3080 33048 3108
rect 28074 3040 28080 3052
rect 28035 3012 28080 3040
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 27522 2932 27528 2984
rect 27580 2972 27586 2984
rect 29917 2975 29975 2981
rect 29917 2972 29929 2975
rect 27580 2944 29929 2972
rect 27580 2932 27586 2944
rect 29917 2941 29929 2944
rect 29963 2972 29975 2975
rect 31726 2972 31754 3080
rect 33042 3068 33048 3080
rect 33100 3068 33106 3120
rect 36004 3108 36032 3148
rect 36170 3136 36176 3148
rect 36228 3136 36234 3188
rect 39117 3179 39175 3185
rect 39117 3145 39129 3179
rect 39163 3176 39175 3179
rect 39850 3176 39856 3188
rect 39163 3148 39856 3176
rect 39163 3145 39175 3148
rect 39117 3139 39175 3145
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 39942 3136 39948 3188
rect 40000 3176 40006 3188
rect 46382 3176 46388 3188
rect 40000 3148 46388 3176
rect 40000 3136 40006 3148
rect 46382 3136 46388 3148
rect 46440 3136 46446 3188
rect 39761 3111 39819 3117
rect 39761 3108 39773 3111
rect 36004 3080 38608 3108
rect 29963 2944 31754 2972
rect 32508 3012 32812 3040
rect 29963 2941 29975 2944
rect 29917 2935 29975 2941
rect 32508 2904 32536 3012
rect 26206 2876 32536 2904
rect 32784 2904 32812 3012
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 36136 3012 36369 3040
rect 36136 3000 36142 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 38470 3040 38476 3052
rect 38431 3012 38476 3040
rect 36357 3003 36415 3009
rect 38470 3000 38476 3012
rect 38528 3000 38534 3052
rect 32861 2975 32919 2981
rect 32861 2941 32873 2975
rect 32907 2972 32919 2975
rect 33226 2972 33232 2984
rect 32907 2944 33232 2972
rect 32907 2941 32919 2944
rect 32861 2935 32919 2941
rect 33226 2932 33232 2944
rect 33284 2932 33290 2984
rect 33502 2972 33508 2984
rect 33463 2944 33508 2972
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 38580 2972 38608 3080
rect 38672 3080 39773 3108
rect 38672 3049 38700 3080
rect 39761 3077 39773 3080
rect 39807 3108 39819 3111
rect 40310 3108 40316 3120
rect 39807 3080 40316 3108
rect 39807 3077 39819 3080
rect 39761 3071 39819 3077
rect 40310 3068 40316 3080
rect 40368 3068 40374 3120
rect 42610 3108 42616 3120
rect 42571 3080 42616 3108
rect 42610 3068 42616 3080
rect 42668 3068 42674 3120
rect 45370 3108 45376 3120
rect 45331 3080 45376 3108
rect 45370 3068 45376 3080
rect 45428 3068 45434 3120
rect 47762 3108 47768 3120
rect 47723 3080 47768 3108
rect 47762 3068 47768 3080
rect 47820 3068 47826 3120
rect 38657 3043 38715 3049
rect 38657 3009 38669 3043
rect 38703 3009 38715 3043
rect 38657 3003 38715 3009
rect 39482 3000 39488 3052
rect 39540 3040 39546 3052
rect 39577 3043 39635 3049
rect 39577 3040 39589 3043
rect 39540 3012 39589 3040
rect 39540 3000 39546 3012
rect 39577 3009 39589 3012
rect 39623 3009 39635 3043
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 39577 3003 39635 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 40037 2975 40095 2981
rect 40037 2972 40049 2975
rect 38580 2944 40049 2972
rect 40037 2941 40049 2944
rect 40083 2972 40095 2975
rect 42978 2972 42984 2984
rect 40083 2944 42984 2972
rect 40083 2941 40095 2944
rect 40037 2935 40095 2941
rect 42978 2932 42984 2944
rect 43036 2932 43042 2984
rect 43162 2972 43168 2984
rect 43123 2944 43168 2972
rect 43162 2932 43168 2944
rect 43220 2932 43226 2984
rect 47029 2975 47087 2981
rect 47029 2941 47041 2975
rect 47075 2972 47087 2975
rect 47670 2972 47676 2984
rect 47075 2944 47676 2972
rect 47075 2941 47087 2944
rect 47029 2935 47087 2941
rect 47670 2932 47676 2944
rect 47728 2932 47734 2984
rect 43254 2904 43260 2916
rect 32784 2876 43260 2904
rect 43254 2864 43260 2876
rect 43312 2864 43318 2916
rect 7432 2808 17172 2836
rect 7432 2796 7438 2808
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 23750 2836 23756 2848
rect 17276 2808 23756 2836
rect 17276 2796 17282 2808
rect 23750 2796 23756 2808
rect 23808 2796 23814 2848
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 32674 2836 32680 2848
rect 23900 2808 32680 2836
rect 23900 2796 23906 2808
rect 32674 2796 32680 2808
rect 32732 2796 32738 2848
rect 32766 2796 32772 2848
rect 32824 2836 32830 2848
rect 40034 2836 40040 2848
rect 32824 2808 40040 2836
rect 32824 2796 32830 2808
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 47857 2839 47915 2845
rect 47857 2836 47869 2839
rect 40184 2808 47869 2836
rect 40184 2796 40190 2808
rect 47857 2805 47869 2808
rect 47903 2805 47915 2839
rect 47857 2799 47915 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 3292 2604 17264 2632
rect 3292 2592 3298 2604
rect 2958 2564 2964 2576
rect 1412 2536 2964 2564
rect 1412 2505 1440 2536
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 5276 2536 8984 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 2866 2496 2872 2508
rect 2827 2468 2872 2496
rect 1397 2459 1455 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5276 2505 5304 2536
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6052 2468 6561 2496
rect 6052 2456 6058 2468
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6914 2496 6920 2508
rect 6779 2468 6920 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7064 2468 7109 2496
rect 7064 2456 7070 2468
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5166 2428 5172 2440
rect 5031 2400 5172 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 2774 2360 2780 2372
rect 1627 2332 2780 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 4172 2292 4200 2323
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 7006 2360 7012 2372
rect 6512 2332 7012 2360
rect 6512 2320 6518 2332
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 4430 2292 4436 2304
rect 2648 2264 4200 2292
rect 4391 2264 4436 2292
rect 2648 2252 2654 2264
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 8956 2292 8984 2536
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9088 2536 9720 2564
rect 9088 2524 9094 2536
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2496 9183 2499
rect 9490 2496 9496 2508
rect 9171 2468 9496 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9692 2505 9720 2536
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2465 9735 2499
rect 15562 2496 15568 2508
rect 15523 2468 15568 2496
rect 9677 2459 9735 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 9309 2363 9367 2369
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 10042 2360 10048 2372
rect 9355 2332 10048 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16172 2332 17141 2360
rect 16172 2320 16178 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17236 2360 17264 2604
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 18196 2604 18613 2632
rect 18196 2592 18202 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 18601 2595 18659 2601
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 20070 2632 20076 2644
rect 19383 2604 20076 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 23017 2635 23075 2641
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 23842 2632 23848 2644
rect 23063 2604 23848 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 26145 2635 26203 2641
rect 26145 2632 26157 2635
rect 23992 2604 26157 2632
rect 23992 2592 23998 2604
rect 26145 2601 26157 2604
rect 26191 2601 26203 2635
rect 26145 2595 26203 2601
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 35759 2635 35817 2641
rect 35759 2632 35771 2635
rect 26936 2604 35771 2632
rect 26936 2592 26942 2604
rect 35759 2601 35771 2604
rect 35805 2601 35817 2635
rect 47857 2635 47915 2641
rect 47857 2632 47869 2635
rect 35759 2595 35817 2601
rect 35866 2604 47869 2632
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2564 17371 2567
rect 25222 2564 25228 2576
rect 17359 2536 25228 2564
rect 17359 2533 17371 2536
rect 17313 2527 17371 2533
rect 25222 2524 25228 2536
rect 25280 2524 25286 2576
rect 25314 2524 25320 2576
rect 25372 2564 25378 2576
rect 35866 2564 35894 2604
rect 47857 2601 47869 2604
rect 47903 2601 47915 2635
rect 47857 2595 47915 2601
rect 40494 2564 40500 2576
rect 25372 2536 35894 2564
rect 40455 2536 40500 2564
rect 25372 2524 25378 2536
rect 40494 2524 40500 2536
rect 40552 2524 40558 2576
rect 43073 2567 43131 2573
rect 43073 2533 43085 2567
rect 43119 2564 43131 2567
rect 45738 2564 45744 2576
rect 43119 2536 45744 2564
rect 43119 2533 43131 2536
rect 43073 2527 43131 2533
rect 45738 2524 45744 2536
rect 45796 2524 45802 2576
rect 20717 2499 20775 2505
rect 20717 2465 20729 2499
rect 20763 2496 20775 2499
rect 24302 2496 24308 2508
rect 20763 2468 24308 2496
rect 20763 2465 20775 2468
rect 20717 2459 20775 2465
rect 24302 2456 24308 2468
rect 24360 2456 24366 2508
rect 24486 2496 24492 2508
rect 24447 2468 24492 2496
rect 24486 2456 24492 2468
rect 24544 2456 24550 2508
rect 25498 2496 25504 2508
rect 25459 2468 25504 2496
rect 25498 2456 25504 2468
rect 25556 2456 25562 2508
rect 28442 2496 28448 2508
rect 28403 2468 28448 2496
rect 28442 2456 28448 2468
rect 28500 2456 28506 2508
rect 30006 2496 30012 2508
rect 29967 2468 30012 2496
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 32030 2456 32036 2508
rect 32088 2496 32094 2508
rect 38381 2499 38439 2505
rect 38381 2496 38393 2499
rect 32088 2468 38393 2496
rect 32088 2456 32094 2468
rect 38381 2465 38393 2468
rect 38427 2465 38439 2499
rect 41322 2496 41328 2508
rect 41283 2468 41328 2496
rect 38381 2459 38439 2465
rect 41322 2456 41328 2468
rect 41380 2456 41386 2508
rect 43625 2499 43683 2505
rect 43625 2465 43637 2499
rect 43671 2496 43683 2499
rect 46014 2496 46020 2508
rect 43671 2468 46020 2496
rect 43671 2465 43683 2468
rect 43625 2459 43683 2465
rect 46014 2456 46020 2468
rect 46072 2456 46078 2508
rect 46201 2499 46259 2505
rect 46201 2465 46213 2499
rect 46247 2496 46259 2499
rect 47026 2496 47032 2508
rect 46247 2468 47032 2496
rect 46247 2465 46259 2468
rect 46201 2459 46259 2465
rect 47026 2456 47032 2468
rect 47084 2456 47090 2508
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 19242 2428 19248 2440
rect 19203 2400 19248 2428
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2428 20499 2431
rect 20622 2428 20628 2440
rect 20487 2400 20628 2428
rect 20487 2397 20499 2400
rect 20441 2391 20499 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 22186 2428 22192 2440
rect 22147 2400 22192 2428
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23198 2428 23204 2440
rect 23155 2400 23204 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 26878 2428 26884 2440
rect 25976 2400 26884 2428
rect 20990 2360 20996 2372
rect 17236 2332 20996 2360
rect 17129 2323 17187 2329
rect 20990 2320 20996 2332
rect 21048 2320 21054 2372
rect 24581 2363 24639 2369
rect 24581 2329 24593 2363
rect 24627 2360 24639 2363
rect 25976 2360 26004 2400
rect 26878 2388 26884 2400
rect 26936 2388 26942 2440
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28350 2428 28356 2440
rect 28215 2400 28356 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 35434 2388 35440 2440
rect 35492 2428 35498 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35492 2400 35541 2428
rect 35492 2388 35498 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41230 2428 41236 2440
rect 41095 2400 41236 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 45462 2428 45468 2440
rect 45423 2400 45468 2428
rect 43901 2391 43959 2397
rect 24627 2332 26004 2360
rect 26053 2363 26111 2369
rect 24627 2329 24639 2332
rect 24581 2323 24639 2329
rect 26053 2329 26065 2363
rect 26099 2329 26111 2363
rect 26053 2323 26111 2329
rect 15194 2292 15200 2304
rect 8956 2264 15200 2292
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 26068 2292 26096 2323
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 27120 2332 27445 2360
rect 27120 2320 27126 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 27617 2363 27675 2369
rect 27617 2329 27629 2363
rect 27663 2360 27675 2363
rect 27663 2332 35894 2360
rect 27663 2329 27675 2332
rect 27617 2323 27675 2329
rect 24544 2264 26096 2292
rect 35866 2292 35894 2332
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 38197 2363 38255 2369
rect 38197 2360 38209 2363
rect 38068 2332 38209 2360
rect 38068 2320 38074 2332
rect 38197 2329 38209 2332
rect 38243 2329 38255 2363
rect 38197 2323 38255 2329
rect 39298 2320 39304 2372
rect 39356 2360 39362 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39356 2332 40325 2360
rect 39356 2320 39362 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 40644 2332 42901 2360
rect 40644 2320 40650 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 43916 2360 43944 2391
rect 45462 2388 45468 2400
rect 45520 2388 45526 2440
rect 45830 2388 45836 2440
rect 45888 2428 45894 2440
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 45888 2400 46489 2428
rect 45888 2388 45894 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 46477 2391 46535 2397
rect 46198 2360 46204 2372
rect 43916 2332 46204 2360
rect 42889 2323 42947 2329
rect 46198 2320 46204 2332
rect 46256 2320 46262 2372
rect 46382 2320 46388 2372
rect 46440 2360 46446 2372
rect 47765 2363 47823 2369
rect 47765 2360 47777 2363
rect 46440 2332 47777 2360
rect 46440 2320 46446 2332
rect 47765 2329 47777 2332
rect 47811 2329 47823 2363
rect 47765 2323 47823 2329
rect 36354 2292 36360 2304
rect 35866 2264 36360 2292
rect 24544 2252 24550 2264
rect 36354 2252 36360 2264
rect 36412 2252 36418 2304
rect 39022 2252 39028 2304
rect 39080 2292 39086 2304
rect 45649 2295 45707 2301
rect 45649 2292 45661 2295
rect 39080 2264 45661 2292
rect 39080 2252 39086 2264
rect 45649 2261 45661 2264
rect 45695 2261 45707 2295
rect 45649 2255 45707 2261
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 25222 2048 25228 2100
rect 25280 2088 25286 2100
rect 29270 2088 29276 2100
rect 25280 2060 29276 2088
rect 25280 2048 25286 2060
rect 29270 2048 29276 2060
rect 29328 2048 29334 2100
rect 4430 1980 4436 2032
rect 4488 2020 4494 2032
rect 29546 2020 29552 2032
rect 4488 1992 29552 2020
rect 4488 1980 4494 1992
rect 29546 1980 29552 1992
rect 29604 1980 29610 2032
<< via1 >>
rect 15292 47404 15344 47456
rect 16488 47404 16540 47456
rect 40040 47404 40092 47456
rect 41236 47404 41288 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 12808 47132 12860 47184
rect 19432 47175 19484 47184
rect 19432 47141 19441 47175
rect 19441 47141 19475 47175
rect 19475 47141 19484 47175
rect 19432 47132 19484 47141
rect 29092 47132 29144 47184
rect 19984 47064 20036 47116
rect 30748 47107 30800 47116
rect 30748 47073 30757 47107
rect 30757 47073 30791 47107
rect 30791 47073 30800 47107
rect 30748 47064 30800 47073
rect 43168 47107 43220 47116
rect 43168 47073 43177 47107
rect 43177 47073 43211 47107
rect 43211 47073 43220 47107
rect 43168 47064 43220 47073
rect 48320 47064 48372 47116
rect 1952 47039 2004 47048
rect 1952 47005 1961 47039
rect 1961 47005 1995 47039
rect 1995 47005 2004 47039
rect 1952 46996 2004 47005
rect 2596 46996 2648 47048
rect 3240 46996 3292 47048
rect 4712 47039 4764 47048
rect 4712 47005 4721 47039
rect 4721 47005 4755 47039
rect 4755 47005 4764 47039
rect 4712 46996 4764 47005
rect 5816 46996 5868 47048
rect 7104 46996 7156 47048
rect 9036 46996 9088 47048
rect 11612 47039 11664 47048
rect 11612 47005 11621 47039
rect 11621 47005 11655 47039
rect 11655 47005 11664 47039
rect 11612 46996 11664 47005
rect 12256 47039 12308 47048
rect 12256 47005 12265 47039
rect 12265 47005 12299 47039
rect 12299 47005 12308 47039
rect 12256 46996 12308 47005
rect 12900 46996 12952 47048
rect 13820 46996 13872 47048
rect 18696 46996 18748 47048
rect 22744 46996 22796 47048
rect 24860 47039 24912 47048
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 28356 46996 28408 47048
rect 29644 46996 29696 47048
rect 31116 46996 31168 47048
rect 38108 46996 38160 47048
rect 42616 47039 42668 47048
rect 42616 47005 42625 47039
rect 42625 47005 42659 47039
rect 42659 47005 42668 47039
rect 42616 46996 42668 47005
rect 44456 46996 44508 47048
rect 47676 46996 47728 47048
rect 4068 46971 4120 46980
rect 4068 46937 4077 46971
rect 4077 46937 4111 46971
rect 4111 46937 4120 46971
rect 4068 46928 4120 46937
rect 4988 46971 5040 46980
rect 4988 46937 4997 46971
rect 4997 46937 5031 46971
rect 5031 46937 5040 46971
rect 4988 46928 5040 46937
rect 7840 46928 7892 46980
rect 11704 46928 11756 46980
rect 13360 46928 13412 46980
rect 14648 46928 14700 46980
rect 2136 46903 2188 46912
rect 2136 46869 2145 46903
rect 2145 46869 2179 46903
rect 2179 46869 2188 46903
rect 2136 46860 2188 46869
rect 2872 46903 2924 46912
rect 2872 46869 2881 46903
rect 2881 46869 2915 46903
rect 2915 46869 2924 46903
rect 2872 46860 2924 46869
rect 6920 46903 6972 46912
rect 6920 46869 6929 46903
rect 6929 46869 6963 46903
rect 6963 46869 6972 46903
rect 9312 46903 9364 46912
rect 6920 46860 6972 46869
rect 9312 46869 9321 46903
rect 9321 46869 9355 46903
rect 9355 46869 9364 46903
rect 9312 46860 9364 46869
rect 16120 46860 16172 46912
rect 17592 46928 17644 46980
rect 28172 46860 28224 46912
rect 39304 46860 39356 46912
rect 40408 46928 40460 46980
rect 43168 46928 43220 46980
rect 45376 46971 45428 46980
rect 45376 46937 45385 46971
rect 45385 46937 45419 46971
rect 45419 46937 45428 46971
rect 45376 46928 45428 46937
rect 47952 46903 48004 46912
rect 47952 46869 47961 46903
rect 47961 46869 47995 46903
rect 47995 46869 48004 46903
rect 47952 46860 48004 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2872 46588 2924 46640
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 24860 46588 24912 46640
rect 28172 46563 28224 46572
rect 28172 46529 28181 46563
rect 28181 46529 28215 46563
rect 28215 46529 28224 46563
rect 28172 46520 28224 46529
rect 38108 46563 38160 46572
rect 38108 46529 38117 46563
rect 38117 46529 38151 46563
rect 38151 46529 38160 46563
rect 38108 46520 38160 46529
rect 47860 46563 47912 46572
rect 47860 46529 47869 46563
rect 47869 46529 47903 46563
rect 47903 46529 47912 46563
rect 47860 46520 47912 46529
rect 3976 46495 4028 46504
rect 3976 46461 3985 46495
rect 3985 46461 4019 46495
rect 4019 46461 4028 46495
rect 3976 46452 4028 46461
rect 5080 46452 5132 46504
rect 3884 46384 3936 46436
rect 12164 46452 12216 46504
rect 1676 46316 1728 46368
rect 10968 46316 11020 46368
rect 13544 46452 13596 46504
rect 14188 46452 14240 46504
rect 14280 46495 14332 46504
rect 14280 46461 14289 46495
rect 14289 46461 14323 46495
rect 14323 46461 14332 46495
rect 19248 46495 19300 46504
rect 14280 46452 14332 46461
rect 19248 46461 19257 46495
rect 19257 46461 19291 46495
rect 19291 46461 19300 46495
rect 19248 46452 19300 46461
rect 20628 46495 20680 46504
rect 18604 46384 18656 46436
rect 20628 46461 20637 46495
rect 20637 46461 20671 46495
rect 20671 46461 20680 46495
rect 20628 46452 20680 46461
rect 24768 46495 24820 46504
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 25136 46495 25188 46504
rect 25136 46461 25145 46495
rect 25145 46461 25179 46495
rect 25179 46461 25188 46495
rect 25136 46452 25188 46461
rect 29368 46495 29420 46504
rect 29368 46461 29377 46495
rect 29377 46461 29411 46495
rect 29411 46461 29420 46495
rect 29368 46452 29420 46461
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 38292 46495 38344 46504
rect 32220 46384 32272 46436
rect 38292 46461 38301 46495
rect 38301 46461 38335 46495
rect 38335 46461 38344 46495
rect 38292 46452 38344 46461
rect 38660 46495 38712 46504
rect 38660 46461 38669 46495
rect 38669 46461 38703 46495
rect 38703 46461 38712 46495
rect 38660 46452 38712 46461
rect 42616 46495 42668 46504
rect 42616 46461 42625 46495
rect 42625 46461 42659 46495
rect 42659 46461 42668 46495
rect 42616 46452 42668 46461
rect 42524 46384 42576 46436
rect 46664 46452 46716 46504
rect 46848 46495 46900 46504
rect 46848 46461 46857 46495
rect 46857 46461 46891 46495
rect 46891 46461 46900 46495
rect 46848 46452 46900 46461
rect 47768 46384 47820 46436
rect 20720 46316 20772 46368
rect 41236 46359 41288 46368
rect 41236 46325 41245 46359
rect 41245 46325 41279 46359
rect 41279 46325 41288 46359
rect 41236 46316 41288 46325
rect 48044 46359 48096 46368
rect 48044 46325 48053 46359
rect 48053 46325 48087 46359
rect 48087 46325 48096 46359
rect 48044 46316 48096 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3976 46112 4028 46164
rect 5080 46155 5132 46164
rect 5080 46121 5089 46155
rect 5089 46121 5123 46155
rect 5123 46121 5132 46155
rect 5080 46112 5132 46121
rect 12164 46155 12216 46164
rect 12164 46121 12173 46155
rect 12173 46121 12207 46155
rect 12207 46121 12216 46155
rect 12164 46112 12216 46121
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14188 46155 14240 46164
rect 14188 46121 14197 46155
rect 14197 46121 14231 46155
rect 14231 46121 14240 46155
rect 14188 46112 14240 46121
rect 18604 46155 18656 46164
rect 18604 46121 18613 46155
rect 18613 46121 18647 46155
rect 18647 46121 18656 46155
rect 18604 46112 18656 46121
rect 19248 46112 19300 46164
rect 24768 46112 24820 46164
rect 32312 46112 32364 46164
rect 38292 46155 38344 46164
rect 38292 46121 38301 46155
rect 38301 46121 38335 46155
rect 38335 46121 38344 46155
rect 38292 46112 38344 46121
rect 20720 46019 20772 46028
rect 1768 45908 1820 45960
rect 11612 45908 11664 45960
rect 14096 45951 14148 45960
rect 14096 45917 14105 45951
rect 14105 45917 14139 45951
rect 14139 45917 14148 45951
rect 18512 45951 18564 45960
rect 14096 45908 14148 45917
rect 18512 45917 18521 45951
rect 18521 45917 18555 45951
rect 18555 45917 18564 45951
rect 18512 45908 18564 45917
rect 20720 45985 20729 46019
rect 20729 45985 20763 46019
rect 20763 45985 20772 46019
rect 20720 45976 20772 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 25504 45976 25556 46028
rect 25780 46019 25832 46028
rect 25780 45985 25789 46019
rect 25789 45985 25823 46019
rect 25823 45985 25832 46019
rect 25780 45976 25832 45985
rect 24584 45951 24636 45960
rect 24584 45917 24593 45951
rect 24593 45917 24627 45951
rect 24627 45917 24636 45951
rect 24584 45908 24636 45917
rect 31760 45951 31812 45960
rect 31760 45917 31769 45951
rect 31769 45917 31803 45951
rect 31803 45917 31812 45951
rect 45008 46044 45060 46096
rect 41236 46019 41288 46028
rect 41236 45985 41245 46019
rect 41245 45985 41279 46019
rect 41279 45985 41288 46019
rect 41236 45976 41288 45985
rect 41880 46019 41932 46028
rect 41880 45985 41889 46019
rect 41889 45985 41923 46019
rect 41923 45985 41932 46019
rect 41880 45976 41932 45985
rect 47032 46019 47084 46028
rect 47032 45985 47041 46019
rect 47041 45985 47075 46019
rect 47075 45985 47084 46019
rect 47032 45976 47084 45985
rect 31760 45908 31812 45917
rect 20720 45840 20772 45892
rect 20904 45883 20956 45892
rect 20904 45849 20913 45883
rect 20913 45849 20947 45883
rect 20947 45849 20956 45883
rect 20904 45840 20956 45849
rect 25412 45883 25464 45892
rect 25412 45849 25421 45883
rect 25421 45849 25455 45883
rect 25455 45849 25464 45883
rect 25412 45840 25464 45849
rect 43812 45908 43864 45960
rect 45744 45908 45796 45960
rect 45836 45908 45888 45960
rect 41420 45883 41472 45892
rect 41420 45849 41429 45883
rect 41429 45849 41463 45883
rect 41463 45849 41472 45883
rect 41420 45840 41472 45849
rect 44272 45840 44324 45892
rect 46480 45883 46532 45892
rect 40776 45772 40828 45824
rect 45652 45772 45704 45824
rect 46480 45849 46489 45883
rect 46489 45849 46523 45883
rect 46523 45849 46532 45883
rect 46480 45840 46532 45849
rect 46848 45772 46900 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 11612 45568 11664 45620
rect 20904 45611 20956 45620
rect 20904 45577 20913 45611
rect 20913 45577 20947 45611
rect 20947 45577 20956 45611
rect 20904 45568 20956 45577
rect 24584 45568 24636 45620
rect 25412 45611 25464 45620
rect 25412 45577 25421 45611
rect 25421 45577 25455 45611
rect 25455 45577 25464 45611
rect 25412 45568 25464 45577
rect 41420 45611 41472 45620
rect 41420 45577 41429 45611
rect 41429 45577 41463 45611
rect 41463 45577 41472 45611
rect 41420 45568 41472 45577
rect 42616 45568 42668 45620
rect 45100 45568 45152 45620
rect 45560 45568 45612 45620
rect 46388 45568 46440 45620
rect 43168 45543 43220 45552
rect 43168 45509 43177 45543
rect 43177 45509 43211 45543
rect 43211 45509 43220 45543
rect 43168 45500 43220 45509
rect 44180 45500 44232 45552
rect 1768 45475 1820 45484
rect 1768 45441 1777 45475
rect 1777 45441 1811 45475
rect 1811 45441 1820 45475
rect 1768 45432 1820 45441
rect 20720 45432 20772 45484
rect 25320 45475 25372 45484
rect 25320 45441 25329 45475
rect 25329 45441 25363 45475
rect 25363 45441 25372 45475
rect 25320 45432 25372 45441
rect 41052 45432 41104 45484
rect 2228 45364 2280 45416
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 44548 45407 44600 45416
rect 44548 45373 44557 45407
rect 44557 45373 44591 45407
rect 44591 45373 44600 45407
rect 44548 45364 44600 45373
rect 45100 45364 45152 45416
rect 45560 45407 45612 45416
rect 45560 45373 45569 45407
rect 45569 45373 45603 45407
rect 45603 45373 45612 45407
rect 46664 45500 46716 45552
rect 46848 45475 46900 45484
rect 46848 45441 46857 45475
rect 46857 45441 46891 45475
rect 46891 45441 46900 45475
rect 46848 45432 46900 45441
rect 45560 45364 45612 45373
rect 47124 45364 47176 45416
rect 46388 45296 46440 45348
rect 38476 45228 38528 45280
rect 47308 45228 47360 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2228 45067 2280 45076
rect 2228 45033 2237 45067
rect 2237 45033 2271 45067
rect 2271 45033 2280 45067
rect 2228 45024 2280 45033
rect 42708 45024 42760 45076
rect 44456 45067 44508 45076
rect 44456 45033 44465 45067
rect 44465 45033 44499 45067
rect 44499 45033 44508 45067
rect 44456 45024 44508 45033
rect 45100 45067 45152 45076
rect 45100 45033 45109 45067
rect 45109 45033 45143 45067
rect 45143 45033 45152 45067
rect 45100 45024 45152 45033
rect 45376 45024 45428 45076
rect 47032 44888 47084 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 2412 44820 2464 44872
rect 45008 44863 45060 44872
rect 45008 44829 45017 44863
rect 45017 44829 45051 44863
rect 45051 44829 45060 44863
rect 45008 44820 45060 44829
rect 45560 44820 45612 44872
rect 46204 44820 46256 44872
rect 47676 44752 47728 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 46480 44480 46532 44532
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 24584 44344 24636 44396
rect 44548 44344 44600 44396
rect 45744 44387 45796 44396
rect 45744 44353 45753 44387
rect 45753 44353 45787 44387
rect 45787 44353 45796 44387
rect 45744 44344 45796 44353
rect 46572 44344 46624 44396
rect 46664 44344 46716 44396
rect 41052 44208 41104 44260
rect 47584 44208 47636 44260
rect 20720 44140 20772 44192
rect 21364 44140 21416 44192
rect 46940 44183 46992 44192
rect 46940 44149 46949 44183
rect 46949 44149 46983 44183
rect 46983 44149 46992 44183
rect 46940 44140 46992 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 46940 43800 46992 43852
rect 48228 43800 48280 43852
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 47032 43299 47084 43308
rect 47032 43265 47041 43299
rect 47041 43265 47075 43299
rect 47075 43265 47084 43299
rect 47032 43256 47084 43265
rect 47768 43299 47820 43308
rect 47768 43265 47777 43299
rect 47777 43265 47811 43299
rect 47811 43265 47820 43299
rect 47768 43256 47820 43265
rect 1952 43188 2004 43240
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 46296 42687 46348 42696
rect 46296 42653 46305 42687
rect 46305 42653 46339 42687
rect 46339 42653 46348 42687
rect 46296 42644 46348 42653
rect 47676 42576 47728 42628
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 47676 42347 47728 42356
rect 47676 42313 47685 42347
rect 47685 42313 47719 42347
rect 47719 42313 47728 42347
rect 47676 42304 47728 42313
rect 46296 42168 46348 42220
rect 46940 42100 46992 42152
rect 47124 42100 47176 42152
rect 1400 41964 1452 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 47768 41624 47820 41676
rect 31760 41556 31812 41608
rect 48136 41599 48188 41608
rect 48136 41565 48145 41599
rect 48145 41565 48179 41599
rect 48179 41565 48188 41599
rect 48136 41556 48188 41565
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 27160 41420 27212 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 26240 41216 26292 41268
rect 27160 41191 27212 41200
rect 27160 41157 27169 41191
rect 27169 41157 27203 41191
rect 27203 41157 27212 41191
rect 27160 41148 27212 41157
rect 46480 41216 46532 41268
rect 14096 41080 14148 41132
rect 46388 41080 46440 41132
rect 47768 41123 47820 41132
rect 47768 41089 47777 41123
rect 47777 41089 47811 41123
rect 47811 41089 47820 41123
rect 47768 41080 47820 41089
rect 26056 41012 26108 41064
rect 42800 41012 42852 41064
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 26056 40579 26108 40588
rect 26056 40545 26065 40579
rect 26065 40545 26099 40579
rect 26099 40545 26108 40579
rect 26056 40536 26108 40545
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 45100 40511 45152 40520
rect 45100 40477 45109 40511
rect 45109 40477 45143 40511
rect 45143 40477 45152 40511
rect 45100 40468 45152 40477
rect 46848 40468 46900 40520
rect 47676 40511 47728 40520
rect 47676 40477 47685 40511
rect 47685 40477 47719 40511
rect 47719 40477 47728 40511
rect 47676 40468 47728 40477
rect 2136 40400 2188 40452
rect 28080 40400 28132 40452
rect 1860 40332 1912 40384
rect 46112 40375 46164 40384
rect 46112 40341 46121 40375
rect 46121 40341 46155 40375
rect 46155 40341 46164 40375
rect 46112 40332 46164 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 45928 40060 45980 40112
rect 46112 40035 46164 40044
rect 46112 40001 46121 40035
rect 46121 40001 46155 40035
rect 46155 40001 46164 40035
rect 46112 39992 46164 40001
rect 47584 40035 47636 40044
rect 47584 40001 47593 40035
rect 47593 40001 47627 40035
rect 47627 40001 47636 40035
rect 47584 39992 47636 40001
rect 42800 39856 42852 39908
rect 46480 39788 46532 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 47676 39516 47728 39568
rect 46480 39491 46532 39500
rect 46480 39457 46489 39491
rect 46489 39457 46523 39491
rect 46523 39457 46532 39491
rect 46480 39448 46532 39457
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 42064 38904 42116 38956
rect 45836 38947 45888 38956
rect 45836 38913 45845 38947
rect 45845 38913 45879 38947
rect 45879 38913 45888 38947
rect 45836 38904 45888 38913
rect 47860 38947 47912 38956
rect 47860 38913 47869 38947
rect 47869 38913 47903 38947
rect 47903 38913 47912 38947
rect 47860 38904 47912 38913
rect 46664 38836 46716 38888
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 45560 38403 45612 38412
rect 45560 38369 45569 38403
rect 45569 38369 45603 38403
rect 45603 38369 45612 38403
rect 45560 38360 45612 38369
rect 46020 38360 46072 38412
rect 45836 38292 45888 38344
rect 46296 38335 46348 38344
rect 46296 38301 46305 38335
rect 46305 38301 46339 38335
rect 46339 38301 46348 38335
rect 46296 38292 46348 38301
rect 47676 38224 47728 38276
rect 48136 38267 48188 38276
rect 48136 38233 48145 38267
rect 48145 38233 48179 38267
rect 48179 38233 48188 38267
rect 48136 38224 48188 38233
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 47676 37995 47728 38004
rect 47676 37961 47685 37995
rect 47685 37961 47719 37995
rect 47719 37961 47728 37995
rect 47676 37952 47728 37961
rect 25320 37884 25372 37936
rect 45836 37859 45888 37868
rect 45836 37825 45845 37859
rect 45845 37825 45879 37859
rect 45879 37825 45888 37859
rect 45836 37816 45888 37825
rect 47492 37816 47544 37868
rect 46204 37791 46256 37800
rect 46204 37757 46213 37791
rect 46213 37757 46247 37791
rect 46247 37757 46256 37791
rect 46204 37748 46256 37757
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 46296 37408 46348 37460
rect 1768 37204 1820 37256
rect 45836 37247 45888 37256
rect 45836 37213 45845 37247
rect 45845 37213 45879 37247
rect 45879 37213 45888 37247
rect 45836 37204 45888 37213
rect 46572 37136 46624 37188
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 46388 36839 46440 36848
rect 46388 36805 46397 36839
rect 46397 36805 46431 36839
rect 46431 36805 46440 36839
rect 46388 36796 46440 36805
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 45836 36771 45888 36780
rect 45836 36737 45845 36771
rect 45845 36737 45879 36771
rect 45879 36737 45888 36771
rect 45836 36728 45888 36737
rect 2228 36660 2280 36712
rect 2780 36703 2832 36712
rect 2780 36669 2789 36703
rect 2789 36669 2823 36703
rect 2823 36669 2832 36703
rect 2780 36660 2832 36669
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 46204 36116 46256 36168
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 1492 35436 1544 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 48136 35071 48188 35080
rect 48136 35037 48145 35071
rect 48145 35037 48179 35071
rect 48179 35037 48188 35071
rect 48136 35028 48188 35037
rect 47124 34892 47176 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 30564 34595 30616 34604
rect 29644 34527 29696 34536
rect 29644 34493 29653 34527
rect 29653 34493 29687 34527
rect 29687 34493 29696 34527
rect 29644 34484 29696 34493
rect 30564 34561 30573 34595
rect 30573 34561 30607 34595
rect 30607 34561 30616 34595
rect 30564 34552 30616 34561
rect 48136 34595 48188 34604
rect 48136 34561 48145 34595
rect 48145 34561 48179 34595
rect 48179 34561 48188 34595
rect 48136 34552 48188 34561
rect 31760 34484 31812 34536
rect 30380 34391 30432 34400
rect 30380 34357 30389 34391
rect 30389 34357 30423 34391
rect 30423 34357 30432 34391
rect 30380 34348 30432 34357
rect 47216 34348 47268 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 45836 34076 45888 34128
rect 24676 34008 24728 34060
rect 32220 34008 32272 34060
rect 47124 34051 47176 34060
rect 47124 34017 47133 34051
rect 47133 34017 47167 34051
rect 47167 34017 47176 34051
rect 47124 34008 47176 34017
rect 1308 33940 1360 33992
rect 20444 33940 20496 33992
rect 21088 33872 21140 33924
rect 21548 33872 21600 33924
rect 24492 33872 24544 33924
rect 30380 33872 30432 33924
rect 31852 33872 31904 33924
rect 47216 33915 47268 33924
rect 47216 33881 47225 33915
rect 47225 33881 47259 33915
rect 47259 33881 47268 33915
rect 47216 33872 47268 33881
rect 1584 33804 1636 33856
rect 22284 33847 22336 33856
rect 22284 33813 22293 33847
rect 22293 33813 22327 33847
rect 22327 33813 22336 33847
rect 22284 33804 22336 33813
rect 23480 33804 23532 33856
rect 24768 33847 24820 33856
rect 24768 33813 24777 33847
rect 24777 33813 24811 33847
rect 24811 33813 24820 33847
rect 24768 33804 24820 33813
rect 31668 33804 31720 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 11704 33600 11756 33652
rect 14648 33532 14700 33584
rect 25688 33532 25740 33584
rect 29644 33532 29696 33584
rect 19432 33464 19484 33516
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 23480 33507 23532 33516
rect 23480 33473 23489 33507
rect 23489 33473 23523 33507
rect 23523 33473 23532 33507
rect 23480 33464 23532 33473
rect 29920 33464 29972 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 2320 33396 2372 33448
rect 22468 33439 22520 33448
rect 22468 33405 22477 33439
rect 22477 33405 22511 33439
rect 22511 33405 22520 33439
rect 22468 33396 22520 33405
rect 23572 33396 23624 33448
rect 23940 33439 23992 33448
rect 23940 33405 23949 33439
rect 23949 33405 23983 33439
rect 23983 33405 23992 33439
rect 23940 33396 23992 33405
rect 20444 33328 20496 33380
rect 19340 33260 19392 33312
rect 21088 33303 21140 33312
rect 21088 33269 21097 33303
rect 21097 33269 21131 33303
rect 21131 33269 21140 33303
rect 21088 33260 21140 33269
rect 22008 33303 22060 33312
rect 22008 33269 22017 33303
rect 22017 33269 22051 33303
rect 22051 33269 22060 33303
rect 22008 33260 22060 33269
rect 27252 33396 27304 33448
rect 28172 33439 28224 33448
rect 28172 33405 28181 33439
rect 28181 33405 28215 33439
rect 28215 33405 28224 33439
rect 28172 33396 28224 33405
rect 29828 33396 29880 33448
rect 31668 33464 31720 33516
rect 47768 33507 47820 33516
rect 47768 33473 47777 33507
rect 47777 33473 47811 33507
rect 47811 33473 47820 33507
rect 47768 33464 47820 33473
rect 32128 33396 32180 33448
rect 24768 33260 24820 33312
rect 29644 33303 29696 33312
rect 29644 33269 29653 33303
rect 29653 33269 29687 33303
rect 29687 33269 29696 33303
rect 29644 33260 29696 33269
rect 29736 33260 29788 33312
rect 30840 33303 30892 33312
rect 30840 33269 30849 33303
rect 30849 33269 30883 33303
rect 30883 33269 30892 33303
rect 30840 33260 30892 33269
rect 47860 33303 47912 33312
rect 47860 33269 47869 33303
rect 47869 33269 47903 33303
rect 47903 33269 47912 33303
rect 47860 33260 47912 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19156 33056 19208 33108
rect 21272 33056 21324 33108
rect 24492 33056 24544 33108
rect 24584 33056 24636 33108
rect 25688 33099 25740 33108
rect 1492 32988 1544 33040
rect 1860 32988 1912 33040
rect 24860 32988 24912 33040
rect 1584 32963 1636 32972
rect 1584 32929 1593 32963
rect 1593 32929 1627 32963
rect 1627 32929 1636 32963
rect 1584 32920 1636 32929
rect 12532 32852 12584 32904
rect 12624 32895 12676 32904
rect 12624 32861 12633 32895
rect 12633 32861 12667 32895
rect 12667 32861 12676 32895
rect 19432 32920 19484 32972
rect 22008 32920 22060 32972
rect 12624 32852 12676 32861
rect 3240 32827 3292 32836
rect 3240 32793 3249 32827
rect 3249 32793 3283 32827
rect 3283 32793 3292 32827
rect 3240 32784 3292 32793
rect 11980 32716 12032 32768
rect 17776 32716 17828 32768
rect 22744 32920 22796 32972
rect 25688 33065 25697 33099
rect 25697 33065 25731 33099
rect 25731 33065 25740 33099
rect 25688 33056 25740 33065
rect 28172 33056 28224 33108
rect 30564 33099 30616 33108
rect 30564 33065 30573 33099
rect 30573 33065 30607 33099
rect 30607 33065 30616 33099
rect 30564 33056 30616 33065
rect 31852 33099 31904 33108
rect 31852 33065 31861 33099
rect 31861 33065 31895 33099
rect 31895 33065 31904 33099
rect 31852 33056 31904 33065
rect 31944 33056 31996 33108
rect 37280 33056 37332 33108
rect 25044 32988 25096 33040
rect 31116 32988 31168 33040
rect 35072 32988 35124 33040
rect 37464 32988 37516 33040
rect 23388 32852 23440 32904
rect 23572 32895 23624 32904
rect 23572 32861 23581 32895
rect 23581 32861 23615 32895
rect 23615 32861 23624 32895
rect 23572 32852 23624 32861
rect 24032 32852 24084 32904
rect 24584 32852 24636 32904
rect 25044 32852 25096 32904
rect 26332 32852 26384 32904
rect 27896 32895 27948 32904
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 27896 32852 27948 32861
rect 27988 32852 28040 32904
rect 29644 32920 29696 32972
rect 28448 32895 28500 32904
rect 28448 32861 28457 32895
rect 28457 32861 28491 32895
rect 28491 32861 28500 32895
rect 30840 32920 30892 32972
rect 28448 32852 28500 32861
rect 29828 32852 29880 32904
rect 30012 32895 30064 32904
rect 30012 32861 30021 32895
rect 30021 32861 30055 32895
rect 30055 32861 30064 32895
rect 30012 32852 30064 32861
rect 31668 32852 31720 32904
rect 31760 32895 31812 32904
rect 31760 32861 31769 32895
rect 31769 32861 31803 32895
rect 31803 32861 31812 32895
rect 36544 32920 36596 32972
rect 31760 32852 31812 32861
rect 32772 32852 32824 32904
rect 36176 32852 36228 32904
rect 46296 32895 46348 32904
rect 46296 32861 46305 32895
rect 46305 32861 46339 32895
rect 46339 32861 46348 32895
rect 46296 32852 46348 32861
rect 19156 32784 19208 32836
rect 21088 32827 21140 32836
rect 21088 32793 21097 32827
rect 21097 32793 21131 32827
rect 21131 32793 21140 32827
rect 21088 32784 21140 32793
rect 24952 32784 25004 32836
rect 40040 32784 40092 32836
rect 47676 32784 47728 32836
rect 48136 32827 48188 32836
rect 48136 32793 48145 32827
rect 48145 32793 48179 32827
rect 48179 32793 48188 32827
rect 48136 32784 48188 32793
rect 22284 32716 22336 32768
rect 22744 32716 22796 32768
rect 28448 32716 28500 32768
rect 28816 32716 28868 32768
rect 32036 32716 32088 32768
rect 33416 32759 33468 32768
rect 33416 32725 33425 32759
rect 33425 32725 33459 32759
rect 33459 32725 33468 32759
rect 33416 32716 33468 32725
rect 36176 32759 36228 32768
rect 36176 32725 36185 32759
rect 36185 32725 36219 32759
rect 36219 32725 36228 32759
rect 36176 32716 36228 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 22468 32512 22520 32564
rect 25044 32512 25096 32564
rect 27896 32512 27948 32564
rect 2320 32487 2372 32496
rect 2320 32453 2329 32487
rect 2329 32453 2363 32487
rect 2363 32453 2372 32487
rect 2320 32444 2372 32453
rect 12716 32444 12768 32496
rect 19340 32487 19392 32496
rect 14556 32376 14608 32428
rect 19340 32453 19349 32487
rect 19349 32453 19383 32487
rect 19383 32453 19392 32487
rect 19340 32444 19392 32453
rect 31944 32512 31996 32564
rect 33416 32512 33468 32564
rect 36176 32512 36228 32564
rect 34060 32444 34112 32496
rect 47676 32555 47728 32564
rect 47676 32521 47685 32555
rect 47685 32521 47719 32555
rect 47719 32521 47728 32555
rect 47676 32512 47728 32521
rect 46664 32444 46716 32496
rect 15660 32419 15712 32428
rect 15660 32385 15669 32419
rect 15669 32385 15703 32419
rect 15703 32385 15712 32419
rect 15660 32376 15712 32385
rect 16396 32376 16448 32428
rect 22284 32376 22336 32428
rect 22560 32376 22612 32428
rect 24216 32376 24268 32428
rect 24768 32376 24820 32428
rect 25412 32376 25464 32428
rect 28632 32376 28684 32428
rect 29736 32376 29788 32428
rect 30012 32376 30064 32428
rect 32220 32419 32272 32428
rect 2412 32308 2464 32360
rect 3240 32351 3292 32360
rect 3240 32317 3249 32351
rect 3249 32317 3283 32351
rect 3283 32317 3292 32351
rect 3240 32308 3292 32317
rect 12624 32308 12676 32360
rect 14464 32308 14516 32360
rect 17592 32308 17644 32360
rect 22468 32308 22520 32360
rect 25136 32308 25188 32360
rect 14188 32240 14240 32292
rect 17776 32240 17828 32292
rect 1400 32172 1452 32224
rect 11704 32215 11756 32224
rect 11704 32181 11713 32215
rect 11713 32181 11747 32215
rect 11747 32181 11756 32215
rect 11704 32172 11756 32181
rect 13176 32215 13228 32224
rect 13176 32181 13185 32215
rect 13185 32181 13219 32215
rect 13219 32181 13228 32215
rect 13176 32172 13228 32181
rect 15200 32172 15252 32224
rect 15476 32215 15528 32224
rect 15476 32181 15485 32215
rect 15485 32181 15519 32215
rect 15519 32181 15528 32215
rect 15476 32172 15528 32181
rect 16764 32215 16816 32224
rect 16764 32181 16773 32215
rect 16773 32181 16807 32215
rect 16807 32181 16816 32215
rect 16764 32172 16816 32181
rect 23480 32172 23532 32224
rect 24676 32172 24728 32224
rect 29644 32308 29696 32360
rect 32220 32385 32229 32419
rect 32229 32385 32263 32419
rect 32263 32385 32272 32419
rect 32220 32376 32272 32385
rect 32128 32308 32180 32360
rect 34520 32308 34572 32360
rect 35072 32376 35124 32428
rect 37464 32419 37516 32428
rect 37464 32385 37473 32419
rect 37473 32385 37507 32419
rect 37507 32385 37516 32419
rect 37464 32376 37516 32385
rect 46848 32376 46900 32428
rect 47216 32376 47268 32428
rect 36176 32351 36228 32360
rect 32036 32240 32088 32292
rect 26332 32172 26384 32224
rect 28816 32215 28868 32224
rect 28816 32181 28825 32215
rect 28825 32181 28859 32215
rect 28859 32181 28868 32215
rect 28816 32172 28868 32181
rect 29920 32172 29972 32224
rect 33232 32172 33284 32224
rect 36176 32317 36185 32351
rect 36185 32317 36219 32351
rect 36219 32317 36228 32351
rect 36176 32308 36228 32317
rect 36360 32351 36412 32360
rect 36360 32317 36369 32351
rect 36369 32317 36403 32351
rect 36403 32317 36412 32351
rect 36360 32308 36412 32317
rect 33876 32172 33928 32224
rect 36084 32172 36136 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 14464 32011 14516 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 11704 31875 11756 31884
rect 11704 31841 11713 31875
rect 11713 31841 11747 31875
rect 11747 31841 11756 31875
rect 11704 31832 11756 31841
rect 11980 31875 12032 31884
rect 11980 31841 11989 31875
rect 11989 31841 12023 31875
rect 12023 31841 12032 31875
rect 11980 31832 12032 31841
rect 12624 31832 12676 31884
rect 14464 31977 14473 32011
rect 14473 31977 14507 32011
rect 14507 31977 14516 32011
rect 14464 31968 14516 31977
rect 14556 31968 14608 32020
rect 16856 31968 16908 32020
rect 17684 31968 17736 32020
rect 21548 31968 21600 32020
rect 32772 32011 32824 32020
rect 32772 31977 32781 32011
rect 32781 31977 32815 32011
rect 32815 31977 32824 32011
rect 32772 31968 32824 31977
rect 34060 32011 34112 32020
rect 34060 31977 34069 32011
rect 34069 31977 34103 32011
rect 34103 31977 34112 32011
rect 34060 31968 34112 31977
rect 36268 31968 36320 32020
rect 46296 31968 46348 32020
rect 14372 31832 14424 31884
rect 15200 31875 15252 31884
rect 15200 31841 15209 31875
rect 15209 31841 15243 31875
rect 15243 31841 15252 31875
rect 15200 31832 15252 31841
rect 15476 31875 15528 31884
rect 15476 31841 15485 31875
rect 15485 31841 15519 31875
rect 15519 31841 15528 31875
rect 15476 31832 15528 31841
rect 16672 31832 16724 31884
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 9312 31696 9364 31748
rect 10784 31696 10836 31748
rect 12440 31696 12492 31748
rect 3976 31628 4028 31680
rect 12808 31628 12860 31680
rect 12900 31628 12952 31680
rect 14188 31764 14240 31816
rect 16764 31764 16816 31816
rect 17316 31832 17368 31884
rect 17592 31807 17644 31816
rect 17592 31773 17601 31807
rect 17601 31773 17635 31807
rect 17635 31773 17644 31807
rect 17592 31764 17644 31773
rect 17684 31807 17736 31816
rect 17684 31773 17693 31807
rect 17693 31773 17727 31807
rect 17727 31773 17736 31807
rect 17684 31764 17736 31773
rect 32220 31900 32272 31952
rect 20996 31832 21048 31884
rect 27252 31875 27304 31884
rect 14648 31696 14700 31748
rect 14464 31628 14516 31680
rect 17040 31696 17092 31748
rect 18144 31696 18196 31748
rect 19156 31764 19208 31816
rect 27252 31841 27261 31875
rect 27261 31841 27295 31875
rect 27295 31841 27304 31875
rect 27252 31832 27304 31841
rect 28540 31832 28592 31884
rect 32036 31832 32088 31884
rect 32496 31832 32548 31884
rect 36084 31875 36136 31884
rect 36084 31841 36093 31875
rect 36093 31841 36127 31875
rect 36127 31841 36136 31875
rect 36084 31832 36136 31841
rect 26332 31764 26384 31816
rect 19432 31696 19484 31748
rect 26240 31696 26292 31748
rect 31760 31764 31812 31816
rect 33968 31807 34020 31816
rect 33968 31773 33977 31807
rect 33977 31773 34011 31807
rect 34011 31773 34020 31807
rect 33968 31764 34020 31773
rect 27988 31696 28040 31748
rect 33232 31739 33284 31748
rect 33232 31705 33241 31739
rect 33241 31705 33275 31739
rect 33275 31705 33284 31739
rect 33232 31696 33284 31705
rect 33324 31696 33376 31748
rect 37372 31696 37424 31748
rect 16948 31628 17000 31680
rect 17776 31671 17828 31680
rect 17776 31637 17785 31671
rect 17785 31637 17819 31671
rect 17819 31637 17828 31671
rect 17776 31628 17828 31637
rect 25596 31628 25648 31680
rect 29184 31628 29236 31680
rect 31024 31628 31076 31680
rect 33600 31628 33652 31680
rect 33876 31628 33928 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1584 31424 1636 31476
rect 2228 31288 2280 31340
rect 7196 31288 7248 31340
rect 9404 31424 9456 31476
rect 12256 31424 12308 31476
rect 12624 31424 12676 31476
rect 12808 31424 12860 31476
rect 8760 31220 8812 31272
rect 11520 31331 11572 31340
rect 11520 31297 11529 31331
rect 11529 31297 11563 31331
rect 11563 31297 11572 31331
rect 11520 31288 11572 31297
rect 12900 31356 12952 31408
rect 13176 31399 13228 31408
rect 13176 31365 13185 31399
rect 13185 31365 13219 31399
rect 13219 31365 13228 31399
rect 13176 31356 13228 31365
rect 14188 31356 14240 31408
rect 14556 31424 14608 31476
rect 15660 31424 15712 31476
rect 16672 31399 16724 31408
rect 16672 31365 16681 31399
rect 16681 31365 16715 31399
rect 16715 31365 16724 31399
rect 16672 31356 16724 31365
rect 17776 31424 17828 31476
rect 23940 31424 23992 31476
rect 18144 31356 18196 31408
rect 26240 31424 26292 31476
rect 27988 31424 28040 31476
rect 28540 31424 28592 31476
rect 36176 31424 36228 31476
rect 37372 31467 37424 31476
rect 37372 31433 37381 31467
rect 37381 31433 37415 31467
rect 37415 31433 37424 31467
rect 37372 31424 37424 31433
rect 12808 31288 12860 31340
rect 16764 31288 16816 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 19248 31288 19300 31340
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 22468 31331 22520 31340
rect 22468 31297 22477 31331
rect 22477 31297 22511 31331
rect 22511 31297 22520 31331
rect 22468 31288 22520 31297
rect 25596 31356 25648 31408
rect 27620 31288 27672 31340
rect 27896 31331 27948 31340
rect 27896 31297 27905 31331
rect 27905 31297 27939 31331
rect 27939 31297 27948 31331
rect 27896 31288 27948 31297
rect 28356 31288 28408 31340
rect 28448 31331 28500 31340
rect 28448 31297 28457 31331
rect 28457 31297 28491 31331
rect 28491 31297 28500 31331
rect 29276 31331 29328 31340
rect 28448 31288 28500 31297
rect 29276 31297 29285 31331
rect 29285 31297 29319 31331
rect 29319 31297 29328 31331
rect 29276 31288 29328 31297
rect 33600 31331 33652 31340
rect 33600 31297 33609 31331
rect 33609 31297 33643 31331
rect 33643 31297 33652 31331
rect 33600 31288 33652 31297
rect 36176 31288 36228 31340
rect 37096 31288 37148 31340
rect 37280 31331 37332 31340
rect 37280 31297 37289 31331
rect 37289 31297 37323 31331
rect 37323 31297 37332 31331
rect 37280 31288 37332 31297
rect 10784 31220 10836 31272
rect 12900 31263 12952 31272
rect 9496 31127 9548 31136
rect 9496 31093 9505 31127
rect 9505 31093 9539 31127
rect 9539 31093 9548 31127
rect 9496 31084 9548 31093
rect 9680 31084 9732 31136
rect 10692 31084 10744 31136
rect 12532 31152 12584 31204
rect 12440 31084 12492 31136
rect 12900 31229 12909 31263
rect 12909 31229 12943 31263
rect 12943 31229 12952 31263
rect 12900 31220 12952 31229
rect 12808 31152 12860 31204
rect 14648 31220 14700 31272
rect 16212 31220 16264 31272
rect 17868 31263 17920 31272
rect 17868 31229 17877 31263
rect 17877 31229 17911 31263
rect 17911 31229 17920 31263
rect 17868 31220 17920 31229
rect 18144 31263 18196 31272
rect 18144 31229 18153 31263
rect 18153 31229 18187 31263
rect 18187 31229 18196 31263
rect 18144 31220 18196 31229
rect 18236 31220 18288 31272
rect 19156 31220 19208 31272
rect 22560 31263 22612 31272
rect 22560 31229 22569 31263
rect 22569 31229 22603 31263
rect 22603 31229 22612 31263
rect 22560 31220 22612 31229
rect 23020 31220 23072 31272
rect 24860 31263 24912 31272
rect 24860 31229 24869 31263
rect 24869 31229 24903 31263
rect 24903 31229 24912 31263
rect 24860 31220 24912 31229
rect 29184 31220 29236 31272
rect 33508 31263 33560 31272
rect 33508 31229 33517 31263
rect 33517 31229 33551 31263
rect 33551 31229 33560 31263
rect 33508 31220 33560 31229
rect 34520 31220 34572 31272
rect 17040 31084 17092 31136
rect 22100 31127 22152 31136
rect 22100 31093 22109 31127
rect 22109 31093 22143 31127
rect 22143 31093 22152 31127
rect 45560 31152 45612 31204
rect 46020 31152 46072 31204
rect 22100 31084 22152 31093
rect 25964 31084 26016 31136
rect 29000 31084 29052 31136
rect 29644 31084 29696 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7840 30880 7892 30932
rect 12900 30923 12952 30932
rect 9496 30812 9548 30864
rect 12900 30889 12909 30923
rect 12909 30889 12943 30923
rect 12943 30889 12952 30923
rect 12900 30880 12952 30889
rect 14188 30923 14240 30932
rect 14188 30889 14197 30923
rect 14197 30889 14231 30923
rect 14231 30889 14240 30923
rect 14188 30880 14240 30889
rect 18144 30880 18196 30932
rect 19248 30880 19300 30932
rect 9680 30787 9732 30796
rect 9680 30753 9689 30787
rect 9689 30753 9723 30787
rect 9723 30753 9732 30787
rect 9680 30744 9732 30753
rect 12440 30676 12492 30728
rect 12716 30676 12768 30728
rect 10692 30608 10744 30660
rect 9404 30540 9456 30592
rect 12624 30608 12676 30660
rect 13268 30676 13320 30728
rect 14648 30676 14700 30728
rect 17040 30676 17092 30728
rect 13360 30608 13412 30660
rect 16856 30608 16908 30660
rect 16212 30583 16264 30592
rect 16212 30549 16221 30583
rect 16221 30549 16255 30583
rect 16255 30549 16264 30583
rect 16212 30540 16264 30549
rect 17868 30812 17920 30864
rect 17592 30787 17644 30796
rect 17592 30753 17601 30787
rect 17601 30753 17635 30787
rect 17635 30753 17644 30787
rect 17592 30744 17644 30753
rect 20444 30787 20496 30796
rect 20444 30753 20453 30787
rect 20453 30753 20487 30787
rect 20487 30753 20496 30787
rect 20444 30744 20496 30753
rect 24860 30880 24912 30932
rect 27620 30880 27672 30932
rect 23204 30812 23256 30864
rect 25228 30812 25280 30864
rect 26148 30812 26200 30864
rect 27896 30880 27948 30932
rect 28356 30880 28408 30932
rect 30104 30880 30156 30932
rect 29000 30812 29052 30864
rect 29276 30812 29328 30864
rect 18236 30676 18288 30728
rect 19248 30719 19300 30728
rect 18144 30608 18196 30660
rect 19248 30685 19257 30719
rect 19257 30685 19291 30719
rect 19291 30685 19300 30719
rect 19248 30676 19300 30685
rect 22652 30719 22704 30728
rect 22652 30685 22661 30719
rect 22661 30685 22695 30719
rect 22695 30685 22704 30719
rect 22652 30676 22704 30685
rect 22744 30676 22796 30728
rect 21180 30608 21232 30660
rect 23480 30676 23532 30728
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 25044 30676 25096 30728
rect 25412 30744 25464 30796
rect 25320 30719 25372 30728
rect 25320 30685 25329 30719
rect 25329 30685 25363 30719
rect 25363 30685 25372 30719
rect 25320 30676 25372 30685
rect 24768 30608 24820 30660
rect 25412 30608 25464 30660
rect 22284 30540 22336 30592
rect 23204 30540 23256 30592
rect 23480 30540 23532 30592
rect 25688 30676 25740 30728
rect 29000 30676 29052 30728
rect 29736 30719 29788 30728
rect 29736 30685 29745 30719
rect 29745 30685 29779 30719
rect 29779 30685 29788 30719
rect 29736 30676 29788 30685
rect 31668 30744 31720 30796
rect 33508 30880 33560 30932
rect 36176 30923 36228 30932
rect 36176 30889 36185 30923
rect 36185 30889 36219 30923
rect 36219 30889 36228 30923
rect 36176 30880 36228 30889
rect 31024 30719 31076 30728
rect 31024 30685 31033 30719
rect 31033 30685 31067 30719
rect 31067 30685 31076 30719
rect 31024 30676 31076 30685
rect 32956 30719 33008 30728
rect 29184 30608 29236 30660
rect 30012 30608 30064 30660
rect 29000 30583 29052 30592
rect 29000 30549 29009 30583
rect 29009 30549 29043 30583
rect 29043 30549 29052 30583
rect 29000 30540 29052 30549
rect 32956 30685 32965 30719
rect 32965 30685 32999 30719
rect 32999 30685 33008 30719
rect 32956 30676 33008 30685
rect 34520 30744 34572 30796
rect 36268 30719 36320 30728
rect 36268 30685 36277 30719
rect 36277 30685 36311 30719
rect 36311 30685 36320 30719
rect 36268 30676 36320 30685
rect 36820 30676 36872 30728
rect 37004 30608 37056 30660
rect 32956 30540 33008 30592
rect 34796 30540 34848 30592
rect 37096 30583 37148 30592
rect 37096 30549 37105 30583
rect 37105 30549 37139 30583
rect 37139 30549 37148 30583
rect 37096 30540 37148 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 17592 30336 17644 30388
rect 22652 30336 22704 30388
rect 24952 30336 25004 30388
rect 11520 30200 11572 30252
rect 13176 30175 13228 30184
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 3700 30064 3752 30116
rect 17040 30268 17092 30320
rect 21180 30311 21232 30320
rect 21180 30277 21189 30311
rect 21189 30277 21223 30311
rect 21223 30277 21232 30311
rect 21180 30268 21232 30277
rect 23020 30311 23072 30320
rect 23020 30277 23029 30311
rect 23029 30277 23063 30311
rect 23063 30277 23072 30311
rect 23020 30268 23072 30277
rect 16948 30200 17000 30252
rect 17316 30243 17368 30252
rect 17316 30209 17325 30243
rect 17325 30209 17359 30243
rect 17359 30209 17368 30243
rect 17316 30200 17368 30209
rect 20996 30200 21048 30252
rect 16856 30132 16908 30184
rect 17316 30064 17368 30116
rect 22468 30200 22520 30252
rect 23204 30243 23256 30252
rect 23204 30209 23213 30243
rect 23213 30209 23247 30243
rect 23247 30209 23256 30243
rect 23204 30200 23256 30209
rect 24676 30268 24728 30320
rect 25044 30268 25096 30320
rect 25688 30243 25740 30252
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 25688 30200 25740 30209
rect 30104 30268 30156 30320
rect 31944 30268 31996 30320
rect 25964 30200 26016 30252
rect 29000 30200 29052 30252
rect 24216 30132 24268 30184
rect 31116 30243 31168 30252
rect 31116 30209 31125 30243
rect 31125 30209 31159 30243
rect 31159 30209 31168 30243
rect 34244 30268 34296 30320
rect 31116 30200 31168 30209
rect 37648 30200 37700 30252
rect 38476 30243 38528 30252
rect 38476 30209 38485 30243
rect 38485 30209 38519 30243
rect 38519 30209 38528 30243
rect 38476 30200 38528 30209
rect 31024 30132 31076 30184
rect 32220 30132 32272 30184
rect 32680 30132 32732 30184
rect 33508 30175 33560 30184
rect 33508 30141 33517 30175
rect 33517 30141 33551 30175
rect 33551 30141 33560 30175
rect 33508 30132 33560 30141
rect 35348 30132 35400 30184
rect 35992 30132 36044 30184
rect 37096 30132 37148 30184
rect 38292 30175 38344 30184
rect 38292 30141 38301 30175
rect 38301 30141 38335 30175
rect 38335 30141 38344 30175
rect 38292 30132 38344 30141
rect 24952 30064 25004 30116
rect 25136 30107 25188 30116
rect 25136 30073 25145 30107
rect 25145 30073 25179 30107
rect 25179 30073 25188 30107
rect 25136 30064 25188 30073
rect 9956 30039 10008 30048
rect 9956 30005 9965 30039
rect 9965 30005 9999 30039
rect 9999 30005 10008 30039
rect 9956 29996 10008 30005
rect 22100 30039 22152 30048
rect 22100 30005 22109 30039
rect 22109 30005 22143 30039
rect 22143 30005 22152 30039
rect 22100 29996 22152 30005
rect 23296 29996 23348 30048
rect 24216 29996 24268 30048
rect 24400 29996 24452 30048
rect 24676 29996 24728 30048
rect 27804 30064 27856 30116
rect 28632 30064 28684 30116
rect 29000 30064 29052 30116
rect 35440 30064 35492 30116
rect 37832 30064 37884 30116
rect 25412 29996 25464 30048
rect 26148 29996 26200 30048
rect 28264 29996 28316 30048
rect 30012 30039 30064 30048
rect 30012 30005 30021 30039
rect 30021 30005 30055 30039
rect 30055 30005 30064 30039
rect 30012 29996 30064 30005
rect 30564 29996 30616 30048
rect 31484 30039 31536 30048
rect 31484 30005 31493 30039
rect 31493 30005 31527 30039
rect 31527 30005 31536 30039
rect 31484 29996 31536 30005
rect 32864 29996 32916 30048
rect 34520 29996 34572 30048
rect 37464 29996 37516 30048
rect 38016 29996 38068 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 13176 29792 13228 29844
rect 13268 29835 13320 29844
rect 13268 29801 13277 29835
rect 13277 29801 13311 29835
rect 13311 29801 13320 29835
rect 13268 29792 13320 29801
rect 8392 29631 8444 29640
rect 8392 29597 8401 29631
rect 8401 29597 8435 29631
rect 8435 29597 8444 29631
rect 8392 29588 8444 29597
rect 8944 29631 8996 29640
rect 8944 29597 8953 29631
rect 8953 29597 8987 29631
rect 8987 29597 8996 29631
rect 8944 29588 8996 29597
rect 11520 29656 11572 29708
rect 13452 29724 13504 29776
rect 20536 29724 20588 29776
rect 23112 29724 23164 29776
rect 24676 29792 24728 29844
rect 25228 29792 25280 29844
rect 28724 29792 28776 29844
rect 29000 29835 29052 29844
rect 29000 29801 29009 29835
rect 29009 29801 29043 29835
rect 29043 29801 29052 29835
rect 29000 29792 29052 29801
rect 31116 29792 31168 29844
rect 31668 29835 31720 29844
rect 31668 29801 31677 29835
rect 31677 29801 31711 29835
rect 31711 29801 31720 29835
rect 31668 29792 31720 29801
rect 34244 29792 34296 29844
rect 35348 29835 35400 29844
rect 35348 29801 35357 29835
rect 35357 29801 35391 29835
rect 35391 29801 35400 29835
rect 35348 29792 35400 29801
rect 35992 29835 36044 29844
rect 35992 29801 36001 29835
rect 36001 29801 36035 29835
rect 36035 29801 36044 29835
rect 35992 29792 36044 29801
rect 36084 29792 36136 29844
rect 37648 29792 37700 29844
rect 17224 29699 17276 29708
rect 17224 29665 17233 29699
rect 17233 29665 17267 29699
rect 17267 29665 17276 29699
rect 17224 29656 17276 29665
rect 18236 29656 18288 29708
rect 12624 29588 12676 29640
rect 12900 29588 12952 29640
rect 13360 29588 13412 29640
rect 16304 29588 16356 29640
rect 17316 29631 17368 29640
rect 17316 29597 17325 29631
rect 17325 29597 17359 29631
rect 17359 29597 17368 29631
rect 17316 29588 17368 29597
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 22560 29588 22612 29640
rect 23296 29631 23348 29640
rect 9956 29520 10008 29572
rect 14556 29563 14608 29572
rect 14556 29529 14565 29563
rect 14565 29529 14599 29563
rect 14599 29529 14608 29563
rect 14556 29520 14608 29529
rect 23296 29597 23305 29631
rect 23305 29597 23339 29631
rect 23339 29597 23348 29631
rect 23296 29588 23348 29597
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 24400 29631 24452 29640
rect 24400 29597 24409 29631
rect 24409 29597 24443 29631
rect 24443 29597 24452 29631
rect 24400 29588 24452 29597
rect 24492 29631 24544 29640
rect 24492 29597 24501 29631
rect 24501 29597 24535 29631
rect 24535 29597 24544 29631
rect 24492 29588 24544 29597
rect 26240 29656 26292 29708
rect 27252 29699 27304 29708
rect 27252 29665 27261 29699
rect 27261 29665 27295 29699
rect 27295 29665 27304 29699
rect 27252 29656 27304 29665
rect 31024 29656 31076 29708
rect 31944 29656 31996 29708
rect 33508 29724 33560 29776
rect 26332 29588 26384 29640
rect 29828 29588 29880 29640
rect 10692 29495 10744 29504
rect 10692 29461 10701 29495
rect 10701 29461 10735 29495
rect 10735 29461 10744 29495
rect 10692 29452 10744 29461
rect 11428 29452 11480 29504
rect 15936 29495 15988 29504
rect 15936 29461 15945 29495
rect 15945 29461 15979 29495
rect 15979 29461 15988 29495
rect 15936 29452 15988 29461
rect 17960 29452 18012 29504
rect 19340 29495 19392 29504
rect 19340 29461 19349 29495
rect 19349 29461 19383 29495
rect 19383 29461 19392 29495
rect 19340 29452 19392 29461
rect 22468 29452 22520 29504
rect 23940 29452 23992 29504
rect 27528 29520 27580 29572
rect 28540 29520 28592 29572
rect 26608 29495 26660 29504
rect 26608 29461 26617 29495
rect 26617 29461 26651 29495
rect 26651 29461 26660 29495
rect 26608 29452 26660 29461
rect 27804 29452 27856 29504
rect 30748 29588 30800 29640
rect 31484 29588 31536 29640
rect 32864 29631 32916 29640
rect 32864 29597 32873 29631
rect 32873 29597 32907 29631
rect 32907 29597 32916 29631
rect 32864 29588 32916 29597
rect 33232 29588 33284 29640
rect 33968 29588 34020 29640
rect 34520 29656 34572 29708
rect 34612 29588 34664 29640
rect 29736 29452 29788 29504
rect 32772 29452 32824 29504
rect 32956 29495 33008 29504
rect 32956 29461 32965 29495
rect 32965 29461 32999 29495
rect 32999 29461 33008 29495
rect 32956 29452 33008 29461
rect 34796 29631 34848 29640
rect 34796 29597 34806 29631
rect 34806 29597 34840 29631
rect 34840 29597 34848 29631
rect 34796 29588 34848 29597
rect 35440 29656 35492 29708
rect 36820 29699 36872 29708
rect 36820 29665 36829 29699
rect 36829 29665 36863 29699
rect 36863 29665 36872 29699
rect 36820 29656 36872 29665
rect 46940 29656 46992 29708
rect 35808 29588 35860 29640
rect 36084 29588 36136 29640
rect 36452 29588 36504 29640
rect 47400 29588 47452 29640
rect 35716 29520 35768 29572
rect 35992 29452 36044 29504
rect 36176 29495 36228 29504
rect 36176 29461 36185 29495
rect 36185 29461 36219 29495
rect 36219 29461 36228 29495
rect 36176 29452 36228 29461
rect 37004 29520 37056 29572
rect 37924 29520 37976 29572
rect 38476 29520 38528 29572
rect 37648 29452 37700 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 8392 29248 8444 29300
rect 13360 29248 13412 29300
rect 17316 29248 17368 29300
rect 20996 29248 21048 29300
rect 23664 29248 23716 29300
rect 25136 29248 25188 29300
rect 27344 29248 27396 29300
rect 28724 29291 28776 29300
rect 8944 29180 8996 29232
rect 18236 29223 18288 29232
rect 7104 29112 7156 29164
rect 8760 29155 8812 29164
rect 8760 29121 8769 29155
rect 8769 29121 8803 29155
rect 8803 29121 8812 29155
rect 8760 29112 8812 29121
rect 11520 29112 11572 29164
rect 15476 29155 15528 29164
rect 15476 29121 15485 29155
rect 15485 29121 15519 29155
rect 15519 29121 15528 29155
rect 15476 29112 15528 29121
rect 17040 29112 17092 29164
rect 11152 29044 11204 29096
rect 12164 29044 12216 29096
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 16212 29044 16264 29096
rect 16856 29044 16908 29096
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 18236 29189 18245 29223
rect 18245 29189 18279 29223
rect 18279 29189 18288 29223
rect 18236 29180 18288 29189
rect 17960 29155 18012 29164
rect 17960 29121 17969 29155
rect 17969 29121 18003 29155
rect 18003 29121 18012 29155
rect 17960 29112 18012 29121
rect 19340 29112 19392 29164
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 23112 29155 23164 29164
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 23112 29112 23164 29121
rect 23572 29087 23624 29096
rect 9036 29019 9088 29028
rect 9036 28985 9045 29019
rect 9045 28985 9079 29019
rect 9079 28985 9088 29019
rect 9036 28976 9088 28985
rect 17960 28976 18012 29028
rect 23572 29053 23581 29087
rect 23581 29053 23615 29087
rect 23615 29053 23624 29087
rect 23572 29044 23624 29053
rect 24400 29044 24452 29096
rect 24676 29112 24728 29164
rect 24952 29155 25004 29164
rect 24952 29121 24961 29155
rect 24961 29121 24995 29155
rect 24995 29121 25004 29155
rect 27436 29180 27488 29232
rect 28724 29257 28733 29291
rect 28733 29257 28767 29291
rect 28767 29257 28776 29291
rect 28724 29248 28776 29257
rect 28816 29248 28868 29300
rect 46848 29248 46900 29300
rect 24952 29112 25004 29121
rect 26332 29112 26384 29164
rect 27068 29112 27120 29164
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27528 29153 27580 29164
rect 27528 29119 27537 29153
rect 27537 29119 27571 29153
rect 27571 29119 27580 29153
rect 27988 29155 28040 29164
rect 27528 29112 27580 29119
rect 27988 29121 27997 29155
rect 27997 29121 28031 29155
rect 28031 29121 28040 29155
rect 27988 29112 28040 29121
rect 24768 29044 24820 29096
rect 26240 28976 26292 29028
rect 28264 29155 28316 29164
rect 28264 29121 28273 29155
rect 28273 29121 28307 29155
rect 28307 29121 28316 29155
rect 28264 29112 28316 29121
rect 29000 29112 29052 29164
rect 30564 29223 30616 29232
rect 30564 29189 30573 29223
rect 30573 29189 30607 29223
rect 30607 29189 30616 29223
rect 30564 29180 30616 29189
rect 28356 29087 28408 29096
rect 28356 29053 28365 29087
rect 28365 29053 28399 29087
rect 28399 29053 28408 29087
rect 28356 29044 28408 29053
rect 28816 29044 28868 29096
rect 10416 28951 10468 28960
rect 10416 28917 10425 28951
rect 10425 28917 10459 28951
rect 10459 28917 10468 28951
rect 10416 28908 10468 28917
rect 15292 28908 15344 28960
rect 17408 28908 17460 28960
rect 22376 28951 22428 28960
rect 22376 28917 22385 28951
rect 22385 28917 22419 28951
rect 22419 28917 22428 28951
rect 22376 28908 22428 28917
rect 24400 28908 24452 28960
rect 25688 28908 25740 28960
rect 28816 28908 28868 28960
rect 28908 28908 28960 28960
rect 30472 28976 30524 29028
rect 30932 29112 30984 29164
rect 32680 29155 32732 29164
rect 32680 29121 32689 29155
rect 32689 29121 32723 29155
rect 32723 29121 32732 29155
rect 32680 29112 32732 29121
rect 34796 29112 34848 29164
rect 30748 29087 30800 29096
rect 30748 29053 30757 29087
rect 30757 29053 30791 29087
rect 30791 29053 30800 29087
rect 30748 29044 30800 29053
rect 33048 29044 33100 29096
rect 34612 29044 34664 29096
rect 35348 29112 35400 29164
rect 38016 29180 38068 29232
rect 38476 29223 38528 29232
rect 38476 29189 38485 29223
rect 38485 29189 38519 29223
rect 38519 29189 38528 29223
rect 38476 29180 38528 29189
rect 37464 29155 37516 29164
rect 37464 29121 37471 29155
rect 37471 29121 37516 29155
rect 37464 29112 37516 29121
rect 35716 29087 35768 29096
rect 35716 29053 35725 29087
rect 35725 29053 35759 29087
rect 35759 29053 35768 29087
rect 35716 29044 35768 29053
rect 35808 29044 35860 29096
rect 37648 29155 37700 29164
rect 37648 29121 37657 29155
rect 37657 29121 37691 29155
rect 37691 29121 37700 29155
rect 37648 29112 37700 29121
rect 37832 29112 37884 29164
rect 34796 28976 34848 29028
rect 37280 28976 37332 29028
rect 37740 28976 37792 29028
rect 37924 29019 37976 29028
rect 37924 28985 37933 29019
rect 37933 28985 37967 29019
rect 37967 28985 37976 29019
rect 37924 28976 37976 28985
rect 30840 28951 30892 28960
rect 30840 28917 30849 28951
rect 30849 28917 30883 28951
rect 30883 28917 30892 28951
rect 30840 28908 30892 28917
rect 32404 28908 32456 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 12164 28747 12216 28756
rect 9496 28611 9548 28620
rect 9496 28577 9505 28611
rect 9505 28577 9539 28611
rect 9539 28577 9548 28611
rect 9496 28568 9548 28577
rect 12164 28713 12173 28747
rect 12173 28713 12207 28747
rect 12207 28713 12216 28747
rect 12164 28704 12216 28713
rect 13176 28704 13228 28756
rect 15476 28704 15528 28756
rect 17316 28704 17368 28756
rect 23664 28704 23716 28756
rect 24676 28704 24728 28756
rect 24952 28704 25004 28756
rect 28540 28704 28592 28756
rect 30840 28747 30892 28756
rect 30840 28713 30849 28747
rect 30849 28713 30883 28747
rect 30883 28713 30892 28747
rect 30840 28704 30892 28713
rect 31024 28747 31076 28756
rect 31024 28713 31033 28747
rect 31033 28713 31067 28747
rect 31067 28713 31076 28747
rect 31024 28704 31076 28713
rect 32404 28747 32456 28756
rect 32404 28713 32413 28747
rect 32413 28713 32447 28747
rect 32447 28713 32456 28747
rect 32404 28704 32456 28713
rect 33508 28704 33560 28756
rect 33784 28747 33836 28756
rect 33784 28713 33793 28747
rect 33793 28713 33827 28747
rect 33827 28713 33836 28747
rect 33784 28704 33836 28713
rect 35992 28704 36044 28756
rect 17408 28679 17460 28688
rect 17408 28645 17417 28679
rect 17417 28645 17451 28679
rect 17451 28645 17460 28679
rect 17408 28636 17460 28645
rect 17776 28636 17828 28688
rect 10416 28611 10468 28620
rect 10416 28577 10425 28611
rect 10425 28577 10459 28611
rect 10459 28577 10468 28611
rect 10416 28568 10468 28577
rect 14556 28568 14608 28620
rect 15292 28568 15344 28620
rect 17224 28568 17276 28620
rect 17316 28568 17368 28620
rect 9588 28543 9640 28552
rect 9588 28509 9597 28543
rect 9597 28509 9631 28543
rect 9631 28509 9640 28543
rect 9588 28500 9640 28509
rect 12624 28543 12676 28552
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 12624 28500 12676 28509
rect 13452 28500 13504 28552
rect 17960 28500 18012 28552
rect 11428 28432 11480 28484
rect 15936 28432 15988 28484
rect 16948 28432 17000 28484
rect 20352 28475 20404 28484
rect 20352 28441 20361 28475
rect 20361 28441 20395 28475
rect 20395 28441 20404 28475
rect 20352 28432 20404 28441
rect 22008 28475 22060 28484
rect 22008 28441 22017 28475
rect 22017 28441 22051 28475
rect 22051 28441 22060 28475
rect 22008 28432 22060 28441
rect 23480 28636 23532 28688
rect 24216 28636 24268 28688
rect 23756 28568 23808 28620
rect 25136 28636 25188 28688
rect 35716 28636 35768 28688
rect 46112 28636 46164 28688
rect 24952 28568 25004 28620
rect 26240 28568 26292 28620
rect 23480 28432 23532 28484
rect 24400 28543 24452 28552
rect 24400 28509 24409 28543
rect 24409 28509 24443 28543
rect 24443 28509 24452 28543
rect 25228 28543 25280 28552
rect 24400 28500 24452 28509
rect 25228 28509 25237 28543
rect 25237 28509 25271 28543
rect 25271 28509 25280 28543
rect 25228 28500 25280 28509
rect 26608 28500 26660 28552
rect 27804 28568 27856 28620
rect 28816 28568 28868 28620
rect 30748 28611 30800 28620
rect 27712 28500 27764 28552
rect 29644 28543 29696 28552
rect 29644 28509 29653 28543
rect 29653 28509 29687 28543
rect 29687 28509 29696 28543
rect 29644 28500 29696 28509
rect 30748 28577 30757 28611
rect 30757 28577 30791 28611
rect 30791 28577 30800 28611
rect 30748 28568 30800 28577
rect 31484 28568 31536 28620
rect 30472 28500 30524 28552
rect 32956 28568 33008 28620
rect 31852 28543 31904 28552
rect 25504 28475 25556 28484
rect 25504 28441 25513 28475
rect 25513 28441 25547 28475
rect 25547 28441 25556 28475
rect 25504 28432 25556 28441
rect 27528 28432 27580 28484
rect 29184 28432 29236 28484
rect 30196 28432 30248 28484
rect 31852 28509 31861 28543
rect 31861 28509 31895 28543
rect 31895 28509 31904 28543
rect 31852 28500 31904 28509
rect 31944 28543 31996 28552
rect 31944 28509 31953 28543
rect 31953 28509 31987 28543
rect 31987 28509 31996 28543
rect 31944 28500 31996 28509
rect 32128 28500 32180 28552
rect 32680 28500 32732 28552
rect 33048 28543 33100 28552
rect 33048 28509 33057 28543
rect 33057 28509 33091 28543
rect 33091 28509 33100 28543
rect 33048 28500 33100 28509
rect 36176 28568 36228 28620
rect 36544 28568 36596 28620
rect 38292 28568 38344 28620
rect 46940 28568 46992 28620
rect 35348 28543 35400 28552
rect 35348 28509 35357 28543
rect 35357 28509 35391 28543
rect 35391 28509 35400 28543
rect 35348 28500 35400 28509
rect 39028 28500 39080 28552
rect 46296 28543 46348 28552
rect 46296 28509 46305 28543
rect 46305 28509 46339 28543
rect 46339 28509 46348 28543
rect 46296 28500 46348 28509
rect 30932 28432 30984 28484
rect 33508 28432 33560 28484
rect 36452 28432 36504 28484
rect 13452 28407 13504 28416
rect 13452 28373 13461 28407
rect 13461 28373 13495 28407
rect 13495 28373 13504 28407
rect 13452 28364 13504 28373
rect 17408 28364 17460 28416
rect 22100 28364 22152 28416
rect 23848 28407 23900 28416
rect 23848 28373 23857 28407
rect 23857 28373 23891 28407
rect 23891 28373 23900 28407
rect 23848 28364 23900 28373
rect 28356 28364 28408 28416
rect 31852 28364 31904 28416
rect 31944 28364 31996 28416
rect 35348 28407 35400 28416
rect 35348 28373 35357 28407
rect 35357 28373 35391 28407
rect 35391 28373 35400 28407
rect 35348 28364 35400 28373
rect 36084 28364 36136 28416
rect 36268 28407 36320 28416
rect 36268 28373 36277 28407
rect 36277 28373 36311 28407
rect 36311 28373 36320 28407
rect 36268 28364 36320 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 16304 28160 16356 28212
rect 16856 28160 16908 28212
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 20352 28160 20404 28212
rect 9680 28092 9732 28144
rect 12900 28092 12952 28144
rect 13452 28092 13504 28144
rect 16948 28135 17000 28144
rect 11428 28024 11480 28076
rect 16948 28101 16957 28135
rect 16957 28101 16991 28135
rect 16991 28101 17000 28135
rect 16948 28092 17000 28101
rect 17960 28092 18012 28144
rect 19340 28092 19392 28144
rect 19432 28024 19484 28076
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 25228 28160 25280 28212
rect 25504 28160 25556 28212
rect 22100 28135 22152 28144
rect 22100 28101 22109 28135
rect 22109 28101 22143 28135
rect 22143 28101 22152 28135
rect 22100 28092 22152 28101
rect 22376 28092 22428 28144
rect 23848 28092 23900 28144
rect 23480 28024 23532 28076
rect 8116 27999 8168 28008
rect 8116 27965 8125 27999
rect 8125 27965 8159 27999
rect 8159 27965 8168 27999
rect 8116 27956 8168 27965
rect 12716 27999 12768 28008
rect 3976 27888 4028 27940
rect 12716 27965 12725 27999
rect 12725 27965 12759 27999
rect 12759 27965 12768 27999
rect 12716 27956 12768 27965
rect 12900 27999 12952 28008
rect 12900 27965 12909 27999
rect 12909 27965 12943 27999
rect 12943 27965 12952 27999
rect 12900 27956 12952 27965
rect 8300 27820 8352 27872
rect 11152 27820 11204 27872
rect 17040 27820 17092 27872
rect 18052 27956 18104 28008
rect 19248 27956 19300 28008
rect 23572 27999 23624 28008
rect 23572 27965 23581 27999
rect 23581 27965 23615 27999
rect 23615 27965 23624 27999
rect 23572 27956 23624 27965
rect 24308 28067 24360 28076
rect 24308 28033 24317 28067
rect 24317 28033 24351 28067
rect 24351 28033 24360 28067
rect 24492 28067 24544 28076
rect 24308 28024 24360 28033
rect 24492 28033 24501 28067
rect 24501 28033 24535 28067
rect 24535 28033 24544 28067
rect 24492 28024 24544 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 25228 28067 25280 28076
rect 24584 28024 24636 28033
rect 25228 28033 25237 28067
rect 25237 28033 25271 28067
rect 25271 28033 25280 28067
rect 25228 28024 25280 28033
rect 25504 28067 25556 28076
rect 25504 28033 25513 28067
rect 25513 28033 25547 28067
rect 25547 28033 25556 28067
rect 25504 28024 25556 28033
rect 30380 28160 30432 28212
rect 31208 28160 31260 28212
rect 31944 28160 31996 28212
rect 35348 28160 35400 28212
rect 31392 28092 31444 28144
rect 27620 28067 27672 28076
rect 24952 27956 25004 28008
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 29828 28024 29880 28076
rect 29920 28024 29972 28076
rect 31116 28067 31168 28076
rect 26240 27888 26292 27940
rect 29644 27888 29696 27940
rect 18052 27820 18104 27872
rect 29828 27863 29880 27872
rect 29828 27829 29837 27863
rect 29837 27829 29871 27863
rect 29871 27829 29880 27863
rect 29828 27820 29880 27829
rect 31116 28033 31125 28067
rect 31125 28033 31159 28067
rect 31159 28033 31168 28067
rect 31116 28024 31168 28033
rect 31024 27956 31076 28008
rect 32220 28024 32272 28076
rect 32312 28024 32364 28076
rect 35992 28067 36044 28076
rect 35992 28033 36001 28067
rect 36001 28033 36035 28067
rect 36035 28033 36044 28067
rect 35992 28024 36044 28033
rect 36084 28024 36136 28076
rect 37740 28024 37792 28076
rect 46572 28024 46624 28076
rect 47584 28067 47636 28076
rect 47584 28033 47593 28067
rect 47593 28033 47627 28067
rect 47627 28033 47636 28067
rect 47584 28024 47636 28033
rect 31576 27956 31628 28008
rect 35808 27956 35860 28008
rect 36176 27999 36228 28008
rect 36176 27965 36185 27999
rect 36185 27965 36219 27999
rect 36219 27965 36228 27999
rect 36176 27956 36228 27965
rect 36360 27956 36412 28008
rect 33508 27888 33560 27940
rect 36268 27888 36320 27940
rect 31024 27820 31076 27872
rect 31208 27863 31260 27872
rect 31208 27829 31217 27863
rect 31217 27829 31251 27863
rect 31251 27829 31260 27863
rect 31208 27820 31260 27829
rect 31300 27820 31352 27872
rect 33416 27863 33468 27872
rect 33416 27829 33425 27863
rect 33425 27829 33459 27863
rect 33459 27829 33468 27863
rect 33416 27820 33468 27829
rect 36360 27820 36412 27872
rect 38016 27863 38068 27872
rect 38016 27829 38025 27863
rect 38025 27829 38059 27863
rect 38059 27829 38068 27863
rect 38016 27820 38068 27829
rect 47032 27863 47084 27872
rect 47032 27829 47041 27863
rect 47041 27829 47075 27863
rect 47075 27829 47084 27863
rect 47032 27820 47084 27829
rect 47676 27863 47728 27872
rect 47676 27829 47685 27863
rect 47685 27829 47719 27863
rect 47719 27829 47728 27863
rect 47676 27820 47728 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8116 27616 8168 27668
rect 12900 27616 12952 27668
rect 9036 27591 9088 27600
rect 9036 27557 9045 27591
rect 9045 27557 9079 27591
rect 9079 27557 9088 27591
rect 9036 27548 9088 27557
rect 9680 27548 9732 27600
rect 10692 27548 10744 27600
rect 17960 27616 18012 27668
rect 25412 27616 25464 27668
rect 25504 27616 25556 27668
rect 27896 27616 27948 27668
rect 18052 27591 18104 27600
rect 18052 27557 18061 27591
rect 18061 27557 18095 27591
rect 18095 27557 18104 27591
rect 18052 27548 18104 27557
rect 19340 27591 19392 27600
rect 19340 27557 19349 27591
rect 19349 27557 19383 27591
rect 19383 27557 19392 27591
rect 19340 27548 19392 27557
rect 9588 27480 9640 27532
rect 23664 27548 23716 27600
rect 23756 27548 23808 27600
rect 24676 27548 24728 27600
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 7564 27412 7616 27421
rect 8852 27412 8904 27464
rect 10048 27412 10100 27464
rect 11152 27455 11204 27464
rect 11152 27421 11161 27455
rect 11161 27421 11195 27455
rect 11195 27421 11204 27455
rect 11152 27412 11204 27421
rect 12624 27412 12676 27464
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 19156 27412 19208 27464
rect 24492 27480 24544 27532
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 24768 27455 24820 27464
rect 23664 27412 23716 27421
rect 24768 27421 24777 27455
rect 24777 27421 24811 27455
rect 24811 27421 24820 27455
rect 24768 27412 24820 27421
rect 26332 27412 26384 27464
rect 31024 27616 31076 27668
rect 36360 27659 36412 27668
rect 36360 27625 36390 27659
rect 36390 27625 36412 27659
rect 36360 27616 36412 27625
rect 31392 27591 31444 27600
rect 31392 27557 31401 27591
rect 31401 27557 31435 27591
rect 31435 27557 31444 27591
rect 31392 27548 31444 27557
rect 31484 27548 31536 27600
rect 34796 27548 34848 27600
rect 41420 27548 41472 27600
rect 42064 27548 42116 27600
rect 31576 27480 31628 27532
rect 32220 27523 32272 27532
rect 32220 27489 32229 27523
rect 32229 27489 32263 27523
rect 32263 27489 32272 27523
rect 32220 27480 32272 27489
rect 32588 27412 32640 27464
rect 33784 27480 33836 27532
rect 36452 27480 36504 27532
rect 47032 27480 47084 27532
rect 48136 27523 48188 27532
rect 48136 27489 48145 27523
rect 48145 27489 48179 27523
rect 48179 27489 48188 27523
rect 48136 27480 48188 27489
rect 8208 27319 8260 27328
rect 8208 27285 8217 27319
rect 8217 27285 8251 27319
rect 8251 27285 8260 27319
rect 8208 27276 8260 27285
rect 9220 27276 9272 27328
rect 24308 27344 24360 27396
rect 29920 27387 29972 27396
rect 29920 27353 29929 27387
rect 29929 27353 29963 27387
rect 29963 27353 29972 27387
rect 29920 27344 29972 27353
rect 32036 27344 32088 27396
rect 10232 27276 10284 27328
rect 11244 27276 11296 27328
rect 11520 27276 11572 27328
rect 26424 27276 26476 27328
rect 30196 27276 30248 27328
rect 33968 27412 34020 27464
rect 37740 27412 37792 27464
rect 35440 27344 35492 27396
rect 38016 27344 38068 27396
rect 47676 27344 47728 27396
rect 33324 27276 33376 27328
rect 33692 27276 33744 27328
rect 38384 27319 38436 27328
rect 38384 27285 38393 27319
rect 38393 27285 38427 27319
rect 38427 27285 38436 27319
rect 38384 27276 38436 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 7564 27072 7616 27124
rect 8024 27072 8076 27124
rect 12532 27072 12584 27124
rect 12716 27072 12768 27124
rect 27896 27115 27948 27124
rect 27896 27081 27905 27115
rect 27905 27081 27939 27115
rect 27939 27081 27948 27115
rect 27896 27072 27948 27081
rect 31300 27072 31352 27124
rect 9036 27004 9088 27056
rect 8208 26936 8260 26988
rect 9128 26936 9180 26988
rect 8300 26800 8352 26852
rect 9220 26800 9272 26852
rect 10232 26936 10284 26988
rect 12256 27004 12308 27056
rect 13084 27004 13136 27056
rect 11520 26979 11572 26988
rect 11520 26945 11529 26979
rect 11529 26945 11563 26979
rect 11563 26945 11572 26979
rect 11520 26936 11572 26945
rect 18144 27004 18196 27056
rect 23572 27004 23624 27056
rect 30196 27047 30248 27056
rect 10048 26911 10100 26920
rect 10048 26877 10057 26911
rect 10057 26877 10091 26911
rect 10091 26877 10100 26911
rect 10048 26868 10100 26877
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 12532 26868 12584 26920
rect 17592 26936 17644 26988
rect 17684 26936 17736 26988
rect 17040 26868 17092 26920
rect 22560 26979 22612 26988
rect 22560 26945 22569 26979
rect 22569 26945 22603 26979
rect 22603 26945 22612 26979
rect 22560 26936 22612 26945
rect 23480 26979 23532 26988
rect 23480 26945 23489 26979
rect 23489 26945 23523 26979
rect 23523 26945 23532 26979
rect 23480 26936 23532 26945
rect 24124 26979 24176 26988
rect 24124 26945 24133 26979
rect 24133 26945 24167 26979
rect 24167 26945 24176 26979
rect 24124 26936 24176 26945
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 27160 26979 27212 26988
rect 27160 26945 27169 26979
rect 27169 26945 27203 26979
rect 27203 26945 27212 26979
rect 27160 26936 27212 26945
rect 27804 26936 27856 26988
rect 20260 26868 20312 26920
rect 21088 26868 21140 26920
rect 23112 26868 23164 26920
rect 23664 26868 23716 26920
rect 29184 26911 29236 26920
rect 29184 26877 29193 26911
rect 29193 26877 29227 26911
rect 29227 26877 29236 26911
rect 29184 26868 29236 26877
rect 30196 27013 30205 27047
rect 30205 27013 30239 27047
rect 30239 27013 30248 27047
rect 30196 27004 30248 27013
rect 30380 27047 30432 27056
rect 30380 27013 30389 27047
rect 30389 27013 30423 27047
rect 30423 27013 30432 27047
rect 30380 27004 30432 27013
rect 33416 27072 33468 27124
rect 33784 27004 33836 27056
rect 29644 26979 29696 26988
rect 29644 26945 29653 26979
rect 29653 26945 29687 26979
rect 29687 26945 29696 26979
rect 29644 26936 29696 26945
rect 33876 26936 33928 26988
rect 38292 26936 38344 26988
rect 44272 26936 44324 26988
rect 31944 26868 31996 26920
rect 7380 26732 7432 26784
rect 8208 26732 8260 26784
rect 8576 26775 8628 26784
rect 8576 26741 8585 26775
rect 8585 26741 8619 26775
rect 8619 26741 8628 26775
rect 8576 26732 8628 26741
rect 9496 26775 9548 26784
rect 9496 26741 9505 26775
rect 9505 26741 9539 26775
rect 9539 26741 9548 26775
rect 9496 26732 9548 26741
rect 17868 26800 17920 26852
rect 32128 26800 32180 26852
rect 12348 26732 12400 26784
rect 15016 26775 15068 26784
rect 15016 26741 15025 26775
rect 15025 26741 15059 26775
rect 15059 26741 15068 26775
rect 15016 26732 15068 26741
rect 19432 26732 19484 26784
rect 22652 26732 22704 26784
rect 22744 26775 22796 26784
rect 22744 26741 22753 26775
rect 22753 26741 22787 26775
rect 22787 26741 22796 26775
rect 23572 26775 23624 26784
rect 22744 26732 22796 26741
rect 23572 26741 23581 26775
rect 23581 26741 23615 26775
rect 23615 26741 23624 26775
rect 23572 26732 23624 26741
rect 24308 26775 24360 26784
rect 24308 26741 24317 26775
rect 24317 26741 24351 26775
rect 24351 26741 24360 26775
rect 24308 26732 24360 26741
rect 25964 26732 26016 26784
rect 29000 26732 29052 26784
rect 32588 26868 32640 26920
rect 33600 26800 33652 26852
rect 37740 26800 37792 26852
rect 33048 26732 33100 26784
rect 34796 26775 34848 26784
rect 34796 26741 34805 26775
rect 34805 26741 34839 26775
rect 34839 26741 34848 26775
rect 34796 26732 34848 26741
rect 38660 26732 38712 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8392 26528 8444 26580
rect 9496 26528 9548 26580
rect 12256 26571 12308 26580
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 12348 26528 12400 26580
rect 17592 26528 17644 26580
rect 22560 26528 22612 26580
rect 22836 26528 22888 26580
rect 24308 26528 24360 26580
rect 9036 26460 9088 26512
rect 7380 26367 7432 26376
rect 7380 26333 7389 26367
rect 7389 26333 7423 26367
rect 7423 26333 7432 26367
rect 7380 26324 7432 26333
rect 8576 26392 8628 26444
rect 15844 26460 15896 26512
rect 8392 26324 8444 26376
rect 9496 26324 9548 26376
rect 12716 26392 12768 26444
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 16488 26435 16540 26444
rect 16488 26401 16497 26435
rect 16497 26401 16531 26435
rect 16531 26401 16540 26435
rect 16488 26392 16540 26401
rect 12532 26324 12584 26376
rect 12900 26324 12952 26376
rect 8944 26299 8996 26308
rect 8944 26265 8971 26299
rect 8971 26265 8996 26299
rect 9128 26299 9180 26308
rect 8944 26256 8996 26265
rect 9128 26265 9137 26299
rect 9137 26265 9171 26299
rect 9171 26265 9180 26299
rect 9128 26256 9180 26265
rect 12992 26256 13044 26308
rect 13912 26324 13964 26376
rect 14464 26324 14516 26376
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 15752 26256 15804 26308
rect 19248 26435 19300 26444
rect 19248 26401 19257 26435
rect 19257 26401 19291 26435
rect 19291 26401 19300 26435
rect 19248 26392 19300 26401
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 22376 26392 22428 26444
rect 27252 26392 27304 26444
rect 31024 26392 31076 26444
rect 17868 26324 17920 26376
rect 25412 26324 25464 26376
rect 18144 26256 18196 26308
rect 21180 26256 21232 26308
rect 21824 26299 21876 26308
rect 21824 26265 21833 26299
rect 21833 26265 21867 26299
rect 21867 26265 21876 26299
rect 21824 26256 21876 26265
rect 22100 26256 22152 26308
rect 24952 26256 25004 26308
rect 25964 26299 26016 26308
rect 25964 26265 25973 26299
rect 25973 26265 26007 26299
rect 26007 26265 26016 26299
rect 25964 26256 26016 26265
rect 26424 26256 26476 26308
rect 29828 26299 29880 26308
rect 29828 26265 29837 26299
rect 29837 26265 29871 26299
rect 29871 26265 29880 26299
rect 29828 26256 29880 26265
rect 30380 26256 30432 26308
rect 31760 26528 31812 26580
rect 33600 26528 33652 26580
rect 33784 26571 33836 26580
rect 33784 26537 33793 26571
rect 33793 26537 33827 26571
rect 33827 26537 33836 26571
rect 33784 26528 33836 26537
rect 31944 26460 31996 26512
rect 47860 26528 47912 26580
rect 36176 26460 36228 26512
rect 32588 26392 32640 26444
rect 33048 26392 33100 26444
rect 37832 26392 37884 26444
rect 40224 26392 40276 26444
rect 31944 26324 31996 26376
rect 33692 26367 33744 26376
rect 33692 26333 33701 26367
rect 33701 26333 33735 26367
rect 33735 26333 33744 26367
rect 33692 26324 33744 26333
rect 34888 26367 34940 26376
rect 34888 26333 34897 26367
rect 34897 26333 34931 26367
rect 34931 26333 34940 26367
rect 34888 26324 34940 26333
rect 41420 26324 41472 26376
rect 45192 26324 45244 26376
rect 31760 26256 31812 26308
rect 37832 26299 37884 26308
rect 37832 26265 37841 26299
rect 37841 26265 37875 26299
rect 37875 26265 37884 26299
rect 37832 26256 37884 26265
rect 38384 26256 38436 26308
rect 43996 26256 44048 26308
rect 46848 26256 46900 26308
rect 7840 26231 7892 26240
rect 7840 26197 7849 26231
rect 7849 26197 7883 26231
rect 7883 26197 7892 26231
rect 7840 26188 7892 26197
rect 8300 26188 8352 26240
rect 9220 26188 9272 26240
rect 9772 26188 9824 26240
rect 11704 26188 11756 26240
rect 13268 26231 13320 26240
rect 13268 26197 13277 26231
rect 13277 26197 13311 26231
rect 13311 26197 13320 26231
rect 13268 26188 13320 26197
rect 26792 26188 26844 26240
rect 38752 26188 38804 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 11796 25984 11848 26036
rect 12900 25984 12952 26036
rect 13268 25984 13320 26036
rect 15752 26027 15804 26036
rect 15752 25993 15761 26027
rect 15761 25993 15795 26027
rect 15795 25993 15804 26027
rect 15752 25984 15804 25993
rect 7840 25916 7892 25968
rect 9036 25916 9088 25968
rect 12716 25916 12768 25968
rect 16856 25916 16908 25968
rect 17868 25984 17920 26036
rect 19616 25959 19668 25968
rect 19616 25925 19625 25959
rect 19625 25925 19659 25959
rect 19659 25925 19668 25959
rect 19616 25916 19668 25925
rect 7104 25848 7156 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 12440 25891 12492 25900
rect 12440 25857 12449 25891
rect 12449 25857 12483 25891
rect 12483 25857 12492 25891
rect 12440 25848 12492 25857
rect 12808 25848 12860 25900
rect 12992 25848 13044 25900
rect 14464 25848 14516 25900
rect 15016 25848 15068 25900
rect 15752 25848 15804 25900
rect 21916 25984 21968 26036
rect 23940 25984 23992 26036
rect 27160 25984 27212 26036
rect 27988 25984 28040 26036
rect 29552 25984 29604 26036
rect 29828 25984 29880 26036
rect 21088 25891 21140 25900
rect 11244 25780 11296 25832
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 22284 25959 22336 25968
rect 22284 25925 22293 25959
rect 22293 25925 22327 25959
rect 22327 25925 22336 25959
rect 22284 25916 22336 25925
rect 23572 25916 23624 25968
rect 22560 25848 22612 25900
rect 24032 25848 24084 25900
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 27804 25916 27856 25968
rect 28724 25916 28776 25968
rect 30196 25984 30248 26036
rect 30380 25984 30432 26036
rect 25136 25848 25188 25900
rect 25780 25891 25832 25900
rect 25780 25857 25789 25891
rect 25789 25857 25823 25891
rect 25823 25857 25832 25891
rect 25780 25848 25832 25857
rect 27344 25891 27396 25900
rect 17132 25780 17184 25832
rect 17776 25823 17828 25832
rect 17776 25789 17785 25823
rect 17785 25789 17819 25823
rect 17819 25789 17828 25823
rect 17776 25780 17828 25789
rect 17960 25823 18012 25832
rect 17960 25789 17969 25823
rect 17969 25789 18003 25823
rect 18003 25789 18012 25823
rect 17960 25780 18012 25789
rect 24124 25780 24176 25832
rect 27344 25857 27353 25891
rect 27353 25857 27387 25891
rect 27387 25857 27396 25891
rect 27344 25848 27396 25857
rect 18144 25712 18196 25764
rect 27160 25780 27212 25832
rect 29000 25848 29052 25900
rect 29460 25891 29512 25900
rect 29460 25857 29469 25891
rect 29469 25857 29503 25891
rect 29503 25857 29512 25891
rect 29460 25848 29512 25857
rect 29644 25848 29696 25900
rect 31944 25848 31996 25900
rect 31024 25780 31076 25832
rect 31300 25823 31352 25832
rect 31300 25789 31309 25823
rect 31309 25789 31343 25823
rect 31343 25789 31352 25823
rect 31300 25780 31352 25789
rect 32588 25916 32640 25968
rect 36176 25984 36228 26036
rect 37832 25984 37884 26036
rect 33508 25959 33560 25968
rect 33508 25925 33517 25959
rect 33517 25925 33551 25959
rect 33551 25925 33560 25959
rect 33508 25916 33560 25925
rect 34796 25916 34848 25968
rect 33692 25848 33744 25900
rect 37740 25891 37792 25900
rect 37740 25857 37749 25891
rect 37749 25857 37783 25891
rect 37783 25857 37792 25891
rect 37740 25848 37792 25857
rect 40408 25916 40460 25968
rect 41052 25959 41104 25968
rect 41052 25925 41061 25959
rect 41061 25925 41095 25959
rect 41095 25925 41104 25959
rect 41052 25916 41104 25925
rect 41144 25916 41196 25968
rect 45652 25916 45704 25968
rect 37924 25891 37976 25900
rect 37924 25857 37933 25891
rect 37933 25857 37967 25891
rect 37967 25857 37976 25891
rect 37924 25848 37976 25857
rect 9220 25644 9272 25696
rect 12072 25644 12124 25696
rect 14832 25687 14884 25696
rect 14832 25653 14841 25687
rect 14841 25653 14875 25687
rect 14875 25653 14884 25687
rect 14832 25644 14884 25653
rect 17040 25687 17092 25696
rect 17040 25653 17049 25687
rect 17049 25653 17083 25687
rect 17083 25653 17092 25687
rect 17040 25644 17092 25653
rect 21824 25644 21876 25696
rect 22192 25644 22244 25696
rect 25964 25644 26016 25696
rect 27344 25644 27396 25696
rect 28080 25687 28132 25696
rect 28080 25653 28089 25687
rect 28089 25653 28123 25687
rect 28123 25653 28132 25687
rect 28080 25644 28132 25653
rect 32404 25644 32456 25696
rect 33048 25644 33100 25696
rect 34520 25823 34572 25832
rect 34520 25789 34529 25823
rect 34529 25789 34563 25823
rect 34563 25789 34572 25823
rect 34520 25780 34572 25789
rect 38200 25848 38252 25900
rect 38752 25891 38804 25900
rect 38752 25857 38761 25891
rect 38761 25857 38795 25891
rect 38795 25857 38804 25891
rect 38752 25848 38804 25857
rect 40224 25891 40276 25900
rect 40224 25857 40233 25891
rect 40233 25857 40267 25891
rect 40267 25857 40276 25891
rect 40224 25848 40276 25857
rect 45560 25848 45612 25900
rect 33692 25644 33744 25696
rect 35532 25644 35584 25696
rect 38292 25644 38344 25696
rect 46480 25644 46532 25696
rect 47768 25687 47820 25696
rect 47768 25653 47777 25687
rect 47777 25653 47811 25687
rect 47811 25653 47820 25687
rect 47768 25644 47820 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 9036 25483 9088 25492
rect 9036 25449 9045 25483
rect 9045 25449 9079 25483
rect 9079 25449 9088 25483
rect 9036 25440 9088 25449
rect 13268 25440 13320 25492
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 7104 25236 7156 25288
rect 9036 25236 9088 25288
rect 9772 25279 9824 25288
rect 9772 25245 9781 25279
rect 9781 25245 9815 25279
rect 9815 25245 9824 25279
rect 9772 25236 9824 25245
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 22100 25440 22152 25492
rect 23480 25440 23532 25492
rect 23940 25440 23992 25492
rect 20076 25372 20128 25424
rect 22744 25372 22796 25424
rect 23112 25372 23164 25424
rect 24860 25372 24912 25424
rect 13912 25304 13964 25356
rect 13820 25236 13872 25288
rect 14832 25304 14884 25356
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 1768 25168 1820 25220
rect 13084 25168 13136 25220
rect 17132 25236 17184 25288
rect 21732 25304 21784 25356
rect 20996 25236 21048 25288
rect 22836 25279 22888 25288
rect 18144 25168 18196 25220
rect 19340 25168 19392 25220
rect 19432 25168 19484 25220
rect 19708 25211 19760 25220
rect 19708 25177 19717 25211
rect 19717 25177 19751 25211
rect 19751 25177 19760 25211
rect 19708 25168 19760 25177
rect 21272 25168 21324 25220
rect 22008 25211 22060 25220
rect 7564 25100 7616 25152
rect 9588 25143 9640 25152
rect 9588 25109 9597 25143
rect 9597 25109 9631 25143
rect 9631 25109 9640 25143
rect 9588 25100 9640 25109
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 14464 25143 14516 25152
rect 14464 25109 14473 25143
rect 14473 25109 14507 25143
rect 14507 25109 14516 25143
rect 14464 25100 14516 25109
rect 15108 25100 15160 25152
rect 22008 25177 22017 25211
rect 22017 25177 22051 25211
rect 22051 25177 22060 25211
rect 22008 25168 22060 25177
rect 22836 25245 22845 25279
rect 22845 25245 22879 25279
rect 22879 25245 22888 25279
rect 22836 25236 22888 25245
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 26240 25440 26292 25492
rect 26884 25440 26936 25492
rect 27160 25483 27212 25492
rect 27160 25449 27169 25483
rect 27169 25449 27203 25483
rect 27203 25449 27212 25483
rect 27160 25440 27212 25449
rect 28080 25440 28132 25492
rect 29736 25372 29788 25424
rect 32312 25372 32364 25424
rect 33140 25372 33192 25424
rect 34520 25440 34572 25492
rect 37924 25440 37976 25492
rect 41144 25372 41196 25424
rect 26240 25304 26292 25356
rect 32404 25347 32456 25356
rect 32404 25313 32413 25347
rect 32413 25313 32447 25347
rect 32447 25313 32456 25347
rect 32404 25304 32456 25313
rect 32496 25347 32548 25356
rect 32496 25313 32505 25347
rect 32505 25313 32539 25347
rect 32539 25313 32548 25347
rect 32496 25304 32548 25313
rect 33692 25304 33744 25356
rect 26792 25279 26844 25288
rect 26792 25245 26801 25279
rect 26801 25245 26835 25279
rect 26835 25245 26844 25279
rect 26792 25236 26844 25245
rect 30104 25236 30156 25288
rect 31944 25236 31996 25288
rect 32956 25236 33008 25288
rect 34060 25279 34112 25288
rect 22744 25168 22796 25220
rect 24308 25168 24360 25220
rect 28632 25168 28684 25220
rect 34060 25245 34069 25279
rect 34069 25245 34103 25279
rect 34103 25245 34112 25279
rect 34060 25236 34112 25245
rect 35532 25304 35584 25356
rect 35440 25236 35492 25288
rect 37464 25304 37516 25356
rect 38292 25304 38344 25356
rect 40316 25304 40368 25356
rect 40776 25347 40828 25356
rect 40776 25313 40785 25347
rect 40785 25313 40819 25347
rect 40819 25313 40828 25347
rect 40776 25304 40828 25313
rect 45744 25304 45796 25356
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 48136 25347 48188 25356
rect 48136 25313 48145 25347
rect 48145 25313 48179 25347
rect 48179 25313 48188 25347
rect 48136 25304 48188 25313
rect 37096 25236 37148 25288
rect 38016 25236 38068 25288
rect 40224 25279 40276 25288
rect 40224 25245 40233 25279
rect 40233 25245 40267 25279
rect 40267 25245 40276 25279
rect 40224 25236 40276 25245
rect 46296 25279 46348 25288
rect 46296 25245 46305 25279
rect 46305 25245 46339 25279
rect 46339 25245 46348 25279
rect 46296 25236 46348 25245
rect 23480 25100 23532 25152
rect 35808 25168 35860 25220
rect 36084 25168 36136 25220
rect 38660 25100 38712 25152
rect 45652 25100 45704 25152
rect 46112 25100 46164 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 12440 24896 12492 24948
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 8944 24760 8996 24812
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 9588 24692 9640 24744
rect 9036 24624 9088 24676
rect 12716 24735 12768 24744
rect 12716 24701 12725 24735
rect 12725 24701 12759 24735
rect 12759 24701 12768 24735
rect 13636 24760 13688 24812
rect 14464 24828 14516 24880
rect 17408 24896 17460 24948
rect 19432 24896 19484 24948
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 15752 24803 15804 24812
rect 13820 24760 13872 24769
rect 15752 24769 15761 24803
rect 15761 24769 15795 24803
rect 15795 24769 15804 24803
rect 15752 24760 15804 24769
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 17868 24760 17920 24812
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 22008 24760 22060 24812
rect 23296 24896 23348 24948
rect 24032 24896 24084 24948
rect 24860 24896 24912 24948
rect 29460 24896 29512 24948
rect 30288 24896 30340 24948
rect 25136 24828 25188 24880
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 23480 24803 23532 24812
rect 22652 24760 22704 24769
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 12716 24692 12768 24701
rect 12532 24624 12584 24676
rect 14096 24692 14148 24744
rect 22100 24692 22152 24744
rect 22192 24692 22244 24744
rect 22468 24735 22520 24744
rect 22468 24701 22477 24735
rect 22477 24701 22511 24735
rect 22511 24701 22520 24735
rect 23940 24760 23992 24812
rect 22468 24692 22520 24701
rect 8852 24556 8904 24608
rect 9956 24556 10008 24608
rect 11612 24599 11664 24608
rect 11612 24565 11621 24599
rect 11621 24565 11655 24599
rect 11655 24565 11664 24599
rect 11612 24556 11664 24565
rect 12900 24556 12952 24608
rect 20352 24624 20404 24676
rect 13820 24556 13872 24608
rect 16856 24556 16908 24608
rect 17500 24556 17552 24608
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 22284 24556 22336 24608
rect 25872 24760 25924 24812
rect 26332 24760 26384 24812
rect 27620 24760 27672 24812
rect 28632 24803 28684 24812
rect 28632 24769 28641 24803
rect 28641 24769 28675 24803
rect 28675 24769 28684 24803
rect 28632 24760 28684 24769
rect 26240 24692 26292 24744
rect 27252 24735 27304 24744
rect 27252 24701 27261 24735
rect 27261 24701 27295 24735
rect 27295 24701 27304 24735
rect 27252 24692 27304 24701
rect 27528 24692 27580 24744
rect 24676 24624 24728 24676
rect 30104 24760 30156 24812
rect 30196 24692 30248 24744
rect 30472 24760 30524 24812
rect 32496 24896 32548 24948
rect 33508 24939 33560 24948
rect 33508 24905 33517 24939
rect 33517 24905 33551 24939
rect 33551 24905 33560 24939
rect 33508 24896 33560 24905
rect 34060 24896 34112 24948
rect 31300 24828 31352 24880
rect 32864 24760 32916 24812
rect 33140 24803 33192 24812
rect 33140 24769 33149 24803
rect 33149 24769 33183 24803
rect 33183 24769 33192 24803
rect 33140 24760 33192 24769
rect 31760 24692 31812 24744
rect 31944 24692 31996 24744
rect 32312 24692 32364 24744
rect 33692 24760 33744 24812
rect 34704 24760 34756 24812
rect 38016 24828 38068 24880
rect 37280 24803 37332 24812
rect 37280 24769 37289 24803
rect 37289 24769 37323 24803
rect 37323 24769 37332 24803
rect 37280 24760 37332 24769
rect 46020 24760 46072 24812
rect 47124 24760 47176 24812
rect 37004 24692 37056 24744
rect 38752 24692 38804 24744
rect 46204 24735 46256 24744
rect 46204 24701 46213 24735
rect 46213 24701 46247 24735
rect 46247 24701 46256 24735
rect 46204 24692 46256 24701
rect 29920 24624 29972 24676
rect 46756 24624 46808 24676
rect 24952 24556 25004 24608
rect 26148 24556 26200 24608
rect 26332 24599 26384 24608
rect 26332 24565 26341 24599
rect 26341 24565 26375 24599
rect 26375 24565 26384 24599
rect 26332 24556 26384 24565
rect 26516 24556 26568 24608
rect 27988 24556 28040 24608
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 30012 24556 30064 24608
rect 31300 24556 31352 24608
rect 32312 24599 32364 24608
rect 32312 24565 32321 24599
rect 32321 24565 32355 24599
rect 32355 24565 32364 24599
rect 32312 24556 32364 24565
rect 32404 24556 32456 24608
rect 32956 24556 33008 24608
rect 36728 24556 36780 24608
rect 37464 24599 37516 24608
rect 37464 24565 37473 24599
rect 37473 24565 37507 24599
rect 37507 24565 37516 24599
rect 37464 24556 37516 24565
rect 46480 24556 46532 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1676 24284 1728 24336
rect 12900 24352 12952 24404
rect 13084 24352 13136 24404
rect 8944 24284 8996 24336
rect 11796 24284 11848 24336
rect 1952 24216 2004 24268
rect 17960 24284 18012 24336
rect 22008 24352 22060 24404
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 26240 24395 26292 24404
rect 22100 24352 22152 24361
rect 22744 24284 22796 24336
rect 9036 24148 9088 24200
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 12532 24148 12584 24200
rect 18144 24216 18196 24268
rect 22008 24216 22060 24268
rect 26240 24361 26249 24395
rect 26249 24361 26283 24395
rect 26283 24361 26292 24395
rect 26240 24352 26292 24361
rect 28816 24395 28868 24404
rect 28816 24361 28825 24395
rect 28825 24361 28859 24395
rect 28859 24361 28868 24395
rect 28816 24352 28868 24361
rect 26976 24284 27028 24336
rect 30656 24352 30708 24404
rect 31944 24352 31996 24404
rect 35440 24352 35492 24404
rect 37280 24352 37332 24404
rect 38292 24352 38344 24404
rect 30748 24284 30800 24336
rect 24032 24216 24084 24268
rect 25872 24216 25924 24268
rect 10140 24080 10192 24132
rect 11612 24080 11664 24132
rect 17040 24080 17092 24132
rect 17316 24080 17368 24132
rect 9588 24012 9640 24064
rect 12992 24012 13044 24064
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 17592 24012 17644 24064
rect 19984 24012 20036 24064
rect 25964 24191 26016 24200
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 26056 24191 26108 24200
rect 26056 24157 26065 24191
rect 26065 24157 26099 24191
rect 26099 24157 26108 24191
rect 26056 24148 26108 24157
rect 26884 24191 26936 24200
rect 20352 24123 20404 24132
rect 20352 24089 20361 24123
rect 20361 24089 20395 24123
rect 20395 24089 20404 24123
rect 20352 24080 20404 24089
rect 21088 24080 21140 24132
rect 21640 24080 21692 24132
rect 26332 24080 26384 24132
rect 20996 24012 21048 24064
rect 22468 24055 22520 24064
rect 22468 24021 22477 24055
rect 22477 24021 22511 24055
rect 22511 24021 22520 24055
rect 22468 24012 22520 24021
rect 24400 24012 24452 24064
rect 25596 24012 25648 24064
rect 26148 24012 26200 24064
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 26884 24148 26936 24157
rect 29460 24148 29512 24200
rect 30012 24191 30064 24200
rect 30012 24157 30021 24191
rect 30021 24157 30055 24191
rect 30055 24157 30064 24191
rect 30012 24148 30064 24157
rect 30288 24148 30340 24200
rect 32864 24284 32916 24336
rect 31300 24191 31352 24200
rect 31300 24157 31309 24191
rect 31309 24157 31343 24191
rect 31343 24157 31352 24191
rect 31300 24148 31352 24157
rect 32404 24191 32456 24200
rect 32404 24157 32413 24191
rect 32413 24157 32447 24191
rect 32447 24157 32456 24191
rect 32404 24148 32456 24157
rect 32772 24148 32824 24200
rect 37096 24327 37148 24336
rect 37096 24293 37105 24327
rect 37105 24293 37139 24327
rect 37139 24293 37148 24327
rect 37096 24284 37148 24293
rect 47768 24284 47820 24336
rect 29828 24012 29880 24064
rect 30748 24012 30800 24064
rect 31668 24080 31720 24132
rect 31300 24012 31352 24064
rect 32128 24012 32180 24064
rect 33876 24148 33928 24200
rect 33508 24080 33560 24132
rect 35900 24123 35952 24132
rect 35900 24089 35909 24123
rect 35909 24089 35943 24123
rect 35943 24089 35952 24123
rect 35900 24080 35952 24089
rect 36084 24123 36136 24132
rect 36084 24089 36093 24123
rect 36093 24089 36127 24123
rect 36127 24089 36136 24123
rect 36084 24080 36136 24089
rect 36360 24080 36412 24132
rect 36728 24080 36780 24132
rect 36176 24055 36228 24064
rect 36176 24021 36185 24055
rect 36185 24021 36219 24055
rect 36219 24021 36228 24055
rect 36176 24012 36228 24021
rect 36544 24012 36596 24064
rect 37004 24148 37056 24200
rect 46480 24259 46532 24268
rect 46480 24225 46489 24259
rect 46489 24225 46523 24259
rect 46523 24225 46532 24259
rect 46480 24216 46532 24225
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 38568 24148 38620 24200
rect 37740 24080 37792 24132
rect 38200 24080 38252 24132
rect 37924 24012 37976 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 11520 23808 11572 23860
rect 15108 23808 15160 23860
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 8760 23672 8812 23724
rect 9588 23672 9640 23724
rect 12716 23740 12768 23792
rect 14280 23740 14332 23792
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 10968 23468 11020 23520
rect 12256 23672 12308 23724
rect 15016 23672 15068 23724
rect 17500 23672 17552 23724
rect 19984 23740 20036 23792
rect 22744 23740 22796 23792
rect 22468 23715 22520 23724
rect 14464 23604 14516 23656
rect 22468 23681 22477 23715
rect 22477 23681 22511 23715
rect 22511 23681 22520 23715
rect 22468 23672 22520 23681
rect 19248 23604 19300 23656
rect 12348 23468 12400 23520
rect 13820 23468 13872 23520
rect 14372 23468 14424 23520
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 16764 23511 16816 23520
rect 16764 23477 16773 23511
rect 16773 23477 16807 23511
rect 16807 23477 16816 23511
rect 16764 23468 16816 23477
rect 18052 23468 18104 23520
rect 22284 23511 22336 23520
rect 22284 23477 22293 23511
rect 22293 23477 22327 23511
rect 22327 23477 22336 23511
rect 22284 23468 22336 23477
rect 23756 23468 23808 23520
rect 24400 23647 24452 23656
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 26056 23808 26108 23860
rect 26424 23808 26476 23860
rect 26884 23808 26936 23860
rect 25872 23740 25924 23792
rect 26148 23672 26200 23724
rect 26332 23672 26384 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 31116 23808 31168 23860
rect 31300 23851 31352 23860
rect 31300 23817 31309 23851
rect 31309 23817 31343 23851
rect 31343 23817 31352 23851
rect 31300 23808 31352 23817
rect 31852 23808 31904 23860
rect 29828 23783 29880 23792
rect 29828 23749 29837 23783
rect 29837 23749 29871 23783
rect 29871 23749 29880 23783
rect 29828 23740 29880 23749
rect 31208 23740 31260 23792
rect 27528 23672 27580 23724
rect 30196 23604 30248 23656
rect 31852 23672 31904 23724
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32312 23808 32364 23860
rect 32496 23808 32548 23860
rect 34796 23808 34848 23860
rect 35900 23808 35952 23860
rect 31116 23604 31168 23656
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 32864 23672 32916 23724
rect 34704 23715 34756 23724
rect 34704 23681 34713 23715
rect 34713 23681 34747 23715
rect 34747 23681 34756 23715
rect 34704 23672 34756 23681
rect 35440 23715 35492 23724
rect 35440 23681 35449 23715
rect 35449 23681 35483 23715
rect 35483 23681 35492 23715
rect 35440 23672 35492 23681
rect 36176 23740 36228 23792
rect 36360 23715 36412 23724
rect 36360 23681 36369 23715
rect 36369 23681 36403 23715
rect 36403 23681 36412 23715
rect 36360 23672 36412 23681
rect 36544 23715 36596 23724
rect 36544 23681 36553 23715
rect 36553 23681 36587 23715
rect 36587 23681 36596 23715
rect 36544 23672 36596 23681
rect 36728 23715 36780 23724
rect 36728 23681 36737 23715
rect 36737 23681 36771 23715
rect 36771 23681 36780 23715
rect 36728 23672 36780 23681
rect 37556 23715 37608 23724
rect 37556 23681 37565 23715
rect 37565 23681 37599 23715
rect 37599 23681 37608 23715
rect 37556 23672 37608 23681
rect 37924 23715 37976 23724
rect 33876 23604 33928 23656
rect 37280 23647 37332 23656
rect 37280 23613 37289 23647
rect 37289 23613 37323 23647
rect 37323 23613 37332 23647
rect 37280 23604 37332 23613
rect 37924 23681 37933 23715
rect 37933 23681 37967 23715
rect 37967 23681 37976 23715
rect 37924 23672 37976 23681
rect 38568 23715 38620 23724
rect 28816 23536 28868 23588
rect 32220 23536 32272 23588
rect 31760 23468 31812 23520
rect 32404 23468 32456 23520
rect 35716 23511 35768 23520
rect 35716 23477 35725 23511
rect 35725 23477 35759 23511
rect 35759 23477 35768 23511
rect 35716 23468 35768 23477
rect 36360 23536 36412 23588
rect 38568 23681 38577 23715
rect 38577 23681 38611 23715
rect 38611 23681 38620 23715
rect 38568 23672 38620 23681
rect 45192 23715 45244 23724
rect 45192 23681 45201 23715
rect 45201 23681 45235 23715
rect 45235 23681 45244 23715
rect 45192 23672 45244 23681
rect 47584 23715 47636 23724
rect 47584 23681 47593 23715
rect 47593 23681 47627 23715
rect 47627 23681 47636 23715
rect 47584 23672 47636 23681
rect 44088 23604 44140 23656
rect 46572 23604 46624 23656
rect 46848 23647 46900 23656
rect 46848 23613 46857 23647
rect 46857 23613 46891 23647
rect 46891 23613 46900 23647
rect 46848 23604 46900 23613
rect 47952 23536 48004 23588
rect 47676 23511 47728 23520
rect 47676 23477 47685 23511
rect 47685 23477 47719 23511
rect 47719 23477 47728 23511
rect 47676 23468 47728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 14464 23264 14516 23316
rect 19340 23307 19392 23316
rect 19340 23273 19349 23307
rect 19349 23273 19383 23307
rect 19383 23273 19392 23307
rect 19340 23264 19392 23273
rect 23756 23307 23808 23316
rect 23756 23273 23765 23307
rect 23765 23273 23799 23307
rect 23799 23273 23808 23307
rect 23756 23264 23808 23273
rect 26976 23264 27028 23316
rect 28908 23264 28960 23316
rect 30288 23307 30340 23316
rect 30288 23273 30297 23307
rect 30297 23273 30331 23307
rect 30331 23273 30340 23307
rect 30288 23264 30340 23273
rect 31208 23307 31260 23316
rect 31208 23273 31217 23307
rect 31217 23273 31251 23307
rect 31251 23273 31260 23307
rect 31208 23264 31260 23273
rect 31852 23264 31904 23316
rect 36452 23264 36504 23316
rect 38568 23264 38620 23316
rect 20 22992 72 23044
rect 14372 23171 14424 23180
rect 11336 23060 11388 23112
rect 9956 22992 10008 23044
rect 10324 22924 10376 22976
rect 10968 22924 11020 22976
rect 12808 23060 12860 23112
rect 13360 23060 13412 23112
rect 14372 23137 14381 23171
rect 14381 23137 14415 23171
rect 14415 23137 14424 23171
rect 14372 23128 14424 23137
rect 15200 23128 15252 23180
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 22008 23171 22060 23180
rect 22008 23137 22017 23171
rect 22017 23137 22051 23171
rect 22051 23137 22060 23171
rect 22008 23128 22060 23137
rect 22376 23128 22428 23180
rect 25596 23171 25648 23180
rect 25596 23137 25605 23171
rect 25605 23137 25639 23171
rect 25639 23137 25648 23171
rect 25596 23128 25648 23137
rect 26792 23128 26844 23180
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 19984 23060 20036 23112
rect 20536 23060 20588 23112
rect 20720 23060 20772 23112
rect 23388 23060 23440 23112
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 30380 23128 30432 23180
rect 31668 23128 31720 23180
rect 34796 23128 34848 23180
rect 47676 23128 47728 23180
rect 30472 23103 30524 23112
rect 30472 23069 30481 23103
rect 30481 23069 30515 23103
rect 30515 23069 30524 23103
rect 30472 23060 30524 23069
rect 30656 23060 30708 23112
rect 33232 23060 33284 23112
rect 34704 23060 34756 23112
rect 41420 23103 41472 23112
rect 41420 23069 41429 23103
rect 41429 23069 41463 23103
rect 41463 23069 41472 23103
rect 41420 23060 41472 23069
rect 46296 23103 46348 23112
rect 11704 22967 11756 22976
rect 11704 22933 11713 22967
rect 11713 22933 11747 22967
rect 11747 22933 11756 22967
rect 11704 22924 11756 22933
rect 12440 22967 12492 22976
rect 12440 22933 12449 22967
rect 12449 22933 12483 22967
rect 12483 22933 12492 22967
rect 12440 22924 12492 22933
rect 14188 22924 14240 22976
rect 15292 22967 15344 22976
rect 15292 22933 15301 22967
rect 15301 22933 15335 22967
rect 15335 22933 15344 22967
rect 15292 22924 15344 22933
rect 18420 22992 18472 23044
rect 22284 23035 22336 23044
rect 22284 23001 22293 23035
rect 22293 23001 22327 23035
rect 22327 23001 22336 23035
rect 22284 22992 22336 23001
rect 26332 22992 26384 23044
rect 27068 22992 27120 23044
rect 35716 22992 35768 23044
rect 37280 22992 37332 23044
rect 37464 22992 37516 23044
rect 41328 22992 41380 23044
rect 46296 23069 46305 23103
rect 46305 23069 46339 23103
rect 46339 23069 46348 23103
rect 46296 23060 46348 23069
rect 47124 22992 47176 23044
rect 48228 22992 48280 23044
rect 19064 22924 19116 22976
rect 20444 22967 20496 22976
rect 20444 22933 20453 22967
rect 20453 22933 20487 22967
rect 20487 22933 20496 22967
rect 20444 22924 20496 22933
rect 33140 22924 33192 22976
rect 34612 22924 34664 22976
rect 34796 22924 34848 22976
rect 41604 22967 41656 22976
rect 41604 22933 41613 22967
rect 41613 22933 41647 22967
rect 41647 22933 41656 22967
rect 41604 22924 41656 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 8024 22627 8076 22636
rect 8024 22593 8033 22627
rect 8033 22593 8067 22627
rect 8067 22593 8076 22627
rect 8024 22584 8076 22593
rect 13084 22720 13136 22772
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 18420 22763 18472 22772
rect 18420 22729 18429 22763
rect 18429 22729 18463 22763
rect 18463 22729 18472 22763
rect 18420 22720 18472 22729
rect 11704 22652 11756 22704
rect 12440 22652 12492 22704
rect 13360 22652 13412 22704
rect 14188 22627 14240 22636
rect 14188 22593 14197 22627
rect 14197 22593 14231 22627
rect 14231 22593 14240 22627
rect 14188 22584 14240 22593
rect 14740 22584 14792 22636
rect 16856 22652 16908 22704
rect 19064 22652 19116 22704
rect 23388 22695 23440 22704
rect 23388 22661 23397 22695
rect 23397 22661 23431 22695
rect 23431 22661 23440 22695
rect 23388 22652 23440 22661
rect 26332 22695 26384 22704
rect 26332 22661 26341 22695
rect 26341 22661 26375 22695
rect 26375 22661 26384 22695
rect 26332 22652 26384 22661
rect 20536 22627 20588 22636
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 11796 22559 11848 22568
rect 3792 22448 3844 22500
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 16580 22448 16632 22500
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 23112 22584 23164 22636
rect 26148 22584 26200 22636
rect 27620 22652 27672 22704
rect 28172 22652 28224 22704
rect 32404 22695 32456 22704
rect 32404 22661 32413 22695
rect 32413 22661 32447 22695
rect 32447 22661 32456 22695
rect 32404 22652 32456 22661
rect 33140 22652 33192 22704
rect 34612 22652 34664 22704
rect 26792 22516 26844 22568
rect 27068 22627 27120 22636
rect 27068 22593 27077 22627
rect 27077 22593 27111 22627
rect 27111 22593 27120 22627
rect 27068 22584 27120 22593
rect 35440 22584 35492 22636
rect 27712 22516 27764 22568
rect 32128 22559 32180 22568
rect 32128 22525 32137 22559
rect 32137 22525 32171 22559
rect 32171 22525 32180 22559
rect 32128 22516 32180 22525
rect 33876 22559 33928 22568
rect 33876 22525 33885 22559
rect 33885 22525 33919 22559
rect 33919 22525 33928 22559
rect 33876 22516 33928 22525
rect 36452 22652 36504 22704
rect 37464 22652 37516 22704
rect 41420 22652 41472 22704
rect 46020 22652 46072 22704
rect 46572 22720 46624 22772
rect 37280 22627 37332 22636
rect 19708 22448 19760 22500
rect 20904 22448 20956 22500
rect 26884 22448 26936 22500
rect 27344 22448 27396 22500
rect 37280 22593 37289 22627
rect 37289 22593 37323 22627
rect 37323 22593 37332 22627
rect 37280 22584 37332 22593
rect 47584 22627 47636 22636
rect 47584 22593 47593 22627
rect 47593 22593 47627 22627
rect 47627 22593 47636 22627
rect 47584 22584 47636 22593
rect 42432 22559 42484 22568
rect 42432 22525 42441 22559
rect 42441 22525 42475 22559
rect 42475 22525 42484 22559
rect 42432 22516 42484 22525
rect 42616 22559 42668 22568
rect 42616 22525 42625 22559
rect 42625 22525 42659 22559
rect 42659 22525 42668 22559
rect 42616 22516 42668 22525
rect 43996 22559 44048 22568
rect 43996 22525 44005 22559
rect 44005 22525 44039 22559
rect 44039 22525 44048 22559
rect 43996 22516 44048 22525
rect 45652 22559 45704 22568
rect 45652 22525 45661 22559
rect 45661 22525 45695 22559
rect 45695 22525 45704 22559
rect 45652 22516 45704 22525
rect 47860 22516 47912 22568
rect 47400 22448 47452 22500
rect 9128 22380 9180 22432
rect 20168 22380 20220 22432
rect 20812 22380 20864 22432
rect 35348 22380 35400 22432
rect 38200 22380 38252 22432
rect 41328 22380 41380 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8852 22176 8904 22228
rect 15936 22176 15988 22228
rect 20444 22176 20496 22228
rect 20904 22176 20956 22228
rect 38200 22176 38252 22228
rect 42616 22176 42668 22228
rect 46296 22176 46348 22228
rect 12624 22151 12676 22160
rect 12624 22117 12633 22151
rect 12633 22117 12667 22151
rect 12667 22117 12676 22151
rect 12624 22108 12676 22117
rect 17040 22151 17092 22160
rect 17040 22117 17049 22151
rect 17049 22117 17083 22151
rect 17083 22117 17092 22151
rect 17040 22108 17092 22117
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 9128 22083 9180 22092
rect 9128 22049 9137 22083
rect 9137 22049 9171 22083
rect 9171 22049 9180 22083
rect 9128 22040 9180 22049
rect 9312 22040 9364 22092
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11336 21972 11388 21981
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 13268 21972 13320 22024
rect 12992 21904 13044 21956
rect 15292 21972 15344 22024
rect 15568 21972 15620 22024
rect 16672 22040 16724 22092
rect 20812 22040 20864 22092
rect 19708 21972 19760 22024
rect 27988 22151 28040 22160
rect 27988 22117 27997 22151
rect 27997 22117 28031 22151
rect 28031 22117 28040 22151
rect 27988 22108 28040 22117
rect 32772 22151 32824 22160
rect 32772 22117 32781 22151
rect 32781 22117 32815 22151
rect 32815 22117 32824 22151
rect 32772 22108 32824 22117
rect 33232 22108 33284 22160
rect 17224 21904 17276 21956
rect 18604 21904 18656 21956
rect 19340 21904 19392 21956
rect 20812 21904 20864 21956
rect 5448 21836 5500 21888
rect 9312 21836 9364 21888
rect 9588 21836 9640 21888
rect 11980 21836 12032 21888
rect 14464 21836 14516 21888
rect 15752 21836 15804 21888
rect 16948 21836 17000 21888
rect 20444 21836 20496 21888
rect 20536 21836 20588 21888
rect 22652 21904 22704 21956
rect 26608 21972 26660 22024
rect 26976 22040 27028 22092
rect 27712 22015 27764 22024
rect 23112 21904 23164 21956
rect 23388 21904 23440 21956
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 26976 21947 27028 21956
rect 26976 21913 26985 21947
rect 26985 21913 27019 21947
rect 27019 21913 27028 21947
rect 28172 21972 28224 22024
rect 29828 22015 29880 22024
rect 29828 21981 29837 22015
rect 29837 21981 29871 22015
rect 29871 21981 29880 22015
rect 29828 21972 29880 21981
rect 26976 21904 27028 21913
rect 26424 21836 26476 21888
rect 27160 21879 27212 21888
rect 27160 21845 27169 21879
rect 27169 21845 27203 21879
rect 27203 21845 27212 21879
rect 27160 21836 27212 21845
rect 27252 21836 27304 21888
rect 29184 21904 29236 21956
rect 29736 21904 29788 21956
rect 30472 22040 30524 22092
rect 30104 22015 30156 22024
rect 30104 21981 30113 22015
rect 30113 21981 30147 22015
rect 30147 21981 30156 22015
rect 30104 21972 30156 21981
rect 28540 21879 28592 21888
rect 28540 21845 28549 21879
rect 28549 21845 28583 21879
rect 28583 21845 28592 21879
rect 28540 21836 28592 21845
rect 29460 21836 29512 21888
rect 30104 21836 30156 21888
rect 32128 22040 32180 22092
rect 33048 22040 33100 22092
rect 34704 22083 34756 22092
rect 34704 22049 34713 22083
rect 34713 22049 34747 22083
rect 34747 22049 34756 22083
rect 34704 22040 34756 22049
rect 35348 22040 35400 22092
rect 35440 22040 35492 22092
rect 42708 22083 42760 22092
rect 42708 22049 42717 22083
rect 42717 22049 42751 22083
rect 42751 22049 42760 22083
rect 42708 22040 42760 22049
rect 46664 22083 46716 22092
rect 46664 22049 46673 22083
rect 46673 22049 46707 22083
rect 46707 22049 46716 22083
rect 46664 22040 46716 22049
rect 33968 21972 34020 22024
rect 35624 21904 35676 21956
rect 41604 21972 41656 22024
rect 42616 21972 42668 22024
rect 45468 22015 45520 22024
rect 45468 21981 45477 22015
rect 45477 21981 45511 22015
rect 45511 21981 45520 22015
rect 45468 21972 45520 21981
rect 42800 21904 42852 21956
rect 45652 21947 45704 21956
rect 45652 21913 45661 21947
rect 45661 21913 45695 21947
rect 45695 21913 45704 21947
rect 45652 21904 45704 21913
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 38936 21879 38988 21888
rect 38936 21845 38945 21879
rect 38945 21845 38979 21879
rect 38979 21845 38988 21879
rect 38936 21836 38988 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12624 21675 12676 21684
rect 12624 21641 12633 21675
rect 12633 21641 12667 21675
rect 12667 21641 12676 21675
rect 12624 21632 12676 21641
rect 12900 21632 12952 21684
rect 16856 21632 16908 21684
rect 17040 21632 17092 21684
rect 20720 21632 20772 21684
rect 27160 21632 27212 21684
rect 3516 21564 3568 21616
rect 8760 21496 8812 21548
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 12992 21496 13044 21548
rect 13728 21539 13780 21548
rect 9128 21428 9180 21480
rect 6920 21360 6972 21412
rect 12716 21428 12768 21480
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 18236 21564 18288 21616
rect 18420 21607 18472 21616
rect 18420 21573 18429 21607
rect 18429 21573 18463 21607
rect 18463 21573 18472 21607
rect 18420 21564 18472 21573
rect 18512 21564 18564 21616
rect 22652 21564 22704 21616
rect 29184 21632 29236 21684
rect 28540 21564 28592 21616
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 13084 21360 13136 21412
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 14924 21428 14976 21480
rect 18328 21428 18380 21480
rect 20812 21496 20864 21548
rect 22192 21496 22244 21548
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 21732 21428 21784 21480
rect 23388 21496 23440 21548
rect 26148 21496 26200 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 32128 21632 32180 21684
rect 35624 21675 35676 21684
rect 35624 21641 35633 21675
rect 35633 21641 35667 21675
rect 35667 21641 35676 21675
rect 35624 21632 35676 21641
rect 44088 21632 44140 21684
rect 45652 21675 45704 21684
rect 45652 21641 45661 21675
rect 45661 21641 45695 21675
rect 45695 21641 45704 21675
rect 45652 21632 45704 21641
rect 29736 21564 29788 21616
rect 38936 21607 38988 21616
rect 38936 21573 38945 21607
rect 38945 21573 38979 21607
rect 38979 21573 38988 21607
rect 38936 21564 38988 21573
rect 42708 21564 42760 21616
rect 26424 21496 26476 21505
rect 32772 21496 32824 21548
rect 33508 21496 33560 21548
rect 37280 21496 37332 21548
rect 42616 21539 42668 21548
rect 42616 21505 42625 21539
rect 42625 21505 42659 21539
rect 42659 21505 42668 21539
rect 42616 21496 42668 21505
rect 27252 21428 27304 21480
rect 27528 21471 27580 21480
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 28264 21428 28316 21480
rect 18512 21360 18564 21412
rect 21456 21360 21508 21412
rect 23020 21360 23072 21412
rect 18236 21292 18288 21344
rect 18788 21335 18840 21344
rect 18788 21301 18797 21335
rect 18797 21301 18831 21335
rect 18831 21301 18840 21335
rect 18788 21292 18840 21301
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 23756 21335 23808 21344
rect 23756 21301 23765 21335
rect 23765 21301 23799 21335
rect 23799 21301 23808 21335
rect 23756 21292 23808 21301
rect 25412 21335 25464 21344
rect 25412 21301 25421 21335
rect 25421 21301 25455 21335
rect 25455 21301 25464 21335
rect 25412 21292 25464 21301
rect 26056 21292 26108 21344
rect 39120 21428 39172 21480
rect 42800 21471 42852 21480
rect 42800 21437 42809 21471
rect 42809 21437 42843 21471
rect 42843 21437 42852 21471
rect 42800 21428 42852 21437
rect 45744 21496 45796 21548
rect 46204 21539 46256 21548
rect 46204 21505 46213 21539
rect 46213 21505 46247 21539
rect 46247 21505 46256 21539
rect 46204 21496 46256 21505
rect 46112 21428 46164 21480
rect 43260 21360 43312 21412
rect 28908 21292 28960 21344
rect 30472 21292 30524 21344
rect 47492 21496 47544 21548
rect 46664 21428 46716 21480
rect 46480 21292 46532 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 9128 21131 9180 21140
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 12716 21131 12768 21140
rect 12716 21097 12725 21131
rect 12725 21097 12759 21131
rect 12759 21097 12768 21131
rect 12716 21088 12768 21097
rect 12900 21088 12952 21140
rect 14464 21131 14516 21140
rect 14464 21097 14473 21131
rect 14473 21097 14507 21131
rect 14507 21097 14516 21131
rect 14464 21088 14516 21097
rect 14924 21088 14976 21140
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 22192 21088 22244 21140
rect 23020 21088 23072 21140
rect 28264 21131 28316 21140
rect 21548 21020 21600 21072
rect 28264 21097 28273 21131
rect 28273 21097 28307 21131
rect 28307 21097 28316 21131
rect 28264 21088 28316 21097
rect 28356 21088 28408 21140
rect 45468 21088 45520 21140
rect 15936 20952 15988 21004
rect 8300 20884 8352 20936
rect 9588 20884 9640 20936
rect 10324 20927 10376 20936
rect 10324 20893 10333 20927
rect 10333 20893 10367 20927
rect 10367 20893 10376 20927
rect 10324 20884 10376 20893
rect 15108 20884 15160 20936
rect 17316 20884 17368 20936
rect 18788 20952 18840 21004
rect 20536 20995 20588 21004
rect 20536 20961 20545 20995
rect 20545 20961 20579 20995
rect 20579 20961 20588 20995
rect 20536 20952 20588 20961
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 11244 20859 11296 20868
rect 11244 20825 11253 20859
rect 11253 20825 11287 20859
rect 11287 20825 11296 20859
rect 11244 20816 11296 20825
rect 11704 20816 11756 20868
rect 13728 20816 13780 20868
rect 18512 20884 18564 20936
rect 19340 20884 19392 20936
rect 21732 20952 21784 21004
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 21824 20884 21876 20936
rect 22008 20884 22060 20936
rect 9772 20791 9824 20800
rect 9772 20757 9781 20791
rect 9781 20757 9815 20791
rect 9815 20757 9824 20791
rect 9772 20748 9824 20757
rect 14280 20791 14332 20800
rect 14280 20757 14305 20791
rect 14305 20757 14332 20791
rect 14280 20748 14332 20757
rect 15292 20748 15344 20800
rect 17960 20748 18012 20800
rect 18420 20816 18472 20868
rect 19616 20816 19668 20868
rect 20076 20816 20128 20868
rect 20720 20816 20772 20868
rect 21548 20816 21600 20868
rect 19984 20748 20036 20800
rect 27528 20952 27580 21004
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 27712 20927 27764 20936
rect 27712 20893 27722 20927
rect 27722 20893 27756 20927
rect 27756 20893 27764 20927
rect 27712 20884 27764 20893
rect 27896 20927 27948 20936
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 27896 20884 27948 20893
rect 28080 20927 28132 20936
rect 28080 20893 28094 20927
rect 28094 20893 28128 20927
rect 28128 20893 28132 20927
rect 28080 20884 28132 20893
rect 25136 20859 25188 20868
rect 25136 20825 25145 20859
rect 25145 20825 25179 20859
rect 25179 20825 25188 20859
rect 25136 20816 25188 20825
rect 25412 20816 25464 20868
rect 22468 20748 22520 20800
rect 24492 20748 24544 20800
rect 26608 20791 26660 20800
rect 26608 20757 26617 20791
rect 26617 20757 26651 20791
rect 26651 20757 26660 20791
rect 26608 20748 26660 20757
rect 27804 20816 27856 20868
rect 28908 20816 28960 20868
rect 29184 21020 29236 21072
rect 42432 21020 42484 21072
rect 30380 20995 30432 21004
rect 30380 20961 30389 20995
rect 30389 20961 30423 20995
rect 30423 20961 30432 20995
rect 30380 20952 30432 20961
rect 30472 20927 30524 20936
rect 30472 20893 30481 20927
rect 30481 20893 30515 20927
rect 30515 20893 30524 20927
rect 30472 20884 30524 20893
rect 42524 20952 42576 21004
rect 46480 20995 46532 21004
rect 46480 20961 46489 20995
rect 46489 20961 46523 20995
rect 46523 20961 46532 20995
rect 46480 20952 46532 20961
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 42616 20884 42668 20936
rect 28356 20748 28408 20800
rect 29000 20748 29052 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 8760 20544 8812 20596
rect 9404 20544 9456 20596
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 14740 20544 14792 20596
rect 17592 20544 17644 20596
rect 8300 20408 8352 20460
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 13176 20476 13228 20528
rect 12900 20408 12952 20460
rect 3976 20272 4028 20324
rect 13728 20408 13780 20460
rect 16580 20408 16632 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17776 20476 17828 20528
rect 18420 20476 18472 20528
rect 17960 20408 18012 20460
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 18236 20383 18288 20392
rect 18236 20349 18245 20383
rect 18245 20349 18279 20383
rect 18279 20349 18288 20383
rect 18236 20340 18288 20349
rect 18696 20340 18748 20392
rect 12624 20272 12676 20324
rect 13084 20272 13136 20324
rect 14280 20272 14332 20324
rect 17316 20272 17368 20324
rect 18972 20272 19024 20324
rect 20720 20544 20772 20596
rect 25136 20544 25188 20596
rect 27712 20544 27764 20596
rect 20904 20519 20956 20528
rect 20904 20485 20913 20519
rect 20913 20485 20947 20519
rect 20947 20485 20956 20519
rect 20904 20476 20956 20485
rect 22376 20476 22428 20528
rect 23756 20476 23808 20528
rect 24492 20519 24544 20528
rect 24492 20485 24501 20519
rect 24501 20485 24535 20519
rect 24535 20485 24544 20519
rect 24492 20476 24544 20485
rect 20076 20340 20128 20392
rect 20444 20383 20496 20392
rect 20444 20349 20453 20383
rect 20453 20349 20487 20383
rect 20487 20349 20496 20383
rect 20444 20340 20496 20349
rect 20812 20408 20864 20460
rect 22468 20451 22520 20460
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 26608 20476 26660 20528
rect 27344 20519 27396 20528
rect 27344 20485 27353 20519
rect 27353 20485 27387 20519
rect 27387 20485 27396 20519
rect 27344 20476 27396 20485
rect 29276 20544 29328 20596
rect 29828 20544 29880 20596
rect 45928 20544 45980 20596
rect 42616 20476 42668 20528
rect 43168 20476 43220 20528
rect 25964 20451 26016 20460
rect 21088 20340 21140 20392
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 26056 20451 26108 20460
rect 26056 20417 26065 20451
rect 26065 20417 26099 20451
rect 26099 20417 26108 20451
rect 26056 20408 26108 20417
rect 27988 20408 28040 20460
rect 29000 20408 29052 20460
rect 29184 20451 29236 20460
rect 29184 20417 29193 20451
rect 29193 20417 29227 20451
rect 29227 20417 29236 20451
rect 29184 20408 29236 20417
rect 29276 20451 29328 20460
rect 29276 20417 29285 20451
rect 29285 20417 29319 20451
rect 29319 20417 29328 20451
rect 45468 20451 45520 20460
rect 29276 20408 29328 20417
rect 45468 20417 45477 20451
rect 45477 20417 45511 20451
rect 45511 20417 45520 20451
rect 45468 20408 45520 20417
rect 46020 20451 46072 20460
rect 46020 20417 46029 20451
rect 46029 20417 46063 20451
rect 46063 20417 46072 20451
rect 46020 20408 46072 20417
rect 28080 20340 28132 20392
rect 29460 20340 29512 20392
rect 45744 20340 45796 20392
rect 12072 20204 12124 20256
rect 12348 20204 12400 20256
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 18144 20204 18196 20256
rect 19432 20204 19484 20256
rect 21640 20204 21692 20256
rect 43168 20247 43220 20256
rect 43168 20213 43177 20247
rect 43177 20213 43211 20247
rect 43211 20213 43220 20247
rect 43168 20204 43220 20213
rect 46480 20204 46532 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 11244 20000 11296 20052
rect 19892 20000 19944 20052
rect 20536 20000 20588 20052
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 22008 20043 22060 20052
rect 22008 20009 22017 20043
rect 22017 20009 22051 20043
rect 22051 20009 22060 20043
rect 22008 20000 22060 20009
rect 22560 20000 22612 20052
rect 25228 20000 25280 20052
rect 25964 20000 26016 20052
rect 27620 20000 27672 20052
rect 40684 20000 40736 20052
rect 45560 20000 45612 20052
rect 17960 19932 18012 19984
rect 18696 19932 18748 19984
rect 9220 19864 9272 19916
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 15292 19907 15344 19916
rect 1768 19796 1820 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 18420 19864 18472 19916
rect 19064 19864 19116 19916
rect 12992 19839 13044 19848
rect 12256 19796 12308 19805
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13268 19796 13320 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 11612 19728 11664 19780
rect 12900 19728 12952 19780
rect 14832 19728 14884 19780
rect 17224 19796 17276 19848
rect 18880 19796 18932 19848
rect 21732 19864 21784 19916
rect 16856 19728 16908 19780
rect 17868 19771 17920 19780
rect 17868 19737 17877 19771
rect 17877 19737 17911 19771
rect 17911 19737 17920 19771
rect 17868 19728 17920 19737
rect 18328 19728 18380 19780
rect 19064 19728 19116 19780
rect 19892 19771 19944 19780
rect 19892 19737 19901 19771
rect 19901 19737 19935 19771
rect 19935 19737 19944 19771
rect 19892 19728 19944 19737
rect 20904 19796 20956 19848
rect 24400 19864 24452 19916
rect 29184 19864 29236 19916
rect 24676 19839 24728 19848
rect 12808 19660 12860 19712
rect 18236 19660 18288 19712
rect 18880 19660 18932 19712
rect 20076 19703 20128 19712
rect 20076 19669 20085 19703
rect 20085 19669 20119 19703
rect 20119 19669 20128 19703
rect 20076 19660 20128 19669
rect 20812 19728 20864 19780
rect 20904 19703 20956 19712
rect 20904 19669 20929 19703
rect 20929 19669 20956 19703
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 25136 19728 25188 19780
rect 28448 19796 28500 19848
rect 30012 19839 30064 19848
rect 30012 19805 30021 19839
rect 30021 19805 30055 19839
rect 30055 19805 30064 19839
rect 30012 19796 30064 19805
rect 45468 19932 45520 19984
rect 46112 19932 46164 19984
rect 46480 19907 46532 19916
rect 46480 19873 46489 19907
rect 46489 19873 46523 19907
rect 46523 19873 46532 19907
rect 46480 19864 46532 19873
rect 45560 19796 45612 19848
rect 46204 19796 46256 19848
rect 45928 19728 45980 19780
rect 47308 19728 47360 19780
rect 20904 19660 20956 19669
rect 22468 19660 22520 19712
rect 46112 19660 46164 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 12992 19456 13044 19508
rect 9404 19431 9456 19440
rect 9404 19397 9413 19431
rect 9413 19397 9447 19431
rect 9447 19397 9456 19431
rect 9404 19388 9456 19397
rect 13084 19388 13136 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 9588 19320 9640 19372
rect 12624 19320 12676 19372
rect 14096 19456 14148 19508
rect 16028 19456 16080 19508
rect 14924 19388 14976 19440
rect 17040 19388 17092 19440
rect 17776 19456 17828 19508
rect 18236 19456 18288 19508
rect 18972 19499 19024 19508
rect 18972 19465 18981 19499
rect 18981 19465 19015 19499
rect 19015 19465 19024 19499
rect 18972 19456 19024 19465
rect 45468 19456 45520 19508
rect 45928 19456 45980 19508
rect 14832 19320 14884 19372
rect 15568 19363 15620 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 9220 19252 9272 19304
rect 13452 19295 13504 19304
rect 3884 19184 3936 19236
rect 3424 19116 3476 19168
rect 12992 19116 13044 19168
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 15568 19329 15577 19363
rect 15577 19329 15611 19363
rect 15611 19329 15620 19363
rect 15568 19320 15620 19329
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19340 19320 19392 19372
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 24584 19320 24636 19372
rect 40684 19388 40736 19440
rect 43168 19320 43220 19372
rect 43904 19320 43956 19372
rect 45560 19388 45612 19440
rect 45744 19320 45796 19372
rect 46112 19363 46164 19372
rect 46112 19329 46121 19363
rect 46121 19329 46155 19363
rect 46155 19329 46164 19363
rect 46112 19320 46164 19329
rect 22376 19252 22428 19304
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 46204 19252 46256 19304
rect 17960 19184 18012 19236
rect 17500 19116 17552 19168
rect 18144 19116 18196 19168
rect 23020 19116 23072 19168
rect 24400 19116 24452 19168
rect 27620 19159 27672 19168
rect 27620 19125 27629 19159
rect 27629 19125 27663 19159
rect 27663 19125 27672 19159
rect 27620 19116 27672 19125
rect 41328 19116 41380 19168
rect 41420 19116 41472 19168
rect 47768 19159 47820 19168
rect 47768 19125 47777 19159
rect 47777 19125 47811 19159
rect 47811 19125 47820 19159
rect 47768 19116 47820 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1952 18912 2004 18964
rect 2320 18912 2372 18964
rect 4804 18844 4856 18896
rect 9220 18819 9272 18828
rect 9220 18785 9229 18819
rect 9229 18785 9263 18819
rect 9263 18785 9272 18819
rect 9220 18776 9272 18785
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 13452 18912 13504 18964
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 14924 18955 14976 18964
rect 14924 18921 14933 18955
rect 14933 18921 14967 18955
rect 14967 18921 14976 18955
rect 14924 18912 14976 18921
rect 12992 18844 13044 18896
rect 17960 18912 18012 18964
rect 18328 18955 18380 18964
rect 18328 18921 18337 18955
rect 18337 18921 18371 18955
rect 18371 18921 18380 18955
rect 18328 18912 18380 18921
rect 18512 18955 18564 18964
rect 18512 18921 18521 18955
rect 18521 18921 18555 18955
rect 18555 18921 18564 18955
rect 18512 18912 18564 18921
rect 19984 18955 20036 18964
rect 19984 18921 19993 18955
rect 19993 18921 20027 18955
rect 20027 18921 20036 18955
rect 19984 18912 20036 18921
rect 20260 18912 20312 18964
rect 20904 18955 20956 18964
rect 20904 18921 20913 18955
rect 20913 18921 20947 18955
rect 20947 18921 20956 18955
rect 20904 18912 20956 18921
rect 17500 18887 17552 18896
rect 17500 18853 17509 18887
rect 17509 18853 17543 18887
rect 17543 18853 17552 18887
rect 17500 18844 17552 18853
rect 32496 18912 32548 18964
rect 46020 18912 46072 18964
rect 22376 18844 22428 18896
rect 28172 18844 28224 18896
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 6552 18708 6604 18760
rect 2044 18640 2096 18692
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 12900 18708 12952 18760
rect 14464 18708 14516 18760
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 26516 18776 26568 18828
rect 27528 18819 27580 18828
rect 27528 18785 27537 18819
rect 27537 18785 27571 18819
rect 27571 18785 27580 18819
rect 27528 18776 27580 18785
rect 12808 18640 12860 18692
rect 17224 18683 17276 18692
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 16948 18572 17000 18624
rect 17224 18649 17233 18683
rect 17233 18649 17267 18683
rect 17267 18649 17276 18683
rect 17224 18640 17276 18649
rect 24400 18751 24452 18760
rect 18144 18683 18196 18692
rect 18144 18649 18153 18683
rect 18153 18649 18187 18683
rect 18187 18649 18196 18683
rect 18144 18640 18196 18649
rect 18052 18572 18104 18624
rect 20628 18640 20680 18692
rect 20720 18683 20772 18692
rect 20720 18649 20745 18683
rect 20745 18649 20772 18683
rect 20720 18640 20772 18649
rect 18696 18572 18748 18624
rect 19984 18572 20036 18624
rect 20996 18572 21048 18624
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 41328 18844 41380 18896
rect 41420 18819 41472 18828
rect 41420 18785 41429 18819
rect 41429 18785 41463 18819
rect 41463 18785 41472 18819
rect 41420 18776 41472 18785
rect 45836 18776 45888 18828
rect 46020 18776 46072 18828
rect 47768 18776 47820 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 41236 18751 41288 18760
rect 41236 18717 41245 18751
rect 41245 18717 41279 18751
rect 41279 18717 41288 18751
rect 41236 18708 41288 18717
rect 45560 18751 45612 18760
rect 45560 18717 45569 18751
rect 45569 18717 45603 18751
rect 45603 18717 45612 18751
rect 45560 18708 45612 18717
rect 45928 18708 45980 18760
rect 27712 18640 27764 18692
rect 22744 18572 22796 18624
rect 24492 18615 24544 18624
rect 24492 18581 24501 18615
rect 24501 18581 24535 18615
rect 24535 18581 24544 18615
rect 24492 18572 24544 18581
rect 24768 18572 24820 18624
rect 30656 18683 30708 18692
rect 29092 18572 29144 18624
rect 30656 18649 30665 18683
rect 30665 18649 30699 18683
rect 30699 18649 30708 18683
rect 30656 18640 30708 18649
rect 47676 18640 47728 18692
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2320 18368 2372 18420
rect 4988 18368 5040 18420
rect 25688 18411 25740 18420
rect 25688 18377 25697 18411
rect 25697 18377 25731 18411
rect 25731 18377 25740 18411
rect 25688 18368 25740 18377
rect 11520 18300 11572 18352
rect 14188 18300 14240 18352
rect 16948 18343 17000 18352
rect 16948 18309 16957 18343
rect 16957 18309 16991 18343
rect 16991 18309 17000 18343
rect 16948 18300 17000 18309
rect 17960 18300 18012 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 14464 18232 14516 18284
rect 15568 18232 15620 18284
rect 19340 18275 19392 18284
rect 19340 18241 19349 18275
rect 19349 18241 19383 18275
rect 19383 18241 19392 18275
rect 19340 18232 19392 18241
rect 19432 18232 19484 18284
rect 20536 18300 20588 18352
rect 23020 18343 23072 18352
rect 23020 18309 23029 18343
rect 23029 18309 23063 18343
rect 23063 18309 23072 18343
rect 23020 18300 23072 18309
rect 24492 18300 24544 18352
rect 30656 18368 30708 18420
rect 40224 18368 40276 18420
rect 47676 18411 47728 18420
rect 47676 18377 47685 18411
rect 47685 18377 47719 18411
rect 47719 18377 47728 18411
rect 47676 18368 47728 18377
rect 19984 18232 20036 18284
rect 20996 18275 21048 18284
rect 20996 18241 21005 18275
rect 21005 18241 21039 18275
rect 21039 18241 21048 18275
rect 20996 18232 21048 18241
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 22744 18275 22796 18284
rect 21824 18232 21876 18241
rect 13360 18164 13412 18216
rect 14280 18164 14332 18216
rect 20444 18164 20496 18216
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 25504 18232 25556 18284
rect 27620 18300 27672 18352
rect 46388 18275 46440 18284
rect 46388 18241 46397 18275
rect 46397 18241 46431 18275
rect 46431 18241 46440 18275
rect 46388 18232 46440 18241
rect 47124 18232 47176 18284
rect 47492 18232 47544 18284
rect 24400 18164 24452 18216
rect 18328 18028 18380 18080
rect 18512 18028 18564 18080
rect 19432 18028 19484 18080
rect 20812 18028 20864 18080
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 21916 18071 21968 18080
rect 21916 18037 21925 18071
rect 21925 18037 21959 18071
rect 21959 18037 21968 18071
rect 21916 18028 21968 18037
rect 22468 18028 22520 18080
rect 28080 18164 28132 18216
rect 28172 18207 28224 18216
rect 28172 18173 28181 18207
rect 28181 18173 28215 18207
rect 28215 18173 28224 18207
rect 28172 18164 28224 18173
rect 27160 18028 27212 18080
rect 46848 18028 46900 18080
rect 47032 18071 47084 18080
rect 47032 18037 47041 18071
rect 47041 18037 47075 18071
rect 47075 18037 47084 18071
rect 47032 18028 47084 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 17960 17824 18012 17876
rect 19340 17824 19392 17876
rect 20996 17824 21048 17876
rect 20812 17731 20864 17740
rect 20812 17697 20821 17731
rect 20821 17697 20855 17731
rect 20855 17697 20864 17731
rect 20812 17688 20864 17697
rect 46664 17756 46716 17808
rect 40224 17731 40276 17740
rect 40224 17697 40233 17731
rect 40233 17697 40267 17731
rect 40267 17697 40276 17731
rect 40224 17688 40276 17697
rect 48044 17688 48096 17740
rect 14832 17620 14884 17672
rect 16580 17620 16632 17672
rect 17684 17620 17736 17672
rect 18052 17620 18104 17672
rect 20444 17620 20496 17672
rect 21916 17620 21968 17672
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 25688 17663 25740 17672
rect 25688 17629 25697 17663
rect 25697 17629 25731 17663
rect 25731 17629 25740 17663
rect 25688 17620 25740 17629
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 27068 17663 27120 17672
rect 27068 17629 27077 17663
rect 27077 17629 27111 17663
rect 27111 17629 27120 17663
rect 27068 17620 27120 17629
rect 45468 17620 45520 17672
rect 47860 17620 47912 17672
rect 19340 17552 19392 17604
rect 28080 17552 28132 17604
rect 40408 17552 40460 17604
rect 48044 17552 48096 17604
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 19156 17484 19208 17536
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20260 17484 20312 17536
rect 20720 17484 20772 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 19340 17280 19392 17332
rect 20628 17280 20680 17332
rect 28264 17280 28316 17332
rect 18420 17212 18472 17264
rect 19432 17212 19484 17264
rect 23664 17255 23716 17264
rect 23664 17221 23673 17255
rect 23673 17221 23707 17255
rect 23707 17221 23716 17255
rect 23664 17212 23716 17221
rect 45468 17212 45520 17264
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 2412 17076 2464 17128
rect 3976 17076 4028 17128
rect 6920 17076 6972 17128
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 23664 17076 23716 17128
rect 24768 17144 24820 17196
rect 25228 17144 25280 17196
rect 25688 17187 25740 17196
rect 25688 17153 25697 17187
rect 25697 17153 25731 17187
rect 25731 17153 25740 17187
rect 25688 17144 25740 17153
rect 26424 17144 26476 17196
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 45744 17144 45796 17196
rect 47584 17187 47636 17196
rect 47584 17153 47593 17187
rect 47593 17153 47627 17187
rect 47627 17153 47636 17187
rect 47584 17144 47636 17153
rect 47860 17144 47912 17196
rect 1400 16940 1452 16992
rect 16672 16940 16724 16992
rect 17960 16940 18012 16992
rect 25504 17076 25556 17128
rect 46204 17119 46256 17128
rect 46204 17085 46213 17119
rect 46213 17085 46247 17119
rect 46247 17085 46256 17119
rect 46204 17076 46256 17085
rect 25412 16940 25464 16992
rect 26148 16940 26200 16992
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 19340 16736 19392 16788
rect 19524 16736 19576 16788
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 46572 16736 46624 16788
rect 25964 16668 26016 16720
rect 19156 16532 19208 16584
rect 23388 16575 23440 16584
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 25964 16575 26016 16584
rect 2136 16464 2188 16516
rect 15016 16464 15068 16516
rect 16948 16507 17000 16516
rect 3424 16396 3476 16448
rect 16948 16473 16957 16507
rect 16957 16473 16991 16507
rect 16991 16473 17000 16507
rect 16948 16464 17000 16473
rect 17960 16464 18012 16516
rect 18696 16507 18748 16516
rect 18696 16473 18705 16507
rect 18705 16473 18739 16507
rect 18739 16473 18748 16507
rect 18696 16464 18748 16473
rect 23480 16439 23532 16448
rect 23480 16405 23489 16439
rect 23489 16405 23523 16439
rect 23523 16405 23532 16439
rect 23480 16396 23532 16405
rect 25228 16464 25280 16516
rect 25964 16541 25973 16575
rect 25973 16541 26007 16575
rect 26007 16541 26016 16575
rect 25964 16532 26016 16541
rect 26148 16575 26200 16584
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 27068 16600 27120 16652
rect 47032 16600 47084 16652
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 25412 16396 25464 16448
rect 26332 16439 26384 16448
rect 26332 16405 26341 16439
rect 26341 16405 26375 16439
rect 26375 16405 26384 16439
rect 26332 16396 26384 16405
rect 40040 16464 40092 16516
rect 47676 16464 47728 16516
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 15016 16235 15068 16244
rect 15016 16201 15025 16235
rect 15025 16201 15059 16235
rect 15059 16201 15068 16235
rect 15016 16192 15068 16201
rect 16948 16192 17000 16244
rect 18512 16192 18564 16244
rect 19156 16124 19208 16176
rect 15108 16056 15160 16108
rect 18696 16056 18748 16108
rect 17316 15988 17368 16040
rect 19984 16056 20036 16108
rect 25504 16192 25556 16244
rect 25964 16192 26016 16244
rect 26240 16235 26292 16244
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 26516 16192 26568 16244
rect 23480 16167 23532 16176
rect 23480 16133 23489 16167
rect 23489 16133 23523 16167
rect 23523 16133 23532 16167
rect 23480 16124 23532 16133
rect 26148 16056 26200 16108
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 27804 16099 27856 16108
rect 27804 16065 27813 16099
rect 27813 16065 27847 16099
rect 27847 16065 27856 16099
rect 27804 16056 27856 16065
rect 40040 16099 40092 16108
rect 40040 16065 40049 16099
rect 40049 16065 40083 16099
rect 40083 16065 40092 16099
rect 40040 16056 40092 16065
rect 45468 16124 45520 16176
rect 46388 16167 46440 16176
rect 46388 16133 46397 16167
rect 46397 16133 46431 16167
rect 46431 16133 46440 16167
rect 46388 16124 46440 16133
rect 47124 16056 47176 16108
rect 47676 16056 47728 16108
rect 20444 15988 20496 16040
rect 2872 15852 2924 15904
rect 18604 15852 18656 15904
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 27160 15920 27212 15972
rect 40500 15988 40552 16040
rect 41880 16031 41932 16040
rect 41880 15997 41889 16031
rect 41889 15997 41923 16031
rect 41923 15997 41932 16031
rect 41880 15988 41932 15997
rect 44088 16031 44140 16040
rect 44088 15997 44097 16031
rect 44097 15997 44131 16031
rect 44131 15997 44140 16031
rect 44088 15988 44140 15997
rect 45468 16031 45520 16040
rect 45468 15997 45477 16031
rect 45477 15997 45511 16031
rect 45511 15997 45520 16031
rect 45468 15988 45520 15997
rect 46204 15988 46256 16040
rect 46940 15988 46992 16040
rect 48044 15988 48096 16040
rect 46664 15920 46716 15972
rect 46848 15852 46900 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 20444 15691 20496 15700
rect 1768 15444 1820 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 19156 15512 19208 15564
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 25504 15691 25556 15700
rect 25504 15657 25513 15691
rect 25513 15657 25547 15691
rect 25547 15657 25556 15691
rect 25504 15648 25556 15657
rect 27712 15648 27764 15700
rect 40500 15691 40552 15700
rect 40500 15657 40509 15691
rect 40509 15657 40543 15691
rect 40543 15657 40552 15691
rect 40500 15648 40552 15657
rect 44088 15648 44140 15700
rect 45744 15691 45796 15700
rect 45744 15657 45753 15691
rect 45753 15657 45787 15691
rect 45787 15657 45796 15691
rect 45744 15648 45796 15657
rect 47124 15648 47176 15700
rect 19984 15623 20036 15632
rect 19984 15589 19993 15623
rect 19993 15589 20027 15623
rect 20027 15589 20036 15623
rect 19984 15580 20036 15589
rect 20536 15512 20588 15564
rect 20260 15444 20312 15496
rect 19340 15376 19392 15428
rect 20536 15376 20588 15428
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 16672 15308 16724 15360
rect 17960 15308 18012 15360
rect 20904 15444 20956 15496
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 25228 15376 25280 15428
rect 26332 15444 26384 15496
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 40316 15444 40368 15496
rect 43536 15444 43588 15496
rect 43904 15487 43956 15496
rect 43904 15453 43913 15487
rect 43913 15453 43947 15487
rect 43947 15453 43956 15487
rect 43904 15444 43956 15453
rect 46388 15512 46440 15564
rect 46664 15487 46716 15496
rect 46664 15453 46673 15487
rect 46673 15453 46707 15487
rect 46707 15453 46716 15487
rect 46664 15444 46716 15453
rect 47032 15487 47084 15496
rect 47032 15453 47041 15487
rect 47041 15453 47075 15487
rect 47075 15453 47084 15487
rect 47032 15444 47084 15453
rect 47676 15444 47728 15496
rect 48044 15487 48096 15496
rect 46296 15376 46348 15428
rect 48044 15453 48053 15487
rect 48053 15453 48087 15487
rect 48087 15453 48096 15487
rect 48044 15444 48096 15453
rect 20812 15308 20864 15360
rect 22100 15308 22152 15360
rect 30564 15308 30616 15360
rect 48044 15308 48096 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3240 15104 3292 15156
rect 17960 15036 18012 15088
rect 19432 15036 19484 15088
rect 21732 15036 21784 15088
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 22836 15036 22888 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 20996 14968 21048 15020
rect 26240 15104 26292 15156
rect 27068 15147 27120 15156
rect 27068 15113 27077 15147
rect 27077 15113 27111 15147
rect 27111 15113 27120 15147
rect 27068 15104 27120 15113
rect 47032 15104 47084 15156
rect 2228 14900 2280 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 17592 14900 17644 14952
rect 19248 14943 19300 14952
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 20536 14832 20588 14884
rect 46388 14968 46440 15020
rect 26516 14900 26568 14952
rect 26792 14900 26844 14952
rect 27712 14900 27764 14952
rect 43720 14943 43772 14952
rect 43720 14909 43729 14943
rect 43729 14909 43763 14943
rect 43763 14909 43772 14943
rect 43720 14900 43772 14909
rect 45100 14943 45152 14952
rect 45100 14909 45109 14943
rect 45109 14909 45143 14943
rect 45143 14909 45152 14943
rect 45100 14900 45152 14909
rect 46756 14968 46808 15020
rect 47768 15011 47820 15020
rect 47768 14977 47777 15011
rect 47777 14977 47811 15011
rect 47811 14977 47820 15011
rect 47768 14968 47820 14977
rect 46848 14900 46900 14952
rect 27804 14832 27856 14884
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 20260 14764 20312 14816
rect 23572 14807 23624 14816
rect 23572 14773 23581 14807
rect 23581 14773 23615 14807
rect 23615 14773 23624 14807
rect 23572 14764 23624 14773
rect 46480 14764 46532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 19432 14560 19484 14612
rect 20076 14560 20128 14612
rect 21364 14560 21416 14612
rect 21732 14603 21784 14612
rect 21732 14569 21741 14603
rect 21741 14569 21775 14603
rect 21775 14569 21784 14603
rect 21732 14560 21784 14569
rect 22836 14560 22888 14612
rect 43720 14560 43772 14612
rect 47768 14560 47820 14612
rect 3516 14492 3568 14544
rect 15200 14467 15252 14476
rect 15200 14433 15209 14467
rect 15209 14433 15243 14467
rect 15243 14433 15252 14467
rect 15200 14424 15252 14433
rect 19984 14492 20036 14544
rect 23572 14424 23624 14476
rect 30564 14467 30616 14476
rect 30564 14433 30573 14467
rect 30573 14433 30607 14467
rect 30607 14433 30616 14467
rect 30564 14424 30616 14433
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 17316 14356 17368 14408
rect 18420 14356 18472 14408
rect 21824 14356 21876 14408
rect 43536 14399 43588 14408
rect 43536 14365 43545 14399
rect 43545 14365 43579 14399
rect 43579 14365 43588 14399
rect 43536 14356 43588 14365
rect 46756 14424 46808 14476
rect 46480 14399 46532 14408
rect 46480 14365 46489 14399
rect 46489 14365 46523 14399
rect 46523 14365 46532 14399
rect 46480 14356 46532 14365
rect 46664 14356 46716 14408
rect 46848 14356 46900 14408
rect 20260 14288 20312 14340
rect 20812 14331 20864 14340
rect 20812 14297 20821 14331
rect 20821 14297 20855 14331
rect 20855 14297 20864 14331
rect 20812 14288 20864 14297
rect 32220 14331 32272 14340
rect 32220 14297 32229 14331
rect 32229 14297 32263 14331
rect 32263 14297 32272 14331
rect 32220 14288 32272 14297
rect 46388 14288 46440 14340
rect 46112 14263 46164 14272
rect 46112 14229 46121 14263
rect 46121 14229 46155 14263
rect 46155 14229 46164 14263
rect 46112 14220 46164 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2136 14016 2188 14068
rect 41052 14016 41104 14068
rect 46756 14016 46808 14068
rect 19248 13948 19300 14000
rect 20904 13991 20956 14000
rect 20904 13957 20913 13991
rect 20913 13957 20947 13991
rect 20947 13957 20956 13991
rect 20904 13948 20956 13957
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 20812 13923 20864 13932
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 20260 13812 20312 13864
rect 43536 13812 43588 13864
rect 45744 13880 45796 13932
rect 46020 13923 46072 13932
rect 46020 13889 46029 13923
rect 46029 13889 46063 13923
rect 46063 13889 46072 13923
rect 46020 13880 46072 13889
rect 46112 13923 46164 13932
rect 46112 13889 46121 13923
rect 46121 13889 46155 13923
rect 46155 13889 46164 13923
rect 46112 13880 46164 13889
rect 46388 13880 46440 13932
rect 46756 13923 46808 13932
rect 46756 13889 46765 13923
rect 46765 13889 46799 13923
rect 46799 13889 46808 13923
rect 46756 13880 46808 13889
rect 45836 13855 45845 13864
rect 45845 13855 45879 13864
rect 45879 13855 45888 13864
rect 45836 13812 45888 13855
rect 46480 13812 46532 13864
rect 3976 13676 4028 13728
rect 5448 13676 5500 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 23388 13268 23440 13320
rect 46112 13311 46164 13320
rect 46112 13277 46121 13311
rect 46121 13277 46155 13311
rect 46155 13277 46164 13311
rect 46112 13268 46164 13277
rect 46664 13311 46716 13320
rect 46664 13277 46673 13311
rect 46673 13277 46707 13311
rect 46707 13277 46716 13311
rect 46664 13268 46716 13277
rect 46940 13268 46992 13320
rect 47492 13243 47544 13252
rect 47492 13209 47501 13243
rect 47501 13209 47535 13243
rect 47535 13209 47544 13243
rect 47492 13200 47544 13209
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20904 13175 20956 13184
rect 20904 13141 20913 13175
rect 20913 13141 20947 13175
rect 20947 13141 20956 13175
rect 20904 13132 20956 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 46664 12971 46716 12980
rect 46664 12937 46673 12971
rect 46673 12937 46707 12971
rect 46707 12937 46716 12971
rect 46664 12928 46716 12937
rect 20260 12860 20312 12912
rect 45836 12860 45888 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 20628 12724 20680 12776
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 45836 12724 45888 12776
rect 45744 12656 45796 12708
rect 34796 12588 34848 12640
rect 45560 12588 45612 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 46020 12384 46072 12436
rect 19432 12248 19484 12300
rect 20904 12248 20956 12300
rect 46940 12316 46992 12368
rect 46480 12291 46532 12300
rect 46480 12257 46489 12291
rect 46489 12257 46523 12291
rect 46523 12257 46532 12291
rect 46480 12248 46532 12257
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 45560 12180 45612 12232
rect 14832 12112 14884 12164
rect 45744 12180 45796 12232
rect 46296 12112 46348 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 46112 11815 46164 11824
rect 46112 11781 46121 11815
rect 46121 11781 46155 11815
rect 46155 11781 46164 11815
rect 46112 11772 46164 11781
rect 46020 11679 46072 11688
rect 46020 11645 46029 11679
rect 46029 11645 46063 11679
rect 46063 11645 46072 11679
rect 46020 11636 46072 11645
rect 46296 11679 46348 11688
rect 46296 11645 46305 11679
rect 46305 11645 46339 11679
rect 46339 11645 46348 11679
rect 46296 11636 46348 11645
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 47676 11024 47728 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 47676 10795 47728 10804
rect 47676 10761 47685 10795
rect 47685 10761 47719 10795
rect 47719 10761 47728 10795
rect 47676 10752 47728 10761
rect 41052 10616 41104 10668
rect 2780 10412 2832 10464
rect 4804 10412 4856 10464
rect 46296 10412 46348 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19064 10072 19116 10124
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 19432 9979 19484 9988
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 20996 9936 21048 9988
rect 47676 9936 47728 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 19432 9596 19484 9648
rect 47676 9639 47728 9648
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 18236 9528 18288 9580
rect 42708 9528 42760 9580
rect 46848 9528 46900 9580
rect 45376 9460 45428 9512
rect 47860 9528 47912 9580
rect 46112 9392 46164 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 47308 8959 47360 8968
rect 47308 8925 47317 8959
rect 47317 8925 47351 8959
rect 47351 8925 47360 8959
rect 47308 8916 47360 8925
rect 47400 8916 47452 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 47768 8551 47820 8560
rect 47768 8517 47777 8551
rect 47777 8517 47811 8551
rect 47811 8517 47820 8551
rect 47768 8508 47820 8517
rect 38016 8304 38068 8356
rect 41880 8236 41932 8288
rect 45560 8236 45612 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 46204 7896 46256 7948
rect 47400 7896 47452 7948
rect 47952 7939 48004 7948
rect 47952 7905 47961 7939
rect 47961 7905 47995 7939
rect 47995 7905 48004 7939
rect 47952 7896 48004 7905
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 48136 7395 48188 7404
rect 48136 7361 48145 7395
rect 48145 7361 48179 7395
rect 48179 7361 48188 7395
rect 48136 7352 48188 7361
rect 47124 7148 47176 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 47124 6851 47176 6860
rect 47124 6817 47133 6851
rect 47133 6817 47167 6851
rect 47167 6817 47176 6851
rect 47124 6808 47176 6817
rect 48044 6851 48096 6860
rect 48044 6817 48053 6851
rect 48053 6817 48087 6851
rect 48087 6817 48096 6851
rect 48044 6808 48096 6817
rect 1860 6672 1912 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 46756 6264 46808 6316
rect 48136 6307 48188 6316
rect 48136 6273 48145 6307
rect 48145 6273 48179 6307
rect 48179 6273 48188 6307
rect 48136 6264 48188 6273
rect 46204 6239 46256 6248
rect 46204 6205 46213 6239
rect 46213 6205 46247 6239
rect 46247 6205 46256 6239
rect 46204 6196 46256 6205
rect 47952 6103 48004 6112
rect 47952 6069 47961 6103
rect 47961 6069 47995 6103
rect 47995 6069 48004 6103
rect 47952 6060 48004 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 41236 5720 41288 5772
rect 47860 5763 47912 5772
rect 47860 5729 47869 5763
rect 47869 5729 47903 5763
rect 47903 5729 47912 5763
rect 47860 5720 47912 5729
rect 46204 5584 46256 5636
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 18328 5176 18380 5228
rect 18972 5176 19024 5228
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 21732 5176 21784 5228
rect 21916 5176 21968 5228
rect 23480 5244 23532 5296
rect 45652 5312 45704 5364
rect 46020 5287 46072 5296
rect 46020 5253 46029 5287
rect 46029 5253 46063 5287
rect 46063 5253 46072 5287
rect 46020 5244 46072 5253
rect 47952 5244 48004 5296
rect 23848 5176 23900 5228
rect 43260 5176 43312 5228
rect 47860 5219 47912 5228
rect 47860 5185 47869 5219
rect 47869 5185 47903 5219
rect 47903 5185 47912 5219
rect 47860 5176 47912 5185
rect 48044 5176 48096 5228
rect 4068 5108 4120 5160
rect 30012 5108 30064 5160
rect 17960 5040 18012 5092
rect 28724 5040 28776 5092
rect 18880 4972 18932 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 21824 4972 21876 5024
rect 22376 4972 22428 5024
rect 23112 4972 23164 5024
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 45928 4972 45980 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 18328 4811 18380 4820
rect 18328 4777 18337 4811
rect 18337 4777 18371 4811
rect 18371 4777 18380 4811
rect 18328 4768 18380 4777
rect 20260 4768 20312 4820
rect 21732 4768 21784 4820
rect 20352 4632 20404 4684
rect 47492 4700 47544 4752
rect 19432 4564 19484 4616
rect 19984 4564 20036 4616
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 45928 4675 45980 4684
rect 45928 4641 45937 4675
rect 45937 4641 45971 4675
rect 45971 4641 45980 4675
rect 45928 4632 45980 4641
rect 46940 4675 46992 4684
rect 46940 4641 46949 4675
rect 46949 4641 46983 4675
rect 46983 4641 46992 4675
rect 46940 4632 46992 4641
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 23112 4607 23164 4616
rect 23112 4573 23121 4607
rect 23121 4573 23155 4607
rect 23155 4573 23164 4607
rect 23112 4564 23164 4573
rect 42432 4564 42484 4616
rect 43812 4564 43864 4616
rect 45192 4564 45244 4616
rect 20076 4496 20128 4548
rect 19340 4471 19392 4480
rect 19340 4437 19349 4471
rect 19349 4437 19383 4471
rect 19383 4437 19392 4471
rect 19340 4428 19392 4437
rect 20536 4428 20588 4480
rect 23112 4428 23164 4480
rect 23756 4428 23808 4480
rect 43076 4428 43128 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 19432 4224 19484 4276
rect 19984 4267 20036 4276
rect 19984 4233 19993 4267
rect 19993 4233 20027 4267
rect 20027 4233 20036 4267
rect 19984 4224 20036 4233
rect 20628 4267 20680 4276
rect 20628 4233 20637 4267
rect 20637 4233 20671 4267
rect 20671 4233 20680 4267
rect 20628 4224 20680 4233
rect 21916 4267 21968 4276
rect 21916 4233 21925 4267
rect 21925 4233 21959 4267
rect 21959 4233 21968 4267
rect 21916 4224 21968 4233
rect 22468 4224 22520 4276
rect 18052 4156 18104 4208
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7104 4088 7156 4140
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7380 4088 7432 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 17960 4088 18012 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 21272 4156 21324 4208
rect 18880 4088 18932 4140
rect 19340 4088 19392 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 21180 4088 21232 4140
rect 21824 4131 21876 4140
rect 21824 4097 21833 4131
rect 21833 4097 21867 4131
rect 21867 4097 21876 4131
rect 21824 4088 21876 4097
rect 22376 4088 22428 4140
rect 23112 4131 23164 4140
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23756 4131 23808 4140
rect 6920 3952 6972 4004
rect 10876 3952 10928 4004
rect 1952 3884 2004 3936
rect 2780 3884 2832 3936
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 11244 3884 11296 3936
rect 18972 3952 19024 4004
rect 19064 3952 19116 4004
rect 22284 4020 22336 4072
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 39488 4224 39540 4276
rect 23296 4020 23348 4072
rect 18052 3884 18104 3936
rect 19248 3884 19300 3936
rect 24676 3952 24728 4004
rect 22008 3884 22060 3936
rect 22744 3884 22796 3936
rect 24492 3884 24544 3936
rect 29368 4020 29420 4072
rect 36268 4020 36320 4072
rect 38568 4088 38620 4140
rect 39212 4131 39264 4140
rect 39212 4097 39221 4131
rect 39221 4097 39255 4131
rect 39255 4097 39264 4131
rect 39856 4131 39908 4140
rect 39212 4088 39264 4097
rect 39856 4097 39865 4131
rect 39865 4097 39899 4131
rect 39899 4097 39908 4131
rect 39856 4088 39908 4097
rect 41236 4156 41288 4208
rect 41052 4088 41104 4140
rect 41420 4088 41472 4140
rect 39396 4020 39448 4072
rect 41144 4063 41196 4072
rect 41144 4029 41153 4063
rect 41153 4029 41187 4063
rect 41187 4029 41196 4063
rect 41144 4020 41196 4029
rect 43076 4199 43128 4208
rect 43076 4165 43085 4199
rect 43085 4165 43119 4199
rect 43119 4165 43128 4199
rect 43076 4156 43128 4165
rect 45652 4224 45704 4276
rect 45928 4224 45980 4276
rect 45008 4088 45060 4140
rect 46020 4156 46072 4208
rect 48320 4088 48372 4140
rect 45836 4020 45888 4072
rect 45928 4063 45980 4072
rect 45928 4029 45937 4063
rect 45937 4029 45971 4063
rect 45971 4029 45980 4063
rect 45928 4020 45980 4029
rect 24860 3952 24912 4004
rect 38384 3884 38436 3936
rect 38476 3884 38528 3936
rect 40040 3952 40092 4004
rect 41052 3884 41104 3936
rect 41328 3927 41380 3936
rect 41328 3893 41337 3927
rect 41337 3893 41371 3927
rect 41371 3893 41380 3927
rect 41328 3884 41380 3893
rect 41420 3884 41472 3936
rect 45468 3884 45520 3936
rect 45560 3884 45612 3936
rect 47768 3884 47820 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7104 3680 7156 3732
rect 3424 3612 3476 3664
rect 10876 3612 10928 3664
rect 10968 3612 11020 3664
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11888 3680 11940 3732
rect 13912 3680 13964 3732
rect 18696 3680 18748 3732
rect 18604 3612 18656 3664
rect 1308 3476 1360 3528
rect 1768 3476 1820 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 7104 3408 7156 3460
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 13728 3476 13780 3528
rect 19984 3680 20036 3732
rect 20168 3680 20220 3732
rect 32128 3680 32180 3732
rect 32772 3680 32824 3732
rect 38936 3680 38988 3732
rect 39212 3723 39264 3732
rect 39212 3689 39221 3723
rect 39221 3689 39255 3723
rect 39255 3689 39264 3723
rect 39212 3680 39264 3689
rect 19432 3612 19484 3664
rect 19984 3544 20036 3596
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 18420 3476 18472 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 15200 3408 15252 3460
rect 15568 3408 15620 3460
rect 17500 3408 17552 3460
rect 19064 3408 19116 3460
rect 19340 3408 19392 3460
rect 20352 3476 20404 3528
rect 21824 3476 21876 3528
rect 22744 3519 22796 3528
rect 22744 3485 22753 3519
rect 22753 3485 22787 3519
rect 22787 3485 22796 3519
rect 22744 3476 22796 3485
rect 23480 3519 23532 3528
rect 23480 3485 23489 3519
rect 23489 3485 23523 3519
rect 23523 3485 23532 3519
rect 23480 3476 23532 3485
rect 21916 3408 21968 3460
rect 24584 3544 24636 3596
rect 26332 3612 26384 3664
rect 47032 3680 47084 3732
rect 39396 3612 39448 3664
rect 42524 3612 42576 3664
rect 45652 3612 45704 3664
rect 47584 3612 47636 3664
rect 26792 3587 26844 3596
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 26332 3476 26384 3528
rect 26424 3476 26476 3528
rect 26792 3553 26801 3587
rect 26801 3553 26835 3587
rect 26835 3553 26844 3587
rect 26792 3544 26844 3553
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 33048 3476 33100 3485
rect 33232 3476 33284 3528
rect 38016 3544 38068 3596
rect 38476 3519 38528 3528
rect 32772 3408 32824 3460
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 11612 3340 11664 3392
rect 13820 3340 13872 3392
rect 13912 3340 13964 3392
rect 18512 3340 18564 3392
rect 19432 3340 19484 3392
rect 22008 3340 22060 3392
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 24860 3340 24912 3392
rect 27528 3340 27580 3392
rect 30932 3340 30984 3392
rect 32220 3340 32272 3392
rect 32680 3340 32732 3392
rect 36176 3408 36228 3460
rect 36268 3408 36320 3460
rect 37832 3408 37884 3460
rect 38476 3485 38485 3519
rect 38485 3485 38519 3519
rect 38519 3485 38528 3519
rect 38476 3476 38528 3485
rect 39488 3476 39540 3528
rect 39764 3544 39816 3596
rect 41328 3587 41380 3596
rect 41328 3553 41337 3587
rect 41337 3553 41371 3587
rect 41371 3553 41380 3587
rect 41328 3544 41380 3553
rect 45468 3544 45520 3596
rect 39948 3476 40000 3528
rect 40316 3519 40368 3528
rect 40316 3485 40325 3519
rect 40325 3485 40359 3519
rect 40359 3485 40368 3519
rect 40316 3476 40368 3485
rect 38476 3340 38528 3392
rect 39488 3340 39540 3392
rect 41144 3408 41196 3460
rect 41328 3408 41380 3460
rect 45376 3476 45428 3528
rect 45652 3521 45704 3528
rect 45652 3487 45661 3521
rect 45661 3487 45695 3521
rect 45695 3487 45704 3521
rect 46296 3519 46348 3528
rect 45652 3476 45704 3487
rect 46296 3485 46305 3519
rect 46305 3485 46339 3519
rect 46339 3485 46348 3519
rect 46296 3476 46348 3485
rect 42984 3408 43036 3460
rect 45560 3408 45612 3460
rect 48964 3408 49016 3460
rect 42340 3340 42392 3392
rect 42616 3340 42668 3392
rect 45376 3340 45428 3392
rect 45468 3340 45520 3392
rect 46296 3340 46348 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 7288 3111 7340 3120
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 17224 3136 17276 3188
rect 17316 3136 17368 3188
rect 18236 3136 18288 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 18604 3136 18656 3188
rect 13912 3111 13964 3120
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 15200 3068 15252 3120
rect 24768 3111 24820 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 6460 3000 6512 3052
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 8484 3000 8536 3052
rect 11060 3000 11112 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 664 2932 716 2984
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 15200 2932 15252 2984
rect 7012 2864 7064 2916
rect 15292 2864 15344 2916
rect 7380 2796 7432 2848
rect 17316 2864 17368 2916
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 32772 3136 32824 3188
rect 36176 3179 36228 3188
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 25136 2975 25188 2984
rect 24860 2864 24912 2916
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 25228 2864 25280 2916
rect 33048 3111 33100 3120
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 27528 2932 27580 2984
rect 33048 3077 33057 3111
rect 33057 3077 33091 3111
rect 33091 3077 33100 3111
rect 33048 3068 33100 3077
rect 36176 3145 36185 3179
rect 36185 3145 36219 3179
rect 36219 3145 36228 3179
rect 36176 3136 36228 3145
rect 39856 3136 39908 3188
rect 39948 3136 40000 3188
rect 46388 3136 46440 3188
rect 36084 3000 36136 3052
rect 38476 3043 38528 3052
rect 38476 3009 38485 3043
rect 38485 3009 38519 3043
rect 38519 3009 38528 3043
rect 38476 3000 38528 3009
rect 33232 2932 33284 2984
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 40316 3068 40368 3120
rect 42616 3111 42668 3120
rect 42616 3077 42625 3111
rect 42625 3077 42659 3111
rect 42659 3077 42668 3111
rect 42616 3068 42668 3077
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 47768 3111 47820 3120
rect 47768 3077 47777 3111
rect 47777 3077 47811 3111
rect 47811 3077 47820 3111
rect 47768 3068 47820 3077
rect 39488 3000 39540 3052
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 42984 2932 43036 2984
rect 43168 2975 43220 2984
rect 43168 2941 43177 2975
rect 43177 2941 43211 2975
rect 43211 2941 43220 2975
rect 43168 2932 43220 2941
rect 47676 2932 47728 2984
rect 43260 2864 43312 2916
rect 17224 2796 17276 2848
rect 23756 2796 23808 2848
rect 23848 2796 23900 2848
rect 32680 2796 32732 2848
rect 32772 2796 32824 2848
rect 40040 2796 40092 2848
rect 40132 2796 40184 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3240 2592 3292 2644
rect 2964 2524 3016 2576
rect 2872 2499 2924 2508
rect 2872 2465 2881 2499
rect 2881 2465 2915 2499
rect 2915 2465 2924 2499
rect 2872 2456 2924 2465
rect 6000 2456 6052 2508
rect 6920 2456 6972 2508
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 5172 2388 5224 2440
rect 2780 2320 2832 2372
rect 2596 2252 2648 2304
rect 6460 2320 6512 2372
rect 7012 2320 7064 2372
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 9036 2524 9088 2576
rect 9496 2456 9548 2508
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 15476 2388 15528 2440
rect 10048 2320 10100 2372
rect 16120 2320 16172 2372
rect 18144 2592 18196 2644
rect 20076 2592 20128 2644
rect 23848 2592 23900 2644
rect 23940 2592 23992 2644
rect 26884 2592 26936 2644
rect 25228 2524 25280 2576
rect 25320 2524 25372 2576
rect 40500 2567 40552 2576
rect 40500 2533 40509 2567
rect 40509 2533 40543 2567
rect 40543 2533 40552 2567
rect 40500 2524 40552 2533
rect 45744 2524 45796 2576
rect 24308 2456 24360 2508
rect 24492 2499 24544 2508
rect 24492 2465 24501 2499
rect 24501 2465 24535 2499
rect 24535 2465 24544 2499
rect 24492 2456 24544 2465
rect 25504 2499 25556 2508
rect 25504 2465 25513 2499
rect 25513 2465 25547 2499
rect 25547 2465 25556 2499
rect 25504 2456 25556 2465
rect 28448 2499 28500 2508
rect 28448 2465 28457 2499
rect 28457 2465 28491 2499
rect 28491 2465 28500 2499
rect 28448 2456 28500 2465
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 32036 2456 32088 2508
rect 41328 2499 41380 2508
rect 41328 2465 41337 2499
rect 41337 2465 41371 2499
rect 41371 2465 41380 2499
rect 41328 2456 41380 2465
rect 46020 2456 46072 2508
rect 47032 2456 47084 2508
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 20628 2388 20680 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 23204 2388 23256 2440
rect 20996 2320 21048 2372
rect 26884 2388 26936 2440
rect 28356 2388 28408 2440
rect 29644 2388 29696 2440
rect 35440 2388 35492 2440
rect 41236 2388 41288 2440
rect 45468 2431 45520 2440
rect 15200 2252 15252 2304
rect 24492 2252 24544 2304
rect 27068 2320 27120 2372
rect 38016 2320 38068 2372
rect 39304 2320 39356 2372
rect 40592 2320 40644 2372
rect 45468 2397 45477 2431
rect 45477 2397 45511 2431
rect 45511 2397 45520 2431
rect 45468 2388 45520 2397
rect 45836 2388 45888 2440
rect 46204 2320 46256 2372
rect 46388 2320 46440 2372
rect 36360 2252 36412 2304
rect 39028 2252 39080 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 25228 2048 25280 2100
rect 29276 2048 29328 2100
rect 4436 1980 4488 2032
rect 29552 1980 29604 2032
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49200 2034 50000
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 4498 49314 4610 50000
rect 4498 49286 4752 49314
rect 4498 49200 4610 49286
rect 32 23050 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 46578 1440 47631
rect 1964 47054 1992 49200
rect 2608 47054 2636 49200
rect 3252 47054 3280 49200
rect 1952 47048 2004 47054
rect 1952 46990 2004 46996
rect 2596 47048 2648 47054
rect 2596 46990 2648 46996
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3698 47016 3754 47025
rect 3698 46951 3754 46960
rect 2136 46912 2188 46918
rect 2136 46854 2188 46860
rect 2872 46912 2924 46918
rect 2872 46854 2924 46860
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1492 35488 1544 35494
rect 1596 35465 1624 35634
rect 1492 35430 1544 35436
rect 1582 35456 1638 35465
rect 1308 33992 1360 33998
rect 1308 33934 1360 33940
rect 1320 32745 1348 33934
rect 1400 33448 1452 33454
rect 1398 33416 1400 33425
rect 1452 33416 1454 33425
rect 1398 33351 1454 33360
rect 1504 33046 1532 35430
rect 1582 35391 1638 35400
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1596 32978 1624 33798
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1306 32736 1362 32745
rect 1306 32671 1362 32680
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1400 25288 1452 25294
rect 1398 25256 1400 25265
rect 1452 25256 1454 25265
rect 1398 25191 1454 25200
rect 1688 24342 1716 46310
rect 1768 45960 1820 45966
rect 1768 45902 1820 45908
rect 1780 45490 1808 45902
rect 1768 45484 1820 45490
rect 1768 45426 1820 45432
rect 1952 43240 2004 43246
rect 1952 43182 2004 43188
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40384 1912 40390
rect 1860 40326 1912 40332
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 1780 36786 1808 37198
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1872 33046 1900 40326
rect 1964 35894 1992 43182
rect 2148 40458 2176 46854
rect 2884 46646 2912 46854
rect 2872 46640 2924 46646
rect 2872 46582 2924 46588
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2792 45422 2820 46271
rect 2228 45416 2280 45422
rect 2228 45358 2280 45364
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 2240 45082 2268 45358
rect 2228 45076 2280 45082
rect 2228 45018 2280 45024
rect 3422 44976 3478 44985
rect 3422 44911 3478 44920
rect 2412 44872 2464 44878
rect 2412 44814 2464 44820
rect 2136 40452 2188 40458
rect 2136 40394 2188 40400
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 1964 35866 2084 35894
rect 1860 33040 1912 33046
rect 1860 32982 1912 32988
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1768 25220 1820 25226
rect 1768 25162 1820 25168
rect 1676 24336 1728 24342
rect 1676 24278 1728 24284
rect 20 23044 72 23050
rect 20 22986 72 22992
rect 1780 20890 1808 25162
rect 1952 24268 2004 24274
rect 1952 24210 2004 24216
rect 1964 23866 1992 24210
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23225 1900 23666
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1780 20862 1900 20890
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1780 19378 1808 19790
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15026 1808 15438
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1872 6730 1900 20862
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18970 1992 19246
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18698 2084 35866
rect 2148 18766 2176 36110
rect 2424 35894 2452 44814
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 2792 36718 2820 36751
rect 2780 36712 2832 36718
rect 2780 36654 2832 36660
rect 2240 35866 2452 35894
rect 2240 31346 2268 35866
rect 2320 33448 2372 33454
rect 2320 33390 2372 33396
rect 2332 32502 2360 33390
rect 3240 32836 3292 32842
rect 3240 32778 3292 32784
rect 2320 32496 2372 32502
rect 2320 32438 2372 32444
rect 3252 32366 3280 32778
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 19145 2268 19246
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2044 18692 2096 18698
rect 2044 18634 2096 18640
rect 2332 18426 2360 18906
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2424 17134 2452 32302
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 16425 1992 16594
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1950 16416 2006 16425
rect 1950 16351 2006 16360
rect 2148 16250 2176 16458
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 14074 2176 14350
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 2148 4146 2176 14010
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10305 2820 10406
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2884 6914 2912 15846
rect 3252 15162 3280 32302
rect 3436 19174 3464 44911
rect 3514 43616 3570 43625
rect 3514 43551 3570 43560
rect 3528 21622 3556 43551
rect 3712 30122 3740 46951
rect 3896 46442 3924 49200
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4724 47054 4752 49286
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49314 13626 50000
rect 13514 49286 13768 49314
rect 13514 49200 13626 49286
rect 5828 47054 5856 49200
rect 7116 47054 7144 49200
rect 4712 47048 4764 47054
rect 4712 46990 4764 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 4068 46980 4120 46986
rect 4068 46922 4120 46928
rect 4988 46980 5040 46986
rect 4988 46922 5040 46928
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 3976 46504 4028 46510
rect 3976 46446 4028 46452
rect 3884 46436 3936 46442
rect 3884 46378 3936 46384
rect 3988 46170 4016 46446
rect 3976 46164 4028 46170
rect 3976 46106 4028 46112
rect 3790 39536 3846 39545
rect 3790 39471 3846 39480
rect 3700 30116 3752 30122
rect 3700 30058 3752 30064
rect 3804 22506 3832 39471
rect 3976 31680 4028 31686
rect 3976 31622 4028 31628
rect 3988 31385 4016 31622
rect 3974 31376 4030 31385
rect 3974 31311 4030 31320
rect 3974 28656 4030 28665
rect 3974 28591 4030 28600
rect 3988 27946 4016 28591
rect 3976 27940 4028 27946
rect 3976 27882 4028 27888
rect 3792 22500 3844 22506
rect 3792 22442 3844 22448
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3988 19825 4016 20266
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3896 18465 3924 19178
rect 3882 18456 3938 18465
rect 3882 18391 3938 18400
rect 3976 17128 4028 17134
rect 3974 17096 3976 17105
rect 4028 17096 4030 17105
rect 3974 17031 4030 17040
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 2792 6886 2912 6914
rect 3436 6905 3464 16390
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 7585 3556 14486
rect 3976 13728 4028 13734
rect 3974 13696 3976 13705
rect 4028 13696 4030 13705
rect 3974 13631 4030 13640
rect 3514 7576 3570 7585
rect 3514 7511 3570 7520
rect 3422 6896 3478 6905
rect 2792 4146 2820 6886
rect 3422 6831 3478 6840
rect 4080 5166 4108 46922
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4816 10470 4844 18838
rect 5000 18426 5028 46922
rect 6920 46912 6972 46918
rect 6920 46854 6972 46860
rect 5080 46504 5132 46510
rect 5080 46446 5132 46452
rect 5092 46170 5120 46446
rect 5080 46164 5132 46170
rect 5080 46106 5132 46112
rect 6932 31754 6960 46854
rect 6932 31726 7052 31754
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5460 13734 5488 21830
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 6564 4146 6592 18702
rect 6932 17134 6960 21354
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 6920 4004 6972 4010
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1320 800 1348 3470
rect 1780 3058 1808 3470
rect 1964 3126 1992 3878
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2792 2378 2820 3878
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 2964 3528 3016 3534
rect 3436 3505 3464 3606
rect 2964 3470 3016 3476
rect 3422 3496 3478 3505
rect 2976 2582 3004 3470
rect 3422 3431 3478 3440
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 2884 785 2912 2450
rect 3252 1465 3280 2586
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 3896 800 3924 3975
rect 6920 3946 6972 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 6656 3602 6684 3878
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 6012 2514 6040 3470
rect 6472 3058 6500 3470
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6932 2514 6960 3946
rect 7024 2922 7052 31726
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7116 25906 7144 29106
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7116 25294 7144 25842
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7208 4146 7236 31282
rect 7852 30938 7880 46922
rect 8404 45554 8432 49200
rect 9048 47054 9076 49200
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9312 46912 9364 46918
rect 9312 46854 9364 46860
rect 8312 45526 8432 45554
rect 7840 30932 7892 30938
rect 7840 30874 7892 30880
rect 8116 28008 8168 28014
rect 8116 27950 8168 27956
rect 8128 27674 8156 27950
rect 8312 27878 8340 45526
rect 9324 31754 9352 46854
rect 10980 46374 11008 49200
rect 11624 47054 11652 49200
rect 12268 47054 12296 49200
rect 12808 47184 12860 47190
rect 12808 47126 12860 47132
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 12256 47048 12308 47054
rect 12256 46990 12308 46996
rect 11704 46980 11756 46986
rect 11704 46922 11756 46928
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 11612 45960 11664 45966
rect 11612 45902 11664 45908
rect 11624 45626 11652 45902
rect 11612 45620 11664 45626
rect 11612 45562 11664 45568
rect 11716 33658 11744 46922
rect 12164 46504 12216 46510
rect 12164 46446 12216 46452
rect 12176 46170 12204 46446
rect 12164 46164 12216 46170
rect 12164 46106 12216 46112
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 11704 32224 11756 32230
rect 11704 32166 11756 32172
rect 11716 31890 11744 32166
rect 11992 31890 12020 32710
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11980 31884 12032 31890
rect 11980 31826 12032 31832
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 10784 31748 10836 31754
rect 10784 31690 10836 31696
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 8392 29640 8444 29646
rect 8392 29582 8444 29588
rect 8404 29306 8432 29582
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8772 29170 8800 31214
rect 9416 30598 9444 31418
rect 10796 31278 10824 31690
rect 12256 31476 12308 31482
rect 12452 31464 12480 31690
rect 12308 31436 12480 31464
rect 12256 31418 12308 31424
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 9496 31136 9548 31142
rect 9496 31078 9548 31084
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 9508 30870 9536 31078
rect 9496 30864 9548 30870
rect 9496 30806 9548 30812
rect 9692 30802 9720 31078
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 10704 30666 10732 31078
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8956 29238 8984 29582
rect 8944 29232 8996 29238
rect 8944 29174 8996 29180
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 9036 29028 9088 29034
rect 9036 28970 9088 28976
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 9048 27606 9076 28970
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 8852 27464 8904 27470
rect 8852 27406 8904 27412
rect 7576 27130 7604 27406
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7392 26382 7420 26726
rect 7380 26376 7432 26382
rect 7380 26318 7432 26324
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7852 25974 7880 26182
rect 7840 25968 7892 25974
rect 7840 25910 7892 25916
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7576 24818 7604 25094
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 8036 22642 8064 27066
rect 8220 26994 8248 27270
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8220 26790 8248 26930
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8312 26246 8340 26794
rect 8576 26784 8628 26790
rect 8576 26726 8628 26732
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8404 26382 8432 26522
rect 8588 26450 8616 26726
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8864 24614 8892 27406
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9036 27056 9088 27062
rect 9036 26998 9088 27004
rect 9048 26518 9076 26998
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9036 26512 9088 26518
rect 9036 26454 9088 26460
rect 8944 26308 8996 26314
rect 9048 26296 9076 26454
rect 9140 26314 9168 26930
rect 9232 26858 9260 27270
rect 9220 26852 9272 26858
rect 9220 26794 9272 26800
rect 8996 26268 9076 26296
rect 9128 26308 9180 26314
rect 8944 26250 8996 26256
rect 9128 26250 9180 26256
rect 9232 26246 9260 26794
rect 9220 26240 9272 26246
rect 9220 26182 9272 26188
rect 9036 25968 9088 25974
rect 9036 25910 9088 25916
rect 9048 25498 9076 25910
rect 9232 25702 9260 26182
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 8944 24812 8996 24818
rect 8944 24754 8996 24760
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 24188 8892 24550
rect 8956 24342 8984 24754
rect 9048 24682 9076 25230
rect 9036 24676 9088 24682
rect 9036 24618 9088 24624
rect 8944 24336 8996 24342
rect 8944 24278 8996 24284
rect 9048 24206 9076 24618
rect 9036 24200 9088 24206
rect 8864 24160 8984 24188
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8772 21554 8800 23666
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8864 22234 8892 22510
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8956 22098 8984 24160
rect 9036 24142 9088 24148
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22098 9168 22374
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9140 21146 9168 21422
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20466 8340 20878
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8772 20466 8800 20538
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 9232 19922 9260 25638
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9324 21894 9352 22034
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9416 20602 9444 30534
rect 11532 30258 11560 31282
rect 12544 31210 12572 32846
rect 12636 32366 12664 32846
rect 12716 32496 12768 32502
rect 12716 32438 12768 32444
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12624 31884 12676 31890
rect 12624 31826 12676 31832
rect 12636 31482 12664 31826
rect 12624 31476 12676 31482
rect 12624 31418 12676 31424
rect 12532 31204 12584 31210
rect 12532 31146 12584 31152
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12452 30734 12480 31078
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12636 30666 12664 31418
rect 12728 30734 12756 32438
rect 12820 31754 12848 47126
rect 12912 47054 12940 49200
rect 13740 47138 13768 49286
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49450 15558 50000
rect 15304 49422 15558 49450
rect 13740 47110 13860 47138
rect 13832 47054 13860 47110
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 13820 47048 13872 47054
rect 13820 46990 13872 46996
rect 13360 46980 13412 46986
rect 13360 46922 13412 46928
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 12820 31726 13032 31754
rect 12808 31680 12860 31686
rect 12808 31622 12860 31628
rect 12900 31680 12952 31686
rect 12900 31622 12952 31628
rect 12820 31482 12848 31622
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 12912 31414 12940 31622
rect 12900 31408 12952 31414
rect 12900 31350 12952 31356
rect 12808 31340 12860 31346
rect 12808 31282 12860 31288
rect 12820 31210 12848 31282
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12912 30938 12940 31214
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12624 30660 12676 30666
rect 12624 30602 12676 30608
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 9968 29578 9996 29990
rect 11532 29714 11560 30194
rect 11520 29708 11572 29714
rect 11520 29650 11572 29656
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10428 28626 10456 28902
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 9508 26790 9536 28562
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9600 27538 9628 28494
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9692 27606 9720 28086
rect 10704 27606 10732 29446
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11164 27878 11192 29038
rect 11440 28490 11468 29446
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 11532 28370 11560 29106
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 12176 28762 12204 29038
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 12636 28558 12664 29582
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 11440 28342 11560 28370
rect 11440 28082 11468 28342
rect 11428 28076 11480 28082
rect 11428 28018 11480 28024
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 10692 27600 10744 27606
rect 10692 27542 10744 27548
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 11164 27470 11192 27814
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 10060 26926 10088 27406
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 10244 26994 10272 27270
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10048 26920 10100 26926
rect 10048 26862 10100 26868
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9508 26382 9536 26522
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 25294 9812 26182
rect 11256 25838 11284 27270
rect 11440 26874 11468 28018
rect 12636 27470 12664 28494
rect 12912 28150 12940 29582
rect 12900 28144 12952 28150
rect 12820 28104 12900 28132
rect 12716 28008 12768 28014
rect 12716 27950 12768 27956
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11532 26994 11560 27270
rect 12728 27130 12756 27950
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11796 26920 11848 26926
rect 11440 26846 11560 26874
rect 11796 26862 11848 26868
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24750 9628 25094
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24206 9996 24550
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9600 23730 9628 24006
rect 10152 23866 10180 24074
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9600 20942 9628 21830
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18834 9260 19246
rect 9416 18834 9444 19382
rect 9600 19378 9628 20878
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 19922 9812 20742
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7116 3738 7144 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 3058 7144 3402
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4448 2038 4476 2246
rect 4436 2032 4488 2038
rect 4436 1974 4488 1980
rect 5184 800 5212 2382
rect 7024 2378 7052 2450
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6472 800 6500 2314
rect 7208 1714 7236 3538
rect 7300 3126 7328 3878
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7392 2854 7420 4082
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 8484 3052 8536 3058
rect 8404 3012 8484 3040
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7116 1686 7236 1714
rect 7116 800 7144 1686
rect 7760 800 7788 2926
rect 8404 800 8432 3012
rect 8484 2994 8536 3000
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 9048 800 9076 2518
rect 9508 2514 9536 3878
rect 9968 3534 9996 22986
rect 10336 22982 10364 24754
rect 11532 23866 11560 26846
rect 11704 26240 11756 26246
rect 11704 26182 11756 26188
rect 11716 25906 11744 26182
rect 11808 26042 11836 26862
rect 12268 26586 12296 26998
rect 12544 26926 12572 27066
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12360 26586 12388 26726
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12728 26450 12756 27066
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12084 25362 12112 25638
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 24138 11652 24550
rect 11808 24342 11836 25230
rect 12452 24954 12480 25842
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12544 24682 12572 26318
rect 12728 25974 12756 26386
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12820 25906 12848 28104
rect 12900 28086 12952 28092
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12912 27674 12940 27950
rect 12900 27668 12952 27674
rect 12900 27610 12952 27616
rect 13004 26874 13032 31726
rect 13188 31414 13216 32166
rect 13372 31754 13400 46922
rect 14200 46594 14228 49200
rect 15304 47462 15332 49422
rect 15446 49200 15558 49422
rect 16090 49200 16202 50000
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49314 27150 50000
rect 26620 49286 27150 49314
rect 15292 47456 15344 47462
rect 15292 47398 15344 47404
rect 14648 46980 14700 46986
rect 14648 46922 14700 46928
rect 14200 46566 14320 46594
rect 14292 46510 14320 46566
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14188 46504 14240 46510
rect 14188 46446 14240 46452
rect 14280 46504 14332 46510
rect 14280 46446 14332 46452
rect 13556 46170 13584 46446
rect 14200 46170 14228 46446
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14188 46164 14240 46170
rect 14188 46106 14240 46112
rect 14096 45960 14148 45966
rect 14096 45902 14148 45908
rect 14108 41138 14136 45902
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 14660 33590 14688 46922
rect 16132 46918 16160 49200
rect 16488 47456 16540 47462
rect 16488 47398 16540 47404
rect 16120 46912 16172 46918
rect 16120 46854 16172 46860
rect 14648 33584 14700 33590
rect 14648 33526 14700 33532
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14188 32292 14240 32298
rect 14188 32234 14240 32240
rect 14200 31822 14228 32234
rect 14476 32026 14504 32302
rect 14568 32026 14596 32370
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15476 32224 15528 32230
rect 15476 32166 15528 32172
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 14372 31884 14424 31890
rect 14372 31826 14424 31832
rect 14188 31816 14240 31822
rect 14188 31758 14240 31764
rect 14384 31754 14412 31826
rect 13372 31726 13492 31754
rect 14384 31726 14504 31754
rect 13176 31408 13228 31414
rect 13176 31350 13228 31356
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13188 29850 13216 30126
rect 13280 29850 13308 30670
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13176 29844 13228 29850
rect 13176 29786 13228 29792
rect 13268 29844 13320 29850
rect 13268 29786 13320 29792
rect 13372 29646 13400 30602
rect 13464 29782 13492 31726
rect 14476 31686 14504 31726
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14568 31482 14596 31962
rect 15212 31890 15240 32166
rect 15488 31890 15516 32166
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 14648 31748 14700 31754
rect 14648 31690 14700 31696
rect 14556 31476 14608 31482
rect 14556 31418 14608 31424
rect 14188 31408 14240 31414
rect 14188 31350 14240 31356
rect 14200 30938 14228 31350
rect 14660 31278 14688 31690
rect 15672 31482 15700 32370
rect 16408 31754 16436 32370
rect 16316 31726 16436 31754
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 16212 31272 16264 31278
rect 16212 31214 16264 31220
rect 14188 30932 14240 30938
rect 14188 30874 14240 30880
rect 14660 30734 14688 31214
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 16224 30598 16252 31214
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13372 29306 13400 29582
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 13188 28762 13216 29038
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 13464 28558 13492 29718
rect 14556 29572 14608 29578
rect 14556 29514 14608 29520
rect 14568 28626 14596 29514
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 15304 28626 15332 28902
rect 15488 28762 15516 29106
rect 15476 28756 15528 28762
rect 15476 28698 15528 28704
rect 14556 28620 14608 28626
rect 14556 28562 14608 28568
rect 15292 28620 15344 28626
rect 15292 28562 15344 28568
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 15948 28490 15976 29446
rect 16224 29102 16252 30534
rect 16316 29646 16344 31726
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16212 29096 16264 29102
rect 16212 29038 16264 29044
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13464 28150 13492 28358
rect 16316 28218 16344 29582
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13096 27062 13124 27406
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 13004 26846 13124 26874
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12912 26042 12940 26318
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12900 26036 12952 26042
rect 12900 25978 12952 25984
rect 13004 25906 13032 26250
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12532 24676 12584 24682
rect 12532 24618 12584 24624
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 12544 24206 12572 24618
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11532 23730 11560 23802
rect 12268 23730 12296 24142
rect 12728 23798 12756 24686
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 10980 22982 11008 23462
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10336 20942 10364 22918
rect 11348 22030 11376 23054
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11716 22710 11744 22918
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11808 21690 11836 22510
rect 12360 22030 12388 23462
rect 12820 23118 12848 25842
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12912 24410 12940 24550
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 13004 24070 13032 25842
rect 13096 25809 13124 26846
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 15028 26450 15056 26726
rect 15844 26512 15896 26518
rect 15844 26454 15896 26460
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 13280 26042 13308 26182
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13082 25800 13138 25809
rect 13082 25735 13138 25744
rect 13280 25498 13308 25978
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13924 25362 13952 26318
rect 14476 25906 14504 26318
rect 15752 26308 15804 26314
rect 15752 26250 15804 26256
rect 15764 26042 15792 26250
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15856 25922 15884 26454
rect 16500 26450 16528 47398
rect 17420 45554 17448 49200
rect 18708 47054 18736 49200
rect 19432 47184 19484 47190
rect 19432 47126 19484 47132
rect 18696 47048 18748 47054
rect 19444 47025 19472 47126
rect 19996 47122 20024 49200
rect 19984 47116 20036 47122
rect 19984 47058 20036 47064
rect 18696 46990 18748 46996
rect 19430 47016 19486 47025
rect 17592 46980 17644 46986
rect 19430 46951 19486 46960
rect 17592 46922 17644 46928
rect 17420 45526 17540 45554
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16672 31884 16724 31890
rect 16672 31826 16724 31832
rect 16684 31414 16712 31826
rect 16776 31822 16804 32166
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16672 31408 16724 31414
rect 16672 31350 16724 31356
rect 16868 31346 16896 31962
rect 17316 31884 17368 31890
rect 17316 31826 17368 31832
rect 17040 31748 17092 31754
rect 17040 31690 17092 31696
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16776 30954 16804 31282
rect 16960 30954 16988 31622
rect 17052 31346 17080 31690
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 16776 30926 16988 30954
rect 17052 30734 17080 31078
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 16856 30660 16908 30666
rect 16856 30602 16908 30608
rect 16868 30190 16896 30602
rect 17052 30326 17080 30670
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 16868 29102 16896 30126
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16868 28218 16896 29038
rect 16960 28490 16988 30194
rect 17052 29170 17080 30262
rect 17328 30258 17356 31826
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17316 30116 17368 30122
rect 17316 30058 17368 30064
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 16948 28484 17000 28490
rect 16948 28426 17000 28432
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16868 25974 16896 28154
rect 16960 28150 16988 28426
rect 16948 28144 17000 28150
rect 16948 28086 17000 28092
rect 17052 27878 17080 29106
rect 17236 28626 17264 29650
rect 17328 29646 17356 30058
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17328 29306 17356 29582
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17328 28762 17356 29038
rect 17408 28960 17460 28966
rect 17408 28902 17460 28908
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17328 28626 17356 28698
rect 17420 28694 17448 28902
rect 17408 28688 17460 28694
rect 17408 28630 17460 28636
rect 17224 28620 17276 28626
rect 17224 28562 17276 28568
rect 17316 28620 17368 28626
rect 17316 28562 17368 28568
rect 17236 28506 17264 28562
rect 17236 28478 17356 28506
rect 17328 28218 17356 28478
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17040 27872 17092 27878
rect 17040 27814 17092 27820
rect 17420 27470 17448 28358
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 15764 25906 15884 25922
rect 16856 25968 16908 25974
rect 16856 25910 16908 25916
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15752 25900 15884 25906
rect 15804 25894 15884 25900
rect 15752 25842 15804 25848
rect 13912 25356 13964 25362
rect 13912 25298 13964 25304
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13096 24410 13124 25162
rect 13832 24818 13860 25230
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13648 24698 13676 24754
rect 13924 24698 13952 25298
rect 14476 25158 14504 25842
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14844 25362 14872 25638
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14108 24750 14136 25094
rect 14476 24886 14504 25094
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 13648 24670 13952 24698
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 13832 24614 13860 24670
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13832 23526 13860 24550
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22710 12480 22918
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11992 21554 12020 21830
rect 12636 21690 12664 22102
rect 13096 22094 13124 22714
rect 13372 22710 13400 23054
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 14200 22642 14228 22918
rect 14292 22778 14320 23734
rect 15028 23730 15056 25842
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15120 24834 15148 25094
rect 15120 24806 15240 24834
rect 15764 24818 15792 25842
rect 17052 25702 17080 26862
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14384 23186 14412 23462
rect 14476 23322 14504 23598
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 13004 22066 13124 22094
rect 13004 21962 13032 22066
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12992 21956 13044 21962
rect 12992 21898 13044 21904
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 21146 12756 21422
rect 12912 21146 12940 21626
rect 13004 21554 13032 21898
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13280 21486 13308 21966
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11256 20058 11284 20810
rect 11716 20602 11744 20810
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 12912 20466 12940 21082
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 12084 19854 12112 20198
rect 12360 19922 12388 20198
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11532 18358 11560 18566
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10888 3670 10916 3946
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 10060 2378 10088 3334
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 10980 800 11008 3606
rect 11256 3602 11284 3878
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11072 3058 11100 3470
rect 11624 3398 11652 19722
rect 12268 18834 12296 19790
rect 12636 19378 12664 20266
rect 12912 19786 12940 20402
rect 13096 20330 13124 21354
rect 13176 20528 13228 20534
rect 13280 20482 13308 21422
rect 13740 20874 13768 21490
rect 14476 21146 14504 21830
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13228 20476 13308 20482
rect 13176 20470 13308 20476
rect 13188 20454 13308 20470
rect 13740 20466 13768 20810
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 13280 19854 13308 20454
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 14292 20330 14320 20742
rect 14752 20602 14780 22578
rect 15028 22094 15056 23666
rect 15120 23118 15148 23802
rect 15212 23526 15240 24806
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23186 15240 23462
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15028 22066 15148 22094
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14936 21146 14964 21422
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 15120 20942 15148 22066
rect 15304 22030 15332 22918
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14292 19854 14320 20266
rect 12992 19848 13044 19854
rect 13268 19848 13320 19854
rect 12992 19790 13044 19796
rect 13096 19808 13268 19836
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12820 18698 12848 19654
rect 12912 18766 12940 19722
rect 13004 19514 13032 19790
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 13096 19446 13124 19808
rect 13268 19790 13320 19796
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18902 13032 19110
rect 13464 18970 13492 19246
rect 14108 18970 14136 19450
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18222 13400 18566
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 14200 17882 14228 18294
rect 14292 18222 14320 19790
rect 14752 19258 14780 20538
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19378 14872 19722
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14752 19230 14872 19258
rect 14844 18766 14872 19230
rect 14936 18970 14964 19382
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14476 18290 14504 18702
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14844 17678 14872 18702
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 16250 15056 16458
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15120 16114 15148 20878
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15304 19922 15332 20742
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15580 19378 15608 21966
rect 15764 21894 15792 24754
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24070 16896 24550
rect 17052 24138 17080 25638
rect 17144 25294 17172 25774
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 17144 24818 17172 25230
rect 17420 24954 17448 26318
rect 17512 25362 17540 45526
rect 17604 41414 17632 46922
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 20640 46510 20668 49200
rect 19248 46504 19300 46510
rect 19248 46446 19300 46452
rect 20628 46504 20680 46510
rect 20628 46446 20680 46452
rect 18604 46436 18656 46442
rect 18604 46378 18656 46384
rect 18616 46170 18644 46378
rect 19260 46170 19288 46446
rect 20720 46368 20772 46374
rect 20720 46310 20772 46316
rect 18604 46164 18656 46170
rect 18604 46106 18656 46112
rect 19248 46164 19300 46170
rect 19248 46106 19300 46112
rect 20732 46034 20760 46310
rect 21284 46034 21312 49200
rect 22744 47048 22796 47054
rect 22744 46990 22796 46996
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 18512 45960 18564 45966
rect 18512 45902 18564 45908
rect 17604 41386 17908 41414
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17604 31822 17632 32302
rect 17788 32298 17816 32710
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17684 32020 17736 32026
rect 17684 31962 17736 31968
rect 17696 31822 17724 31962
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17604 30394 17632 30738
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17696 26994 17724 31758
rect 17788 31686 17816 32234
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17788 31482 17816 31622
rect 17776 31476 17828 31482
rect 17776 31418 17828 31424
rect 17880 31362 17908 41386
rect 18524 31754 18552 45902
rect 20720 45892 20772 45898
rect 20720 45834 20772 45840
rect 20904 45892 20956 45898
rect 20904 45834 20956 45840
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 20732 45490 20760 45834
rect 20916 45626 20944 45834
rect 20904 45620 20956 45626
rect 20904 45562 20956 45568
rect 20720 45484 20772 45490
rect 20720 45426 20772 45432
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 20732 44198 20760 45426
rect 20720 44192 20772 44198
rect 20720 44134 20772 44140
rect 21364 44192 21416 44198
rect 21364 44134 21416 44140
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 21376 41414 21404 44134
rect 19574 41372 19882 41392
rect 21376 41386 21496 41414
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19168 32842 19196 33050
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 19352 32502 19380 33254
rect 19444 32978 19472 33458
rect 20456 33386 20484 33934
rect 21088 33924 21140 33930
rect 21088 33866 21140 33872
rect 20444 33380 20496 33386
rect 20444 33322 20496 33328
rect 19432 32972 19484 32978
rect 19432 32914 19484 32920
rect 19340 32496 19392 32502
rect 19340 32438 19392 32444
rect 19156 31816 19208 31822
rect 19156 31758 19208 31764
rect 18144 31748 18196 31754
rect 18524 31726 18644 31754
rect 18144 31690 18196 31696
rect 18156 31414 18184 31690
rect 17788 31334 17908 31362
rect 18144 31408 18196 31414
rect 18144 31350 18196 31356
rect 17788 28694 17816 31334
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 17880 30870 17908 31214
rect 18156 30938 18184 31214
rect 18144 30932 18196 30938
rect 18144 30874 18196 30880
rect 17868 30864 17920 30870
rect 17868 30806 17920 30812
rect 18248 30734 18276 31214
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 18144 30660 18196 30666
rect 18144 30602 18196 30608
rect 18156 29646 18184 30602
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17972 29170 18000 29446
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 17776 28688 17828 28694
rect 17776 28630 17828 28636
rect 17972 28558 18000 28970
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17972 28234 18000 28494
rect 17972 28206 18092 28234
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 17972 27674 18000 28086
rect 18064 28014 18092 28206
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 18064 27606 18092 27814
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18052 27464 18104 27470
rect 18156 27418 18184 29582
rect 18248 29238 18276 29650
rect 18236 29232 18288 29238
rect 18236 29174 18288 29180
rect 18104 27412 18184 27418
rect 18052 27406 18184 27412
rect 18064 27390 18184 27406
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17604 26586 17632 26930
rect 17868 26852 17920 26858
rect 17868 26794 17920 26800
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17880 26382 17908 26794
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17880 26042 17908 26318
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16776 23186 16804 23462
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15948 21010 15976 22170
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 16592 20466 16620 22442
rect 16684 22098 16712 22510
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16868 21690 16896 22646
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16960 21554 16988 21830
rect 17052 21690 17080 22102
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17236 21146 17264 21898
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17328 20942 17356 24074
rect 17512 23730 17540 24550
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17604 20942 17632 24006
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17604 20602 17632 20878
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 17788 20534 17816 25774
rect 17880 24818 17908 25978
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17972 24342 18000 25774
rect 17960 24336 18012 24342
rect 17960 24278 18012 24284
rect 18064 23526 18092 27390
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18156 26314 18184 26998
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 18156 25770 18184 26250
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 18156 25226 18184 25706
rect 18144 25220 18196 25226
rect 18144 25162 18196 25168
rect 18156 24274 18184 25162
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19514 16068 20198
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15580 18290 15608 19314
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 16592 17678 16620 20402
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16658 16712 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15502 15148 16050
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 15212 14482 15240 15302
rect 16684 15026 16712 15302
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 3738 11928 4082
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13924 3618 13952 3674
rect 13832 3590 13952 3618
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 13740 3058 13768 3470
rect 13832 3398 13860 3590
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13924 3126 13952 3334
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14200 800 14228 2926
rect 14844 800 14872 12106
rect 16868 3777 16896 19722
rect 17052 19446 17080 20198
rect 17236 19854 17264 20402
rect 17316 20324 17368 20330
rect 17316 20266 17368 20272
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17236 18698 17264 19790
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18358 16988 18566
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16960 16250 16988 16458
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17328 16046 17356 20266
rect 17788 19514 17816 20470
rect 17972 20466 18000 20742
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17972 19802 18000 19926
rect 17880 19786 18000 19802
rect 17868 19780 18000 19786
rect 17920 19774 18000 19780
rect 17868 19722 17920 19728
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18902 17540 19110
rect 17972 18970 18000 19178
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 18064 18630 18092 23462
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18432 22778 18460 22986
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18432 21622 18460 22714
rect 18616 21962 18644 31726
rect 19168 31278 19196 31758
rect 19444 31754 19472 32914
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19432 31748 19484 31754
rect 19432 31690 19484 31696
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 19260 30938 19288 31282
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 19260 29646 19288 30670
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19260 28098 19288 29582
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19352 29170 19380 29446
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19168 28070 19288 28098
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 19168 27470 19196 28070
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19156 27464 19208 27470
rect 19156 27406 19208 27412
rect 19260 26450 19288 27950
rect 19352 27606 19380 28086
rect 19444 28082 19472 31690
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 20456 30802 20484 33322
rect 21100 33318 21128 33866
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 21284 33114 21312 33458
rect 21272 33108 21324 33114
rect 21272 33050 21324 33056
rect 21086 32872 21142 32881
rect 21086 32807 21088 32816
rect 21140 32807 21142 32816
rect 21088 32778 21140 32784
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 21008 30258 21036 31826
rect 21180 30660 21232 30666
rect 21180 30602 21232 30608
rect 21192 30326 21220 30602
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 20548 29170 20576 29718
rect 21008 29306 21036 30194
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 20364 28218 20392 28426
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 26450 19472 26726
rect 19248 26444 19300 26450
rect 19248 26386 19300 26392
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19616 25968 19668 25974
rect 19614 25936 19616 25945
rect 19668 25936 19670 25945
rect 19614 25871 19670 25880
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 19706 25256 19762 25265
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19432 25220 19484 25226
rect 19706 25191 19708 25200
rect 19432 25162 19484 25168
rect 19760 25191 19762 25200
rect 19708 25162 19760 25168
rect 19352 23712 19380 25162
rect 19444 24954 19472 25162
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23798 20024 24006
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19352 23684 19472 23712
rect 19248 23656 19300 23662
rect 19300 23604 19380 23610
rect 19248 23598 19380 23604
rect 19260 23582 19380 23598
rect 19352 23322 19380 23582
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19076 22710 19104 22918
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18420 21616 18472 21622
rect 18420 21558 18472 21564
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18248 21350 18276 21558
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18248 20398 18276 21286
rect 18340 20890 18368 21422
rect 18524 21418 18552 21558
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18524 20942 18552 21354
rect 18512 20936 18564 20942
rect 18340 20874 18460 20890
rect 18512 20878 18564 20884
rect 18340 20868 18472 20874
rect 18340 20862 18420 20868
rect 18340 20466 18368 20862
rect 18420 20810 18472 20816
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 19174 18184 20198
rect 18248 19718 18276 20334
rect 18340 19786 18368 20402
rect 18432 19922 18460 20470
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18236 19712 18288 19718
rect 18432 19666 18460 19858
rect 18236 19654 18288 19660
rect 18340 19638 18460 19666
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18248 18986 18276 19450
rect 18156 18958 18276 18986
rect 18340 18970 18368 19638
rect 18524 18970 18552 20878
rect 18328 18964 18380 18970
rect 18156 18698 18184 18958
rect 18328 18906 18380 18912
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17972 17882 18000 18294
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18064 17678 18092 18566
rect 18340 18086 18368 18906
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17696 17202 17724 17614
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17270 18460 17478
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17328 14414 17356 15982
rect 17696 15502 17724 17138
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17972 16522 18000 16934
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 18524 16250 18552 18022
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18616 15910 18644 21898
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18800 21010 18828 21286
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19352 20942 19380 21898
rect 19444 21536 19472 23684
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19720 22030 19748 22442
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19616 21548 19668 21554
rect 19444 21508 19616 21536
rect 19616 21490 19668 21496
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19990 18736 20334
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18708 18630 18736 19926
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18892 19718 18920 19790
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18892 19378 18920 19654
rect 18984 19514 19012 20266
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19076 19786 19104 19858
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 16522 18736 18566
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16114 18736 16458
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15094 18000 15302
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17604 14618 17632 14894
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 18432 14414 18460 14758
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 19076 10130 19104 19722
rect 19352 19378 19380 20878
rect 19628 20874 19656 21490
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19996 20806 20024 23054
rect 20088 20874 20116 25366
rect 20180 22438 20208 28018
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20076 20868 20128 20874
rect 20076 20810 20128 20816
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19444 18290 19472 20198
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19904 19786 19932 19994
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 18970 20024 20742
rect 20088 20398 20116 20810
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19996 18630 20024 18906
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19352 17882 19380 18226
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19168 16590 19196 17478
rect 19352 17338 19380 17546
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 16794 19380 17274
rect 19444 17270 19472 18022
rect 19996 17542 20024 18226
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19536 16794 19564 17070
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 16182 19196 16526
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19168 15570 19196 16118
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 13938 19196 15506
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19352 14906 19380 15370
rect 19444 15094 19472 15846
rect 19996 15638 20024 16050
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19260 14006 19288 14894
rect 19352 14878 19472 14906
rect 19444 14618 19472 14878
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19444 12306 19472 14554
rect 19996 14550 20024 15574
rect 20088 14618 20116 19654
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19444 9654 19472 9930
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4146 18000 5034
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 18064 3942 18092 4150
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 16854 3768 16910 3777
rect 16854 3703 16910 3712
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15212 3126 15240 3402
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2310 15240 2926
rect 15304 2922 15332 3470
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 15292 2916 15344 2922
rect 15292 2858 15344 2864
rect 15580 2514 15608 3402
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17236 2854 17264 3130
rect 17328 2922 17356 3130
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15488 800 15516 2382
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 800 16160 2314
rect 17512 1986 17540 3402
rect 18156 2650 18184 4082
rect 18248 3194 18276 9522
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18340 4826 18368 5170
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18892 4146 18920 4966
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18984 4010 19012 5170
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 20180 4570 20208 22374
rect 20272 22094 20300 26862
rect 21008 25294 21036 29242
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21100 25906 21128 26862
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21008 24818 21036 25230
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20364 24138 20392 24618
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 21008 24070 21036 24754
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21100 24138 21128 24550
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 22234 20484 22918
rect 20548 22642 20576 23054
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20272 22066 20392 22094
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20272 17542 20300 18906
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 14822 20300 15438
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20272 14346 20300 14758
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20272 13870 20300 14282
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 12918 20300 13126
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20364 12434 20392 22066
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20456 21554 20484 21830
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20548 21010 20576 21830
rect 20732 21690 20760 23054
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20824 22098 20852 22374
rect 20916 22234 20944 22442
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20812 21956 20864 21962
rect 20812 21898 20864 21904
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20824 21554 20852 21898
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20456 18222 20484 20334
rect 20548 20058 20576 20946
rect 20824 20942 20852 21490
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20732 20602 20760 20810
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20732 19802 20760 20538
rect 20824 20466 20852 20878
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20916 19854 20944 20470
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21100 20058 21128 20334
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20904 19848 20956 19854
rect 20732 19786 20852 19802
rect 20904 19790 20956 19796
rect 20732 19780 20864 19786
rect 20732 19774 20812 19780
rect 20732 18698 20760 19774
rect 20812 19722 20864 19728
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 18970 20944 19654
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 17678 20484 18158
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15706 20484 15982
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20548 15570 20576 18294
rect 20640 17338 20668 18634
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 18290 21036 18566
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20824 17746 20852 18022
rect 21008 17882 21036 18022
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 17218 20760 17478
rect 20640 17190 20760 17218
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20548 14890 20576 15370
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20640 12782 20668 17190
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20824 14346 20852 15302
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20824 13938 20852 14282
rect 20916 14006 20944 15438
rect 21008 15026 21036 15846
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20364 12406 20484 12434
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20272 4826 20300 5170
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20364 4690 20392 4966
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4146 19380 4422
rect 19444 4282 19472 4558
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 4282 20024 4558
rect 20076 4548 20128 4554
rect 20180 4542 20392 4570
rect 20076 4490 20128 4496
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18432 3194 18460 3470
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18524 2446 18552 3334
rect 18616 3194 18644 3606
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 17420 1958 17540 1986
rect 17420 800 17448 1958
rect 18708 800 18736 3674
rect 19076 3466 19104 3946
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 19260 2446 19288 3878
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19444 3534 19472 3606
rect 19996 3602 20024 3674
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3058 19380 3402
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3074 19472 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19340 3052 19392 3058
rect 19444 3046 19564 3074
rect 19340 2994 19392 3000
rect 19536 2990 19564 3046
rect 19524 2984 19576 2990
rect 19338 2952 19394 2961
rect 19524 2926 19576 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19338 2887 19394 2896
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19352 800 19380 2887
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2926
rect 20088 2650 20116 4490
rect 20166 3768 20222 3777
rect 20166 3703 20168 3712
rect 20220 3703 20222 3712
rect 20168 3674 20220 3680
rect 20364 3534 20392 4542
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20456 2961 20484 12406
rect 20916 12306 20944 13126
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 20536 4616 20588 4622
rect 20588 4576 20668 4604
rect 20536 4558 20588 4564
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4146 20576 4422
rect 20640 4282 20668 4576
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20442 2952 20498 2961
rect 20442 2887 20498 2896
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20640 800 20668 2382
rect 21008 2378 21036 9930
rect 21192 4146 21220 26250
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21284 25226 21312 25842
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21468 21418 21496 41386
rect 21548 33924 21600 33930
rect 21548 33866 21600 33872
rect 21560 32026 21588 33866
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 32978 22048 33254
rect 22008 32972 22060 32978
rect 22008 32914 22060 32920
rect 22296 32774 22324 33798
rect 22468 33448 22520 33454
rect 22468 33390 22520 33396
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22296 32434 22324 32710
rect 22480 32570 22508 33390
rect 22756 32978 22784 46990
rect 24872 46646 24900 46990
rect 24860 46640 24912 46646
rect 24860 46582 24912 46588
rect 25148 46510 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 25136 46504 25188 46510
rect 25136 46446 25188 46452
rect 24780 46170 24808 46446
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 25516 46034 25544 46990
rect 25792 46034 25820 49200
rect 25504 46028 25556 46034
rect 25504 45970 25556 45976
rect 25780 46028 25832 46034
rect 25780 45970 25832 45976
rect 24584 45960 24636 45966
rect 24584 45902 24636 45908
rect 24596 45626 24624 45902
rect 25412 45892 25464 45898
rect 25412 45834 25464 45840
rect 25424 45626 25452 45834
rect 24584 45620 24636 45626
rect 24584 45562 24636 45568
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 24596 44402 24624 45562
rect 26620 45554 26648 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 30902 49314 31014 50000
rect 30760 49286 31014 49314
rect 28368 47054 28396 49200
rect 29092 47184 29144 47190
rect 29092 47126 29144 47132
rect 28356 47048 28408 47054
rect 28356 46990 28408 46996
rect 28172 46912 28224 46918
rect 28172 46854 28224 46860
rect 28184 46578 28212 46854
rect 28172 46572 28224 46578
rect 28172 46514 28224 46520
rect 26252 45526 26648 45554
rect 25320 45484 25372 45490
rect 25320 45426 25372 45432
rect 24584 44396 24636 44402
rect 24584 44338 24636 44344
rect 25332 37942 25360 45426
rect 26252 41274 26280 45526
rect 27160 41472 27212 41478
rect 27160 41414 27212 41420
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 27172 41206 27200 41414
rect 27160 41200 27212 41206
rect 27160 41142 27212 41148
rect 26056 41064 26108 41070
rect 26056 41006 26108 41012
rect 26068 40594 26096 41006
rect 26056 40588 26108 40594
rect 26056 40530 26108 40536
rect 28080 40452 28132 40458
rect 28080 40394 28132 40400
rect 25320 37936 25372 37942
rect 25320 37878 25372 37884
rect 24676 34060 24728 34066
rect 24676 34002 24728 34008
rect 24492 33924 24544 33930
rect 24492 33866 24544 33872
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23492 33522 23520 33798
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23572 33448 23624 33454
rect 23572 33390 23624 33396
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 22744 32972 22796 32978
rect 22744 32914 22796 32920
rect 23584 32910 23612 33390
rect 23388 32904 23440 32910
rect 23572 32904 23624 32910
rect 23440 32864 23520 32892
rect 23388 32846 23440 32852
rect 22744 32768 22796 32774
rect 22742 32736 22744 32745
rect 22796 32736 22798 32745
rect 22742 32671 22798 32680
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22284 32428 22336 32434
rect 22284 32370 22336 32376
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 21548 32020 21600 32026
rect 21548 31962 21600 31968
rect 22480 31346 22508 32302
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22112 30054 22140 31078
rect 22296 30598 22324 31282
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22480 30410 22508 31282
rect 22572 31278 22600 32370
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22756 30734 22784 32671
rect 23492 32230 23520 32864
rect 23572 32846 23624 32852
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23952 31482 23980 33390
rect 24504 33114 24532 33866
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24596 32910 24624 33050
rect 24032 32904 24084 32910
rect 24032 32846 24084 32852
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 23020 31272 23072 31278
rect 23020 31214 23072 31220
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 22480 30382 22600 30410
rect 22664 30394 22692 30670
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22480 29510 22508 30194
rect 22572 29646 22600 30382
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 23032 30326 23060 31214
rect 23204 30864 23256 30870
rect 23204 30806 23256 30812
rect 23216 30598 23244 30806
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 23492 30598 23520 30670
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 23216 30258 23244 30534
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23296 30048 23348 30054
rect 23296 29990 23348 29996
rect 23112 29776 23164 29782
rect 23112 29718 23164 29724
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22006 28520 22062 28529
rect 22006 28455 22008 28464
rect 22060 28455 22062 28464
rect 22008 28426 22060 28432
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22112 28150 22140 28358
rect 22388 28150 22416 28902
rect 22100 28144 22152 28150
rect 22100 28086 22152 28092
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 21836 25702 21864 26250
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 21824 25696 21876 25702
rect 21824 25638 21876 25644
rect 21732 25356 21784 25362
rect 21928 25344 21956 25978
rect 22112 25498 22140 26250
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 21784 25316 21956 25344
rect 21732 25298 21784 25304
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 22020 24818 22048 25162
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22020 24410 22048 24754
rect 22204 24750 22232 25638
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22112 24410 22140 24686
rect 22296 24614 22324 25910
rect 22284 24608 22336 24614
rect 22284 24550 22336 24556
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21456 21412 21508 21418
rect 21456 21354 21508 21360
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21560 20874 21588 21014
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21652 20262 21680 24074
rect 22020 23186 22048 24210
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22008 23180 22060 23186
rect 22008 23122 22060 23128
rect 22296 23050 22324 23462
rect 22388 23186 22416 26386
rect 22480 24750 22508 29446
rect 23124 29170 23152 29718
rect 23308 29646 23336 29990
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23492 28694 23520 30534
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23584 29102 23612 29582
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23572 29096 23624 29102
rect 23572 29038 23624 29044
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23492 28082 23520 28426
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23584 28014 23612 29038
rect 23676 28762 23704 29242
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23676 27606 23704 28698
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23768 27606 23796 28562
rect 23848 28416 23900 28422
rect 23848 28358 23900 28364
rect 23860 28150 23888 28358
rect 23848 28144 23900 28150
rect 23848 28086 23900 28092
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 22572 26586 22600 26930
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23730 22508 24006
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 22572 22930 22600 25842
rect 22664 24818 22692 26726
rect 22756 25430 22784 26726
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22756 25226 22784 25366
rect 22848 25294 22876 26522
rect 23124 25430 23152 26862
rect 23492 25498 23520 26930
rect 23584 26790 23612 26998
rect 23676 26926 23704 27406
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23584 25974 23612 26726
rect 23952 26042 23980 29446
rect 23940 26036 23992 26042
rect 23940 25978 23992 25984
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 23952 25498 23980 25978
rect 24044 25906 24072 32846
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24228 30190 24256 32370
rect 24688 32230 24716 34002
rect 24768 33856 24820 33862
rect 24768 33798 24820 33804
rect 24780 33318 24808 33798
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 24768 33312 24820 33318
rect 24768 33254 24820 33260
rect 24780 32434 24808 33254
rect 25700 33114 25728 33526
rect 27252 33448 27304 33454
rect 27252 33390 27304 33396
rect 25688 33108 25740 33114
rect 25688 33050 25740 33056
rect 24860 33040 24912 33046
rect 25044 33040 25096 33046
rect 24912 32988 25044 32994
rect 24860 32982 25096 32988
rect 24872 32966 25084 32982
rect 25044 32904 25096 32910
rect 24950 32872 25006 32881
rect 25044 32846 25096 32852
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 24950 32807 24952 32816
rect 25004 32807 25006 32816
rect 24952 32778 25004 32784
rect 25056 32570 25084 32846
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 24768 32428 24820 32434
rect 24768 32370 24820 32376
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24860 31272 24912 31278
rect 24860 31214 24912 31220
rect 24872 30938 24900 31214
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 24768 30660 24820 30666
rect 24768 30602 24820 30608
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24228 30054 24256 30126
rect 24688 30054 24716 30262
rect 24216 30048 24268 30054
rect 24216 29990 24268 29996
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24412 29646 24440 29990
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 24400 29640 24452 29646
rect 24400 29582 24452 29588
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29186 24532 29582
rect 24412 29158 24532 29186
rect 24688 29170 24716 29786
rect 24676 29164 24728 29170
rect 24412 29102 24440 29158
rect 24676 29106 24728 29112
rect 24400 29096 24452 29102
rect 24400 29038 24452 29044
rect 24412 28966 24440 29038
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24216 28688 24268 28694
rect 24216 28630 24268 28636
rect 24228 27282 24256 28630
rect 24412 28558 24440 28902
rect 24688 28762 24716 29106
rect 24780 29102 24808 30602
rect 24964 30394 24992 30670
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 25056 30326 25084 30670
rect 25044 30320 25096 30326
rect 25044 30262 25096 30268
rect 25148 30122 25176 32302
rect 25228 30864 25280 30870
rect 25228 30806 25280 30812
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 25136 30116 25188 30122
rect 25136 30058 25188 30064
rect 24964 29170 24992 30058
rect 25148 29306 25176 30058
rect 25240 29850 25268 30806
rect 25424 30802 25452 32370
rect 26344 32230 26372 32846
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26344 31822 26372 32166
rect 27264 31890 27292 33390
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 27988 32904 28040 32910
rect 27988 32846 28040 32852
rect 27908 32570 27936 32846
rect 28000 32745 28028 32846
rect 27986 32736 28042 32745
rect 27986 32671 28042 32680
rect 27896 32564 27948 32570
rect 27896 32506 27948 32512
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26240 31748 26292 31754
rect 26240 31690 26292 31696
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25608 31414 25636 31622
rect 26252 31482 26280 31690
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24676 28756 24728 28762
rect 24676 28698 24728 28704
rect 24400 28552 24452 28558
rect 24452 28512 24532 28540
rect 24400 28494 24452 28500
rect 24504 28082 24532 28512
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24320 27402 24348 28018
rect 24504 27538 24532 28018
rect 24492 27532 24544 27538
rect 24492 27474 24544 27480
rect 24308 27396 24360 27402
rect 24308 27338 24360 27344
rect 24228 27254 24348 27282
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 23112 25424 23164 25430
rect 23112 25366 23164 25372
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 22744 25220 22796 25226
rect 22744 25162 22796 25168
rect 23308 24954 23336 25230
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23492 24818 23520 25094
rect 24044 24954 24072 25842
rect 24136 25838 24164 26930
rect 24320 26790 24348 27254
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 24320 26586 24348 26726
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24306 26344 24362 26353
rect 24306 26279 24362 26288
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 24320 25226 24348 26279
rect 24308 25220 24360 25226
rect 24308 25162 24360 25168
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22756 23798 22784 24278
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23322 23796 23462
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 22296 22902 22600 22930
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21744 21010 21772 21422
rect 22204 21146 22232 21490
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21744 19922 21772 20946
rect 21824 20936 21876 20942
rect 22008 20936 22060 20942
rect 21876 20884 22008 20890
rect 21824 20878 22060 20884
rect 21836 20862 22048 20878
rect 22020 20058 22048 20862
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21836 17202 21864 18226
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 17678 21956 18022
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 14618 21404 15438
rect 21732 15088 21784 15094
rect 21732 15030 21784 15036
rect 21744 14618 21772 15030
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21836 14414 21864 17138
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 15094 22140 15302
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21284 4214 21312 12718
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21744 4826 21772 5170
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21836 4146 21864 4966
rect 21928 4282 21956 5170
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 22296 4078 22324 22902
rect 23400 22710 23428 23054
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23124 21962 23152 22578
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 22664 21622 22692 21898
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 23400 21554 23428 21898
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 20534 22416 21286
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22480 20466 22508 20742
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22572 20058 22600 21490
rect 23020 21412 23072 21418
rect 23020 21354 23072 21360
rect 23032 21146 23060 21354
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 23768 20534 23796 21286
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22480 19378 22508 19654
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22388 18902 22416 19246
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22480 18086 22508 19314
rect 22572 19310 22600 19994
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18290 22784 18566
rect 23032 18358 23060 19110
rect 23020 18352 23072 18358
rect 23020 18294 23072 18300
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 23662 17912 23718 17921
rect 23662 17847 23718 17856
rect 23676 17270 23704 17847
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 22848 14618 22876 15030
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 23400 13326 23428 16526
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23492 16182 23520 16390
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23584 14482 23612 14758
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 22388 4146 22416 4966
rect 23124 4622 23152 4966
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 22480 4282 22508 4558
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 23124 4146 23152 4422
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22008 3936 22060 3942
rect 22006 3904 22008 3913
rect 22744 3936 22796 3942
rect 22060 3904 22062 3913
rect 22744 3878 22796 3884
rect 22006 3839 22062 3848
rect 22756 3534 22784 3878
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 21836 3058 21864 3470
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 21928 800 21956 3402
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22020 2990 22048 3334
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22204 2446 22232 3334
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22572 800 22600 2926
rect 23216 2446 23244 4966
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23308 1442 23336 4014
rect 23492 3534 23520 5238
rect 23676 4026 23704 17070
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 4146 23796 4422
rect 23860 4146 23888 5170
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23676 3998 23888 4026
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23860 2854 23888 3998
rect 23756 2848 23808 2854
rect 23754 2816 23756 2825
rect 23848 2848 23900 2854
rect 23808 2816 23810 2825
rect 23848 2790 23900 2796
rect 23754 2751 23810 2760
rect 23860 2650 23888 2790
rect 23952 2650 23980 24754
rect 24044 24274 24072 24890
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24412 23662 24440 24006
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24596 23508 24624 28018
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24688 26024 24716 27542
rect 24780 27470 24808 29038
rect 24964 28762 24992 29106
rect 24952 28756 25004 28762
rect 24952 28698 25004 28704
rect 24964 28626 24992 28698
rect 25148 28694 25176 29242
rect 25136 28688 25188 28694
rect 25136 28630 25188 28636
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24964 28014 24992 28562
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25240 28218 25268 28494
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24688 25996 24808 26024
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24688 24682 24716 25842
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24412 23480 24624 23508
rect 24412 19922 24440 23480
rect 24780 22094 24808 25996
rect 24872 25906 24900 26930
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24872 25430 24900 25842
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24872 24954 24900 25366
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 24964 24614 24992 26250
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25148 25265 25176 25842
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25148 24886 25176 25191
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24596 22066 24808 22094
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24504 20534 24532 20742
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24596 19378 24624 22066
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25148 20602 25176 20810
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25240 20058 25268 28018
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18766 24440 19110
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24412 18222 24440 18702
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18358 24532 18566
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24688 6914 24716 19790
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24780 17202 24808 18566
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 25148 6914 25176 19722
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25240 16522 25268 17138
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 25240 15434 25268 16458
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 24320 6886 24716 6914
rect 24964 6886 25176 6914
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24320 2514 24348 6886
rect 24676 4004 24728 4010
rect 24676 3946 24728 3952
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24504 2514 24532 3878
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24596 3058 24624 3538
rect 24688 3534 24716 3946
rect 24872 3913 24900 3946
rect 24858 3904 24914 3913
rect 24858 3839 24914 3848
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24780 3126 24808 3334
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24872 2922 24900 3334
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24964 2825 24992 6886
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24950 2816 25006 2825
rect 24950 2751 25006 2760
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 24492 2508 24544 2514
rect 24492 2450 24544 2456
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 23216 1414 23336 1442
rect 23216 800 23244 1414
rect 24504 800 24532 2246
rect 25148 800 25176 2926
rect 25240 2922 25268 15370
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 25332 2582 25360 30670
rect 25424 30666 25452 30738
rect 25688 30728 25740 30734
rect 25688 30670 25740 30676
rect 25412 30660 25464 30666
rect 25412 30602 25464 30608
rect 25700 30258 25728 30670
rect 25976 30258 26004 31078
rect 26148 30864 26200 30870
rect 26148 30806 26200 30812
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25424 27674 25452 29990
rect 25700 28966 25728 30194
rect 26160 30054 26188 30806
rect 26148 30048 26200 30054
rect 26148 29990 26200 29996
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26252 29034 26280 29650
rect 26344 29646 26372 31758
rect 27264 29714 27292 31826
rect 27988 31748 28040 31754
rect 27988 31690 28040 31696
rect 28000 31482 28028 31690
rect 27988 31476 28040 31482
rect 27988 31418 28040 31424
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27632 30938 27660 31282
rect 27908 30938 27936 31282
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 27252 29708 27304 29714
rect 27252 29650 27304 29656
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26344 29170 26372 29582
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 26608 29504 26660 29510
rect 26608 29446 26660 29452
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 26240 29028 26292 29034
rect 26240 28970 26292 28976
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 26252 28626 26280 28970
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25516 28218 25544 28426
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25516 27674 25544 28018
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 25412 27668 25464 27674
rect 25412 27610 25464 27616
rect 25504 27668 25556 27674
rect 25504 27610 25556 27616
rect 25424 26382 25452 27610
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25976 26314 26004 26726
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25792 25809 25820 25842
rect 25778 25800 25834 25809
rect 25778 25735 25834 25744
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24274 25912 24754
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25608 23186 25636 24006
rect 25884 23798 25912 24210
rect 25976 24206 26004 25638
rect 26252 25498 26280 27882
rect 26344 27470 26372 29106
rect 26620 28558 26648 29446
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27356 29170 27384 29242
rect 27436 29232 27488 29238
rect 27436 29174 27488 29180
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26436 26314 26464 27270
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26240 25492 26292 25498
rect 26240 25434 26292 25440
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26252 24750 26280 25298
rect 26804 25294 26832 26182
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 26344 24698 26372 24754
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26068 23866 26096 24142
rect 26160 24070 26188 24550
rect 26252 24410 26280 24686
rect 26344 24670 26464 24698
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26344 24138 26372 24550
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26436 23866 26464 24670
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 26148 23724 26200 23730
rect 26332 23724 26384 23730
rect 26200 23684 26280 23712
rect 26148 23666 26200 23672
rect 26252 23610 26280 23684
rect 26436 23712 26464 23802
rect 26384 23684 26464 23712
rect 26332 23666 26384 23672
rect 26528 23610 26556 24550
rect 26252 23582 26556 23610
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26344 22710 26372 22986
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 26160 21554 26188 22578
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26436 21554 26464 21830
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 25424 20874 25452 21286
rect 25412 20868 25464 20874
rect 25412 20810 25464 20816
rect 26068 20466 26096 21286
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 25976 20058 26004 20402
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26528 18834 26556 23582
rect 26804 23186 26832 25230
rect 26896 24290 26924 25434
rect 26976 24336 27028 24342
rect 26896 24284 26976 24290
rect 26896 24278 27028 24284
rect 26896 24262 27016 24278
rect 26896 24206 26924 24262
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26792 23180 26844 23186
rect 26792 23122 26844 23128
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26804 22386 26832 22510
rect 26896 22506 26924 23802
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26988 23322 27016 23666
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 27080 23202 27108 29106
rect 27448 28370 27476 29174
rect 27540 29170 27568 29514
rect 27632 29322 27660 30874
rect 27804 30116 27856 30122
rect 27804 30058 27856 30064
rect 27816 29510 27844 30058
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27632 29294 27752 29322
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27540 28490 27568 29106
rect 27724 28558 27752 29294
rect 27816 28626 27844 29446
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27804 28620 27856 28626
rect 27804 28562 27856 28568
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27448 28342 27660 28370
rect 27632 28082 27660 28342
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 27172 26042 27200 26930
rect 27252 26444 27304 26450
rect 27252 26386 27304 26392
rect 27160 26036 27212 26042
rect 27160 25978 27212 25984
rect 27160 25832 27212 25838
rect 27160 25774 27212 25780
rect 27172 25498 27200 25774
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 27264 24750 27292 26386
rect 27344 25900 27396 25906
rect 27344 25842 27396 25848
rect 27356 25702 27384 25842
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27632 24818 27660 28018
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27528 24744 27580 24750
rect 27528 24686 27580 24692
rect 27540 23730 27568 24686
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 26988 23174 27108 23202
rect 26884 22500 26936 22506
rect 26884 22442 26936 22448
rect 26988 22386 27016 23174
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27080 22642 27108 22986
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 26804 22358 27016 22386
rect 26988 22098 27016 22358
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26608 22024 26660 22030
rect 27080 21978 27108 22578
rect 27344 22500 27396 22506
rect 27344 22442 27396 22448
rect 26660 21972 27108 21978
rect 26608 21966 27108 21972
rect 26620 21956 27108 21966
rect 26620 21950 26976 21956
rect 26620 20806 26648 21950
rect 27028 21950 27108 21956
rect 26976 21898 27028 21904
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27172 21690 27200 21830
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27264 21486 27292 21830
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26620 20534 26648 20742
rect 27356 20534 27384 22442
rect 27540 21486 27568 23666
rect 27724 23202 27752 28494
rect 27816 26994 27844 28562
rect 27896 27668 27948 27674
rect 27896 27610 27948 27616
rect 27908 27130 27936 27610
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27804 26988 27856 26994
rect 27804 26930 27856 26936
rect 27816 25974 27844 26930
rect 27804 25968 27856 25974
rect 27804 25910 27856 25916
rect 27632 23174 27752 23202
rect 27632 22710 27660 23174
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27724 22574 27752 23054
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27724 22030 27752 22510
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27724 21570 27752 21966
rect 27724 21542 27844 21570
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27540 21010 27568 21422
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27632 20058 27660 20878
rect 27724 20602 27752 20878
rect 27816 20874 27844 21542
rect 27908 20942 27936 27066
rect 28000 26042 28028 29106
rect 27988 26036 28040 26042
rect 27988 25978 28040 25984
rect 28092 25786 28120 40394
rect 28172 33448 28224 33454
rect 28172 33390 28224 33396
rect 28184 33114 28212 33390
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 28448 32904 28500 32910
rect 28448 32846 28500 32852
rect 28460 32774 28488 32846
rect 28448 32768 28500 32774
rect 28262 32736 28318 32745
rect 28448 32710 28500 32716
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 28262 32671 28318 32680
rect 28276 30818 28304 32671
rect 28460 31346 28488 32710
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28552 31482 28580 31826
rect 28540 31476 28592 31482
rect 28540 31418 28592 31424
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28368 30938 28396 31282
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 28276 30790 28396 30818
rect 28264 30048 28316 30054
rect 28264 29990 28316 29996
rect 28276 29170 28304 29990
rect 28264 29164 28316 29170
rect 28264 29106 28316 29112
rect 28368 29102 28396 30790
rect 28356 29096 28408 29102
rect 28356 29038 28408 29044
rect 28368 28422 28396 29038
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28460 26353 28488 31282
rect 28644 30122 28672 32370
rect 28828 32230 28856 32710
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 29012 30870 29040 31078
rect 29000 30864 29052 30870
rect 29000 30806 29052 30812
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 29012 30598 29040 30670
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 29012 30258 29040 30534
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 29000 30116 29052 30122
rect 29000 30058 29052 30064
rect 29012 29850 29040 30058
rect 28724 29844 28776 29850
rect 28724 29786 28776 29792
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28552 28762 28580 29514
rect 28736 29306 28764 29786
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 28828 29102 28856 29242
rect 29012 29170 29040 29786
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 28816 29096 28868 29102
rect 28816 29038 28868 29044
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28540 28756 28592 28762
rect 28540 28698 28592 28704
rect 28828 28626 28856 28902
rect 28816 28620 28868 28626
rect 28816 28562 28868 28568
rect 28446 26344 28502 26353
rect 28446 26279 28502 26288
rect 28724 25968 28776 25974
rect 28724 25910 28776 25916
rect 28000 25758 28120 25786
rect 28000 24614 28028 25758
rect 28080 25696 28132 25702
rect 28080 25638 28132 25644
rect 28092 25498 28120 25638
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 28632 25220 28684 25226
rect 28632 25162 28684 25168
rect 28644 24818 28672 25162
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28172 22704 28224 22710
rect 28172 22646 28224 22652
rect 27988 22160 28040 22166
rect 27988 22102 28040 22108
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 28000 20466 28028 22102
rect 28184 22030 28212 22646
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28552 21622 28580 21830
rect 28540 21616 28592 21622
rect 28540 21558 28592 21564
rect 28264 21480 28316 21486
rect 28264 21422 28316 21428
rect 28276 21146 28304 21422
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28356 21140 28408 21146
rect 28356 21082 28408 21088
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 28092 20398 28120 20878
rect 28368 20806 28396 21082
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25516 17678 25544 18226
rect 25700 17678 25728 18362
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 25516 17134 25544 17614
rect 25700 17202 25728 17614
rect 26436 17202 26464 17614
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 25424 16454 25452 16934
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25976 16590 26004 16662
rect 26160 16590 26188 16934
rect 27080 16658 27108 17614
rect 27172 17202 27200 18022
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25424 15502 25452 16390
rect 25976 16250 26004 16526
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 25516 15706 25544 16186
rect 26160 16114 26188 16526
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25424 2774 25452 15438
rect 26252 15162 26280 16186
rect 26344 15502 26372 16390
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26528 14958 26556 16186
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27080 15162 27108 16050
rect 27160 15972 27212 15978
rect 27160 15914 27212 15920
rect 27172 15502 27200 15914
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 26344 3534 26372 3606
rect 26804 3602 26832 14894
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 25424 2746 25544 2774
rect 25228 2576 25280 2582
rect 25228 2518 25280 2524
rect 25320 2576 25372 2582
rect 25320 2518 25372 2524
rect 25240 2106 25268 2518
rect 25516 2514 25544 2746
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25228 2100 25280 2106
rect 25228 2042 25280 2048
rect 26436 800 26464 3470
rect 27540 3398 27568 18770
rect 27632 18358 27660 19110
rect 28172 18896 28224 18902
rect 28172 18838 28224 18844
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27724 15706 27752 18634
rect 28184 18222 28212 18838
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 28172 18216 28224 18222
rect 28172 18158 28224 18164
rect 28092 17610 28120 18158
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 27804 16108 27856 16114
rect 27804 16050 27856 16056
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27724 14958 27752 15642
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27816 14890 27844 16050
rect 27804 14884 27856 14890
rect 27804 14826 27856 14832
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27540 2990 27568 3334
rect 28092 3058 28120 17546
rect 28276 17338 28304 18702
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26896 2446 26924 2586
rect 28460 2514 28488 19790
rect 28736 5098 28764 25910
rect 28828 24614 28856 28562
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28828 24410 28856 24550
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28828 23594 28856 24346
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 28920 23322 28948 28902
rect 29000 26784 29052 26790
rect 29000 26726 29052 26732
rect 29012 25906 29040 26726
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28920 20874 28948 21286
rect 28908 20868 28960 20874
rect 28908 20810 28960 20816
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 29012 20466 29040 20742
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29104 18630 29132 47126
rect 29656 47054 29684 49200
rect 30760 47122 30788 49286
rect 30902 49200 31014 49286
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36698 49200 36810 50000
rect 37342 49200 37454 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 39918 49314 40030 50000
rect 39592 49286 40030 49314
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 31116 47048 31168 47054
rect 31116 46990 31168 46996
rect 29368 46504 29420 46510
rect 29368 46446 29420 46452
rect 29184 31680 29236 31686
rect 29184 31622 29236 31628
rect 29196 31278 29224 31622
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29184 31272 29236 31278
rect 29184 31214 29236 31220
rect 29196 30666 29224 31214
rect 29288 30870 29316 31282
rect 29276 30864 29328 30870
rect 29276 30806 29328 30812
rect 29184 30660 29236 30666
rect 29184 30602 29236 30608
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 29196 26926 29224 28426
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 29196 21962 29224 26862
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29196 21842 29224 21898
rect 29196 21814 29316 21842
rect 29184 21684 29236 21690
rect 29184 21626 29236 21632
rect 29196 21078 29224 21626
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 29288 20602 29316 21814
rect 29276 20596 29328 20602
rect 29276 20538 29328 20544
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 29196 19922 29224 20402
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 28724 5092 28776 5098
rect 28724 5034 28776 5040
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27080 800 27108 2314
rect 28368 800 28396 2382
rect 29288 2106 29316 20402
rect 29380 4078 29408 46446
rect 30564 34604 30616 34610
rect 30564 34546 30616 34552
rect 29644 34536 29696 34542
rect 29644 34478 29696 34484
rect 29656 33590 29684 34478
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 30392 33930 30420 34342
rect 30380 33924 30432 33930
rect 30380 33866 30432 33872
rect 29644 33584 29696 33590
rect 29644 33526 29696 33532
rect 29920 33516 29972 33522
rect 29920 33458 29972 33464
rect 29828 33448 29880 33454
rect 29828 33390 29880 33396
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29656 32978 29684 33254
rect 29644 32972 29696 32978
rect 29644 32914 29696 32920
rect 29656 32366 29684 32914
rect 29748 32434 29776 33254
rect 29840 32910 29868 33390
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29644 31136 29696 31142
rect 29644 31078 29696 31084
rect 29656 28558 29684 31078
rect 29736 30728 29788 30734
rect 29736 30670 29788 30676
rect 29748 29510 29776 30670
rect 29840 29646 29868 32846
rect 29932 32230 29960 33458
rect 30576 33114 30604 34546
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30564 33108 30616 33114
rect 30564 33050 30616 33056
rect 30852 32978 30880 33254
rect 31128 33046 31156 46990
rect 32232 46442 32260 49200
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 32312 46504 32364 46510
rect 32312 46446 32364 46452
rect 32220 46436 32272 46442
rect 32220 46378 32272 46384
rect 32324 46170 32352 46446
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 32312 46164 32364 46170
rect 32312 46106 32364 46112
rect 31760 45960 31812 45966
rect 31760 45902 31812 45908
rect 31772 41614 31800 45902
rect 38028 45554 38056 49200
rect 38108 47048 38160 47054
rect 38108 46990 38160 46996
rect 38120 46578 38148 46990
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 38672 46510 38700 49200
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38292 46504 38344 46510
rect 38292 46446 38344 46452
rect 38660 46504 38712 46510
rect 38660 46446 38712 46452
rect 38304 46170 38332 46446
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 39592 45554 39620 49286
rect 39918 49200 40030 49286
rect 40562 49200 40674 50000
rect 41206 49200 41318 50000
rect 41850 49200 41962 50000
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 43782 49200 43894 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 45714 49200 45826 50000
rect 46358 49200 46470 50000
rect 47002 49200 47114 50000
rect 47646 49200 47758 50000
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 41248 47462 41276 49200
rect 40040 47456 40092 47462
rect 40040 47398 40092 47404
rect 41236 47456 41288 47462
rect 41236 47398 41288 47404
rect 37292 45526 38056 45554
rect 38856 45526 39620 45554
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 31760 41608 31812 41614
rect 31760 41550 31812 41556
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 31760 34536 31812 34542
rect 31760 34478 31812 34484
rect 31668 33856 31720 33862
rect 31668 33798 31720 33804
rect 31680 33522 31708 33798
rect 31668 33516 31720 33522
rect 31668 33458 31720 33464
rect 31116 33040 31168 33046
rect 31116 32982 31168 32988
rect 30840 32972 30892 32978
rect 30840 32914 30892 32920
rect 31680 32910 31708 33458
rect 31772 32910 31800 34478
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 32220 34060 32272 34066
rect 32220 34002 32272 34008
rect 31852 33924 31904 33930
rect 31852 33866 31904 33872
rect 31864 33114 31892 33866
rect 32128 33448 32180 33454
rect 32128 33390 32180 33396
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 31944 33108 31996 33114
rect 31944 33050 31996 33056
rect 30012 32904 30064 32910
rect 30012 32846 30064 32852
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 30024 32434 30052 32846
rect 30012 32428 30064 32434
rect 30012 32370 30064 32376
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29644 28552 29696 28558
rect 29696 28512 29776 28540
rect 29644 28494 29696 28500
rect 29644 27940 29696 27946
rect 29644 27882 29696 27888
rect 29656 26994 29684 27882
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29552 26036 29604 26042
rect 29552 25978 29604 25984
rect 29460 25900 29512 25906
rect 29460 25842 29512 25848
rect 29472 24954 29500 25842
rect 29460 24948 29512 24954
rect 29460 24890 29512 24896
rect 29472 24206 29500 24890
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29564 22094 29592 25978
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 29472 22066 29592 22094
rect 29472 21894 29500 22066
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29472 20398 29500 21830
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29656 6914 29684 25842
rect 29748 25430 29776 28512
rect 29840 28082 29868 29582
rect 29932 28082 29960 32166
rect 31772 31822 31800 32846
rect 31956 32570 31984 33050
rect 32036 32768 32088 32774
rect 32036 32710 32088 32716
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 32048 32298 32076 32710
rect 32140 32366 32168 33390
rect 32232 32434 32260 34002
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 37292 33114 37320 45526
rect 38476 45280 38528 45286
rect 38476 45222 38528 45228
rect 37280 33108 37332 33114
rect 37280 33050 37332 33056
rect 35072 33040 35124 33046
rect 35072 32982 35124 32988
rect 37464 33040 37516 33046
rect 37464 32982 37516 32988
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 32036 32292 32088 32298
rect 32036 32234 32088 32240
rect 32048 31890 32076 32234
rect 32232 31958 32260 32370
rect 32784 32026 32812 32846
rect 33416 32768 33468 32774
rect 33416 32710 33468 32716
rect 33428 32570 33456 32710
rect 33416 32564 33468 32570
rect 33416 32506 33468 32512
rect 34060 32496 34112 32502
rect 34060 32438 34112 32444
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 32772 32020 32824 32026
rect 32772 31962 32824 31968
rect 32220 31952 32272 31958
rect 32220 31894 32272 31900
rect 32036 31884 32088 31890
rect 32036 31826 32088 31832
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31024 31680 31076 31686
rect 31024 31622 31076 31628
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30012 30660 30064 30666
rect 30012 30602 30064 30608
rect 30024 30054 30052 30602
rect 30116 30326 30144 30874
rect 31036 30734 31064 31622
rect 31668 30796 31720 30802
rect 31668 30738 31720 30744
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 30104 30320 30156 30326
rect 30104 30262 30156 30268
rect 31036 30190 31064 30670
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 31024 30184 31076 30190
rect 31024 30126 31076 30132
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30564 30048 30616 30054
rect 30564 29990 30616 29996
rect 30576 29238 30604 29990
rect 31128 29850 31156 30194
rect 31484 30048 31536 30054
rect 31484 29990 31536 29996
rect 31116 29844 31168 29850
rect 31116 29786 31168 29792
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 30748 29640 30800 29646
rect 30748 29582 30800 29588
rect 30564 29232 30616 29238
rect 30564 29174 30616 29180
rect 30760 29102 30788 29582
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30748 29096 30800 29102
rect 30748 29038 30800 29044
rect 30472 29028 30524 29034
rect 30472 28970 30524 28976
rect 30484 28558 30512 28970
rect 30760 28626 30788 29038
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 30852 28762 30880 28902
rect 30840 28756 30892 28762
rect 30840 28698 30892 28704
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30944 28490 30972 29106
rect 31036 28762 31064 29650
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 30196 28484 30248 28490
rect 30196 28426 30248 28432
rect 30932 28484 30984 28490
rect 30932 28426 30984 28432
rect 29828 28076 29880 28082
rect 29828 28018 29880 28024
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29932 27962 29960 28018
rect 29840 27934 29960 27962
rect 29840 27878 29868 27934
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 29920 27396 29972 27402
rect 29920 27338 29972 27344
rect 29828 26308 29880 26314
rect 29828 26250 29880 26256
rect 29840 26042 29868 26250
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 29736 25424 29788 25430
rect 29736 25366 29788 25372
rect 29932 24682 29960 27338
rect 30208 27334 30236 28426
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 30208 27062 30236 27270
rect 30392 27062 30420 28154
rect 31128 28082 31156 29786
rect 31496 29646 31524 29990
rect 31680 29850 31708 30738
rect 31944 30320 31996 30326
rect 31944 30262 31996 30268
rect 31668 29844 31720 29850
rect 31668 29786 31720 29792
rect 31956 29714 31984 30262
rect 32232 30190 32260 31894
rect 32496 31884 32548 31890
rect 32496 31826 32548 31832
rect 32220 30184 32272 30190
rect 32220 30126 32272 30132
rect 31944 29708 31996 29714
rect 31944 29650 31996 29656
rect 31484 29640 31536 29646
rect 31484 29582 31536 29588
rect 31484 28620 31536 28626
rect 31484 28562 31536 28568
rect 31208 28212 31260 28218
rect 31208 28154 31260 28160
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31024 28008 31076 28014
rect 31024 27950 31076 27956
rect 31036 27878 31064 27950
rect 31220 27878 31248 28154
rect 31392 28144 31444 28150
rect 31392 28086 31444 28092
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 31208 27872 31260 27878
rect 31208 27814 31260 27820
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31036 27674 31064 27814
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 30196 27056 30248 27062
rect 30196 26998 30248 27004
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 30392 26466 30420 26998
rect 30300 26438 30420 26466
rect 31036 26450 31064 27610
rect 31312 27130 31340 27814
rect 31404 27606 31432 28086
rect 31496 27606 31524 28562
rect 31956 28558 31984 29650
rect 32404 28960 32456 28966
rect 32404 28902 32456 28908
rect 32416 28762 32444 28902
rect 32404 28756 32456 28762
rect 32404 28698 32456 28704
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 32128 28552 32180 28558
rect 32128 28494 32180 28500
rect 31864 28422 31892 28494
rect 31956 28422 31984 28494
rect 31852 28416 31904 28422
rect 31852 28358 31904 28364
rect 31944 28416 31996 28422
rect 31944 28358 31996 28364
rect 31576 28008 31628 28014
rect 31576 27950 31628 27956
rect 31392 27600 31444 27606
rect 31392 27542 31444 27548
rect 31484 27600 31536 27606
rect 31484 27542 31536 27548
rect 31588 27538 31616 27950
rect 31576 27532 31628 27538
rect 31576 27474 31628 27480
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 31024 26444 31076 26450
rect 30196 26036 30248 26042
rect 30300 26024 30328 26438
rect 31024 26386 31076 26392
rect 30380 26308 30432 26314
rect 30380 26250 30432 26256
rect 30392 26042 30420 26250
rect 30248 25996 30328 26024
rect 30380 26036 30432 26042
rect 30196 25978 30248 25984
rect 30380 25978 30432 25984
rect 31036 25838 31064 26386
rect 31312 25838 31340 27066
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 31772 26314 31800 26522
rect 31760 26308 31812 26314
rect 31760 26250 31812 26256
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30116 24818 30144 25230
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 30300 24834 30328 24890
rect 31312 24886 31340 25774
rect 31300 24880 31352 24886
rect 30300 24818 30512 24834
rect 31300 24822 31352 24828
rect 30104 24812 30156 24818
rect 30300 24812 30524 24818
rect 30300 24806 30472 24812
rect 30104 24754 30156 24760
rect 30472 24754 30524 24760
rect 29920 24676 29972 24682
rect 29920 24618 29972 24624
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 30024 24206 30052 24550
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29840 23798 29868 24006
rect 29828 23792 29880 23798
rect 29828 23734 29880 23740
rect 30010 23624 30066 23633
rect 30116 23610 30144 24754
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 31760 24744 31812 24750
rect 31760 24686 31812 24692
rect 30208 23662 30236 24686
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 30656 24404 30708 24410
rect 30656 24346 30708 24352
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30066 23582 30144 23610
rect 30196 23656 30248 23662
rect 30196 23598 30248 23604
rect 30010 23559 30066 23568
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29736 21956 29788 21962
rect 29736 21898 29788 21904
rect 29748 21622 29776 21898
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29840 20602 29868 21966
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 30024 19854 30052 23559
rect 30300 23322 30328 24142
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30116 21894 30144 21966
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 30392 21010 30420 23122
rect 30668 23118 30696 24346
rect 30748 24336 30800 24342
rect 30748 24278 30800 24284
rect 30760 24070 30788 24278
rect 31312 24206 31340 24550
rect 31300 24200 31352 24206
rect 31300 24142 31352 24148
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 30748 24064 30800 24070
rect 30746 24032 30748 24041
rect 31300 24064 31352 24070
rect 30800 24032 30802 24041
rect 31300 24006 31352 24012
rect 30746 23967 30802 23976
rect 31312 23866 31340 24006
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31128 23662 31156 23802
rect 31208 23792 31260 23798
rect 31208 23734 31260 23740
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31220 23322 31248 23734
rect 31208 23316 31260 23322
rect 31208 23258 31260 23264
rect 31680 23186 31708 24074
rect 31772 23526 31800 24686
rect 31864 23866 31892 28358
rect 31956 28218 31984 28358
rect 31944 28212 31996 28218
rect 31944 28154 31996 28160
rect 32140 27418 32168 28494
rect 32220 28076 32272 28082
rect 32220 28018 32272 28024
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32232 27538 32260 28018
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32036 27396 32088 27402
rect 32140 27390 32260 27418
rect 32036 27338 32088 27344
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 31956 26518 31984 26862
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 31956 25906 31984 26318
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 31956 25294 31984 25842
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 31956 24750 31984 25230
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 32048 24562 32076 27338
rect 32128 26852 32180 26858
rect 32128 26794 32180 26800
rect 32140 26489 32168 26794
rect 32126 26480 32182 26489
rect 32126 26415 32182 26424
rect 31956 24534 32076 24562
rect 31956 24410 31984 24534
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 32232 24290 32260 27390
rect 32324 25430 32352 28018
rect 32404 25696 32456 25702
rect 32404 25638 32456 25644
rect 32312 25424 32364 25430
rect 32312 25366 32364 25372
rect 32416 25362 32444 25638
rect 32508 25362 32536 31826
rect 33244 31754 33272 32166
rect 33232 31748 33284 31754
rect 33232 31690 33284 31696
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32968 30598 32996 30670
rect 32956 30592 33008 30598
rect 32956 30534 33008 30540
rect 32680 30184 32732 30190
rect 32680 30126 32732 30132
rect 32692 29170 32720 30126
rect 32864 30048 32916 30054
rect 32864 29990 32916 29996
rect 32876 29646 32904 29990
rect 32864 29640 32916 29646
rect 32864 29582 32916 29588
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32956 29504 33008 29510
rect 32956 29446 33008 29452
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32680 28552 32732 28558
rect 32680 28494 32732 28500
rect 32588 27464 32640 27470
rect 32588 27406 32640 27412
rect 32600 26926 32628 27406
rect 32588 26920 32640 26926
rect 32588 26862 32640 26868
rect 32600 26450 32628 26862
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32692 26353 32720 28494
rect 32678 26344 32734 26353
rect 32678 26279 32734 26288
rect 32588 25968 32640 25974
rect 32588 25910 32640 25916
rect 32404 25356 32456 25362
rect 32404 25298 32456 25304
rect 32496 25356 32548 25362
rect 32496 25298 32548 25304
rect 32496 24948 32548 24954
rect 32496 24890 32548 24896
rect 32312 24744 32364 24750
rect 32312 24686 32364 24692
rect 32324 24614 32352 24686
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32048 24262 32260 24290
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 31864 23322 31892 23666
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 30472 23112 30524 23118
rect 30472 23054 30524 23060
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30484 22098 30512 23054
rect 30472 22092 30524 22098
rect 30472 22034 30524 22040
rect 30484 21350 30512 22034
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30484 20942 30512 21286
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30012 19848 30064 19854
rect 30012 19790 30064 19796
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30668 18426 30696 18634
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30576 14482 30604 15302
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 29564 6886 29684 6914
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29276 2100 29328 2106
rect 29276 2042 29328 2048
rect 29564 2038 29592 6886
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 30024 2514 30052 5102
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29552 2032 29604 2038
rect 29552 1974 29604 1980
rect 29656 800 29684 2382
rect 30944 800 30972 3334
rect 32048 2514 32076 24262
rect 32416 24206 32444 24550
rect 32404 24200 32456 24206
rect 32404 24142 32456 24148
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32140 23730 32168 24006
rect 32508 23866 32536 24890
rect 32312 23860 32364 23866
rect 32312 23802 32364 23808
rect 32496 23860 32548 23866
rect 32496 23802 32548 23808
rect 32324 23746 32352 23802
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32232 23718 32352 23746
rect 32232 23594 32260 23718
rect 32220 23588 32272 23594
rect 32220 23530 32272 23536
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32416 22710 32444 23462
rect 32404 22704 32456 22710
rect 32404 22646 32456 22652
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32140 22098 32168 22510
rect 32128 22092 32180 22098
rect 32600 22094 32628 25910
rect 32692 23730 32720 26279
rect 32784 24206 32812 29446
rect 32968 28626 32996 29446
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 33060 28558 33088 29038
rect 33048 28552 33100 28558
rect 33048 28494 33100 28500
rect 33048 26784 33100 26790
rect 33048 26726 33100 26732
rect 33060 26450 33088 26726
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33060 25702 33088 26386
rect 33048 25696 33100 25702
rect 33048 25638 33100 25644
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32876 24342 32904 24754
rect 32968 24614 32996 25230
rect 32956 24608 33008 24614
rect 32956 24550 33008 24556
rect 32864 24336 32916 24342
rect 32864 24278 32916 24284
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32864 23724 32916 23730
rect 32864 23666 32916 23672
rect 32876 23633 32904 23666
rect 32862 23624 32918 23633
rect 32862 23559 32918 23568
rect 32772 22160 32824 22166
rect 32772 22102 32824 22108
rect 32128 22034 32180 22040
rect 32508 22066 32628 22094
rect 32140 21690 32168 22034
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32508 18970 32536 22066
rect 32784 21554 32812 22102
rect 33060 22098 33088 25638
rect 33140 25424 33192 25430
rect 33140 25366 33192 25372
rect 33152 24818 33180 25366
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33244 23118 33272 29582
rect 33336 27334 33364 31690
rect 33888 31686 33916 32166
rect 34072 32026 34100 32438
rect 35084 32434 35112 32982
rect 36544 32972 36596 32978
rect 36544 32914 36596 32920
rect 36176 32904 36228 32910
rect 36228 32852 36308 32858
rect 36176 32846 36308 32852
rect 36188 32830 36308 32846
rect 36176 32768 36228 32774
rect 36176 32710 36228 32716
rect 36188 32570 36216 32710
rect 36176 32564 36228 32570
rect 36176 32506 36228 32512
rect 35072 32428 35124 32434
rect 35072 32370 35124 32376
rect 34520 32360 34572 32366
rect 34520 32302 34572 32308
rect 36176 32360 36228 32366
rect 36176 32302 36228 32308
rect 34060 32020 34112 32026
rect 34060 31962 34112 31968
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33600 31680 33652 31686
rect 33600 31622 33652 31628
rect 33876 31680 33928 31686
rect 33876 31622 33928 31628
rect 33612 31346 33640 31622
rect 33600 31340 33652 31346
rect 33600 31282 33652 31288
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33520 30938 33548 31214
rect 33508 30932 33560 30938
rect 33508 30874 33560 30880
rect 33508 30184 33560 30190
rect 33508 30126 33560 30132
rect 33520 29782 33548 30126
rect 33508 29776 33560 29782
rect 33508 29718 33560 29724
rect 33520 28762 33548 29718
rect 33980 29646 34008 31758
rect 34532 31278 34560 32302
rect 36084 32224 36136 32230
rect 36084 32166 36136 32172
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 36096 31890 36124 32166
rect 36084 31884 36136 31890
rect 36084 31826 36136 31832
rect 36188 31482 36216 32302
rect 36280 32026 36308 32830
rect 36360 32360 36412 32366
rect 36360 32302 36412 32308
rect 36268 32020 36320 32026
rect 36268 31962 36320 31968
rect 36176 31476 36228 31482
rect 36176 31418 36228 31424
rect 36176 31340 36228 31346
rect 36176 31282 36228 31288
rect 34520 31272 34572 31278
rect 34520 31214 34572 31220
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 36188 30938 36216 31282
rect 36176 30932 36228 30938
rect 36176 30874 36228 30880
rect 34520 30796 34572 30802
rect 34520 30738 34572 30744
rect 34244 30320 34296 30326
rect 34244 30262 34296 30268
rect 34256 29850 34284 30262
rect 34532 30054 34560 30738
rect 36280 30734 36308 31962
rect 36268 30728 36320 30734
rect 36268 30670 36320 30676
rect 34796 30592 34848 30598
rect 34796 30534 34848 30540
rect 34520 30048 34572 30054
rect 34520 29990 34572 29996
rect 34244 29844 34296 29850
rect 34244 29786 34296 29792
rect 34532 29714 34560 29990
rect 34520 29708 34572 29714
rect 34520 29650 34572 29656
rect 34808 29646 34836 30534
rect 35348 30184 35400 30190
rect 35348 30126 35400 30132
rect 35992 30184 36044 30190
rect 35992 30126 36044 30132
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 35360 29850 35388 30126
rect 35440 30116 35492 30122
rect 35440 30058 35492 30064
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35452 29714 35480 30058
rect 36004 29850 36032 30126
rect 35992 29844 36044 29850
rect 35992 29786 36044 29792
rect 36084 29844 36136 29850
rect 36084 29786 36136 29792
rect 35440 29708 35492 29714
rect 35440 29650 35492 29656
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 34624 29102 34652 29582
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 34612 29096 34664 29102
rect 34612 29038 34664 29044
rect 34808 29034 34836 29106
rect 34796 29028 34848 29034
rect 34796 28970 34848 28976
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33520 27946 33548 28426
rect 33508 27940 33560 27946
rect 33508 27882 33560 27888
rect 33416 27872 33468 27878
rect 33416 27814 33468 27820
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 33428 27130 33456 27814
rect 33416 27124 33468 27130
rect 33416 27066 33468 27072
rect 33520 25974 33548 27882
rect 33796 27538 33824 28698
rect 34808 27606 34836 28970
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35360 28558 35388 29106
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 35360 28218 35388 28358
rect 35348 28212 35400 28218
rect 35348 28154 35400 28160
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27600 34848 27606
rect 34796 27542 34848 27548
rect 33784 27532 33836 27538
rect 33784 27474 33836 27480
rect 33968 27464 34020 27470
rect 33968 27406 34020 27412
rect 33692 27328 33744 27334
rect 33692 27270 33744 27276
rect 33704 27146 33732 27270
rect 33704 27118 33916 27146
rect 33600 26852 33652 26858
rect 33600 26794 33652 26800
rect 33612 26586 33640 26794
rect 33600 26580 33652 26586
rect 33600 26522 33652 26528
rect 33704 26382 33732 27118
rect 33784 27056 33836 27062
rect 33784 26998 33836 27004
rect 33796 26586 33824 26998
rect 33888 26994 33916 27118
rect 33876 26988 33928 26994
rect 33876 26930 33928 26936
rect 33784 26580 33836 26586
rect 33784 26522 33836 26528
rect 33692 26376 33744 26382
rect 33692 26318 33744 26324
rect 33508 25968 33560 25974
rect 33508 25910 33560 25916
rect 33704 25906 33732 26318
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33692 25696 33744 25702
rect 33692 25638 33744 25644
rect 33704 25362 33732 25638
rect 33692 25356 33744 25362
rect 33692 25298 33744 25304
rect 33508 24948 33560 24954
rect 33508 24890 33560 24896
rect 33520 24138 33548 24890
rect 33704 24818 33732 25298
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33508 24132 33560 24138
rect 33508 24074 33560 24080
rect 33888 23662 33916 24142
rect 33876 23656 33928 23662
rect 33876 23598 33928 23604
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33140 22976 33192 22982
rect 33140 22918 33192 22924
rect 33152 22710 33180 22918
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 33244 22166 33272 23054
rect 33888 22574 33916 23598
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 33232 22160 33284 22166
rect 33232 22102 33284 22108
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 33980 22030 34008 27406
rect 35452 27402 35480 29650
rect 36096 29646 36124 29786
rect 35808 29640 35860 29646
rect 35808 29582 35860 29588
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 35716 29572 35768 29578
rect 35716 29514 35768 29520
rect 35728 29102 35756 29514
rect 35820 29102 35848 29582
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 36176 29504 36228 29510
rect 36176 29446 36228 29452
rect 35716 29096 35768 29102
rect 35716 29038 35768 29044
rect 35808 29096 35860 29102
rect 35808 29038 35860 29044
rect 35728 28694 35756 29038
rect 35716 28688 35768 28694
rect 35716 28630 35768 28636
rect 35820 28014 35848 29038
rect 36004 28762 36032 29446
rect 35992 28756 36044 28762
rect 35992 28698 36044 28704
rect 36188 28626 36216 29446
rect 36176 28620 36228 28626
rect 36176 28562 36228 28568
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 36268 28416 36320 28422
rect 36268 28358 36320 28364
rect 36096 28082 36124 28358
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 35808 28008 35860 28014
rect 35808 27950 35860 27956
rect 35440 27396 35492 27402
rect 35440 27338 35492 27344
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34808 25974 34836 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34888 26376 34940 26382
rect 34888 26318 34940 26324
rect 34796 25968 34848 25974
rect 34796 25910 34848 25916
rect 34520 25832 34572 25838
rect 34900 25786 34928 26318
rect 34520 25774 34572 25780
rect 34532 25498 34560 25774
rect 34808 25758 34928 25786
rect 34520 25492 34572 25498
rect 34520 25434 34572 25440
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 34072 24954 34100 25230
rect 34060 24948 34112 24954
rect 34060 24890 34112 24896
rect 34704 24812 34756 24818
rect 34704 24754 34756 24760
rect 34716 23730 34744 24754
rect 34808 23866 34836 25758
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 35452 25294 35480 27338
rect 35532 25696 35584 25702
rect 35532 25638 35584 25644
rect 35544 25362 35572 25638
rect 35532 25356 35584 25362
rect 35532 25298 35584 25304
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35820 25226 35848 27950
rect 35808 25220 35860 25226
rect 35808 25162 35860 25168
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 34796 23860 34848 23866
rect 34796 23802 34848 23808
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 34808 23186 34836 23802
rect 35452 23730 35480 24346
rect 35900 24132 35952 24138
rect 35900 24074 35952 24080
rect 35912 23866 35940 24074
rect 35900 23860 35952 23866
rect 35900 23802 35952 23808
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34796 23180 34848 23186
rect 34796 23122 34848 23128
rect 34704 23112 34756 23118
rect 34704 23054 34756 23060
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34624 22710 34652 22918
rect 34612 22704 34664 22710
rect 34612 22646 34664 22652
rect 34716 22098 34744 23054
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34704 22092 34756 22098
rect 34704 22034 34756 22040
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 33520 21554 33548 21830
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 33508 21548 33560 21554
rect 33508 21490 33560 21496
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32220 14340 32272 14346
rect 32220 14282 32272 14288
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 32140 1850 32168 3674
rect 32232 3398 32260 14282
rect 34808 12646 34836 22918
rect 35452 22642 35480 23666
rect 35716 23520 35768 23526
rect 35716 23462 35768 23468
rect 35728 23050 35756 23462
rect 35716 23044 35768 23050
rect 35716 22986 35768 22992
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 35348 22432 35400 22438
rect 35348 22374 35400 22380
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35360 22098 35388 22374
rect 35452 22098 35480 22578
rect 35348 22092 35400 22098
rect 35348 22034 35400 22040
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35624 21956 35676 21962
rect 35624 21898 35676 21904
rect 35636 21690 35664 21898
rect 35624 21684 35676 21690
rect 35624 21626 35676 21632
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 36004 16574 36032 28018
rect 36176 28008 36228 28014
rect 36176 27950 36228 27956
rect 36188 26518 36216 27950
rect 36280 27946 36308 28358
rect 36372 28014 36400 32302
rect 36452 29640 36504 29646
rect 36452 29582 36504 29588
rect 36464 28490 36492 29582
rect 36556 28626 36584 32914
rect 37476 32434 37504 32982
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37372 31748 37424 31754
rect 37372 31690 37424 31696
rect 37384 31482 37412 31690
rect 37372 31476 37424 31482
rect 37372 31418 37424 31424
rect 37096 31340 37148 31346
rect 37096 31282 37148 31288
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 36820 30728 36872 30734
rect 36820 30670 36872 30676
rect 36832 29714 36860 30670
rect 37004 30660 37056 30666
rect 37004 30602 37056 30608
rect 36820 29708 36872 29714
rect 36820 29650 36872 29656
rect 37016 29578 37044 30602
rect 37108 30598 37136 31282
rect 37096 30592 37148 30598
rect 37096 30534 37148 30540
rect 37108 30190 37136 30534
rect 37096 30184 37148 30190
rect 37096 30126 37148 30132
rect 37004 29572 37056 29578
rect 37004 29514 37056 29520
rect 37016 29458 37044 29514
rect 37016 29430 37136 29458
rect 36544 28620 36596 28626
rect 36544 28562 36596 28568
rect 36452 28484 36504 28490
rect 36452 28426 36504 28432
rect 36360 28008 36412 28014
rect 36360 27950 36412 27956
rect 36268 27940 36320 27946
rect 36268 27882 36320 27888
rect 36360 27872 36412 27878
rect 36360 27814 36412 27820
rect 36372 27674 36400 27814
rect 36360 27668 36412 27674
rect 36360 27610 36412 27616
rect 36464 27538 36492 28426
rect 36452 27532 36504 27538
rect 36452 27474 36504 27480
rect 36176 26512 36228 26518
rect 36176 26454 36228 26460
rect 36188 26042 36216 26454
rect 36176 26036 36228 26042
rect 36176 25978 36228 25984
rect 36084 25220 36136 25226
rect 36084 25162 36136 25168
rect 36096 24138 36124 25162
rect 36556 24426 36584 28562
rect 37108 25294 37136 29430
rect 37292 29034 37320 31282
rect 38488 30258 38516 45222
rect 38856 35894 38884 45526
rect 38856 35866 39160 35894
rect 37648 30252 37700 30258
rect 37648 30194 37700 30200
rect 38476 30252 38528 30258
rect 38476 30194 38528 30200
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37476 29170 37504 29990
rect 37660 29850 37688 30194
rect 38292 30184 38344 30190
rect 38292 30126 38344 30132
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 37648 29844 37700 29850
rect 37648 29786 37700 29792
rect 37660 29510 37688 29786
rect 37648 29504 37700 29510
rect 37648 29446 37700 29452
rect 37660 29170 37688 29446
rect 37844 29170 37872 30058
rect 38016 30048 38068 30054
rect 38016 29990 38068 29996
rect 37924 29572 37976 29578
rect 37924 29514 37976 29520
rect 37464 29164 37516 29170
rect 37464 29106 37516 29112
rect 37648 29164 37700 29170
rect 37648 29106 37700 29112
rect 37832 29164 37884 29170
rect 37832 29106 37884 29112
rect 37936 29034 37964 29514
rect 38028 29238 38056 29990
rect 38016 29232 38068 29238
rect 38016 29174 38068 29180
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 37740 29028 37792 29034
rect 37740 28970 37792 28976
rect 37924 29028 37976 29034
rect 37924 28970 37976 28976
rect 37752 28082 37780 28970
rect 38304 28626 38332 30126
rect 38476 29572 38528 29578
rect 38476 29514 38528 29520
rect 38488 29238 38516 29514
rect 38476 29232 38528 29238
rect 38476 29174 38528 29180
rect 38292 28620 38344 28626
rect 38292 28562 38344 28568
rect 37740 28076 37792 28082
rect 37740 28018 37792 28024
rect 37752 27470 37780 28018
rect 38016 27872 38068 27878
rect 38016 27814 38068 27820
rect 37740 27464 37792 27470
rect 37740 27406 37792 27412
rect 38028 27402 38056 27814
rect 38016 27396 38068 27402
rect 38016 27338 38068 27344
rect 38304 26994 38332 28562
rect 39028 28552 39080 28558
rect 39028 28494 39080 28500
rect 38384 27328 38436 27334
rect 38384 27270 38436 27276
rect 38292 26988 38344 26994
rect 38292 26930 38344 26936
rect 37740 26852 37792 26858
rect 37740 26794 37792 26800
rect 37752 25906 37780 26794
rect 37830 26480 37886 26489
rect 37830 26415 37832 26424
rect 37884 26415 37886 26424
rect 37832 26386 37884 26392
rect 37832 26308 37884 26314
rect 37832 26250 37884 26256
rect 37844 26042 37872 26250
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 37740 25900 37792 25906
rect 37740 25842 37792 25848
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 38200 25900 38252 25906
rect 38200 25842 38252 25848
rect 37464 25356 37516 25362
rect 37464 25298 37516 25304
rect 37096 25288 37148 25294
rect 37096 25230 37148 25236
rect 37004 24744 37056 24750
rect 37004 24686 37056 24692
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36464 24398 36584 24426
rect 36084 24132 36136 24138
rect 36084 24074 36136 24080
rect 36360 24132 36412 24138
rect 36360 24074 36412 24080
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 36188 23798 36216 24006
rect 36176 23792 36228 23798
rect 36176 23734 36228 23740
rect 36372 23730 36400 24074
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36372 23594 36400 23666
rect 36360 23588 36412 23594
rect 36360 23530 36412 23536
rect 36464 23322 36492 24398
rect 36740 24138 36768 24550
rect 37016 24206 37044 24686
rect 37108 24342 37136 25230
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 37292 24410 37320 24754
rect 37476 24614 37504 25298
rect 37752 25242 37780 25842
rect 37936 25498 37964 25842
rect 37924 25492 37976 25498
rect 37924 25434 37976 25440
rect 37568 25214 37780 25242
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 37464 24608 37516 24614
rect 37464 24550 37516 24556
rect 37280 24404 37332 24410
rect 37280 24346 37332 24352
rect 37096 24336 37148 24342
rect 37096 24278 37148 24284
rect 37004 24200 37056 24206
rect 37004 24142 37056 24148
rect 36728 24132 36780 24138
rect 36728 24074 36780 24080
rect 36544 24064 36596 24070
rect 36544 24006 36596 24012
rect 36556 23730 36584 24006
rect 36740 23730 36768 24074
rect 37568 23730 37596 25214
rect 38028 24886 38056 25230
rect 38016 24880 38068 24886
rect 38016 24822 38068 24828
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37752 24041 37780 24074
rect 37924 24064 37976 24070
rect 37738 24032 37794 24041
rect 37924 24006 37976 24012
rect 37738 23967 37794 23976
rect 37936 23730 37964 24006
rect 36544 23724 36596 23730
rect 36544 23666 36596 23672
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 37556 23724 37608 23730
rect 37556 23666 37608 23672
rect 37924 23724 37976 23730
rect 37924 23666 37976 23672
rect 37280 23656 37332 23662
rect 37280 23598 37332 23604
rect 36452 23316 36504 23322
rect 36452 23258 36504 23264
rect 36464 22710 36492 23258
rect 37292 23050 37320 23598
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 37464 23044 37516 23050
rect 37464 22986 37516 22992
rect 37476 22710 37504 22986
rect 36452 22704 36504 22710
rect 36452 22646 36504 22652
rect 37464 22704 37516 22710
rect 37464 22646 37516 22652
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37292 21554 37320 22578
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 36004 16546 36400 16574
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 12640 34848 12646
rect 34796 12582 34848 12588
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32784 3466 32812 3674
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 32772 3460 32824 3466
rect 32772 3402 32824 3408
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32692 2854 32720 3334
rect 32772 3188 32824 3194
rect 32772 3130 32824 3136
rect 32784 2854 32812 3130
rect 33060 3126 33088 3470
rect 33048 3120 33100 3126
rect 33048 3062 33100 3068
rect 33244 2990 33272 3470
rect 36280 3466 36308 4014
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 36268 3460 36320 3466
rect 36268 3402 36320 3408
rect 36188 3194 36216 3402
rect 36176 3188 36228 3194
rect 36176 3130 36228 3136
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 32680 2848 32732 2854
rect 32680 2790 32732 2796
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 32140 1822 32260 1850
rect 32232 800 32260 1822
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 800 35480 2382
rect 36096 800 36124 2994
rect 36372 2310 36400 16546
rect 38028 8362 38056 24822
rect 38212 24138 38240 25842
rect 38304 25702 38332 26930
rect 38396 26314 38424 27270
rect 38660 26784 38712 26790
rect 38660 26726 38712 26732
rect 38384 26308 38436 26314
rect 38384 26250 38436 26256
rect 38292 25696 38344 25702
rect 38292 25638 38344 25644
rect 38304 25362 38332 25638
rect 38292 25356 38344 25362
rect 38292 25298 38344 25304
rect 38304 24410 38332 25298
rect 38672 25158 38700 26726
rect 38752 26240 38804 26246
rect 38752 26182 38804 26188
rect 38764 25906 38792 26182
rect 38752 25900 38804 25906
rect 38752 25842 38804 25848
rect 38660 25152 38712 25158
rect 38660 25094 38712 25100
rect 38764 24750 38792 25842
rect 38752 24744 38804 24750
rect 38752 24686 38804 24692
rect 38292 24404 38344 24410
rect 38292 24346 38344 24352
rect 38568 24200 38620 24206
rect 38568 24142 38620 24148
rect 38200 24132 38252 24138
rect 38200 24074 38252 24080
rect 38580 23730 38608 24142
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38580 23322 38608 23666
rect 38568 23316 38620 23322
rect 38568 23258 38620 23264
rect 38200 22432 38252 22438
rect 38200 22374 38252 22380
rect 38212 22234 38240 22374
rect 38200 22228 38252 22234
rect 38200 22170 38252 22176
rect 38936 21888 38988 21894
rect 38936 21830 38988 21836
rect 38948 21622 38976 21830
rect 38936 21616 38988 21622
rect 38936 21558 38988 21564
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 38016 3596 38068 3602
rect 38016 3538 38068 3544
rect 38028 3482 38056 3538
rect 37844 3466 38056 3482
rect 37832 3460 38056 3466
rect 37884 3454 38056 3460
rect 37832 3402 37884 3408
rect 38396 2961 38424 3878
rect 38488 3534 38516 3878
rect 38476 3528 38528 3534
rect 38476 3470 38528 3476
rect 38476 3392 38528 3398
rect 38580 3346 38608 4082
rect 38934 3768 38990 3777
rect 38934 3703 38936 3712
rect 38988 3703 38990 3712
rect 38936 3674 38988 3680
rect 38528 3340 38608 3346
rect 38476 3334 38608 3340
rect 38488 3318 38608 3334
rect 38488 3058 38516 3318
rect 38476 3052 38528 3058
rect 38476 2994 38528 3000
rect 38382 2952 38438 2961
rect 38382 2887 38438 2896
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 38028 800 38056 2314
rect 39040 2310 39068 28494
rect 39132 21486 39160 35866
rect 40052 32842 40080 47398
rect 40408 46980 40460 46986
rect 40408 46922 40460 46928
rect 40040 32836 40092 32842
rect 40040 32778 40092 32784
rect 40224 26444 40276 26450
rect 40224 26386 40276 26392
rect 40236 25906 40264 26386
rect 40420 25974 40448 46922
rect 41236 46368 41288 46374
rect 41236 46310 41288 46316
rect 41248 46034 41276 46310
rect 41892 46034 41920 49200
rect 42536 46442 42564 49200
rect 43180 47122 43208 49200
rect 43168 47116 43220 47122
rect 43168 47058 43220 47064
rect 42616 47048 42668 47054
rect 42616 46990 42668 46996
rect 42628 46594 42656 46990
rect 43168 46980 43220 46986
rect 43168 46922 43220 46928
rect 42628 46566 42748 46594
rect 42616 46504 42668 46510
rect 42616 46446 42668 46452
rect 42524 46436 42576 46442
rect 42524 46378 42576 46384
rect 41236 46028 41288 46034
rect 41236 45970 41288 45976
rect 41880 46028 41932 46034
rect 41880 45970 41932 45976
rect 41420 45892 41472 45898
rect 41420 45834 41472 45840
rect 40776 45824 40828 45830
rect 40776 45766 40828 45772
rect 40408 25968 40460 25974
rect 40408 25910 40460 25916
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 40236 25294 40264 25842
rect 40788 25362 40816 45766
rect 41432 45626 41460 45834
rect 42628 45626 42656 46446
rect 41420 45620 41472 45626
rect 41420 45562 41472 45568
rect 42616 45620 42668 45626
rect 42616 45562 42668 45568
rect 41052 45484 41104 45490
rect 41052 45426 41104 45432
rect 41064 44266 41092 45426
rect 42720 45082 42748 46566
rect 43180 45558 43208 46922
rect 43824 45966 43852 49200
rect 44468 47410 44496 49200
rect 44192 47382 44496 47410
rect 43812 45960 43864 45966
rect 43812 45902 43864 45908
rect 44192 45558 44220 47382
rect 44456 47048 44508 47054
rect 44456 46990 44508 46996
rect 44272 45892 44324 45898
rect 44272 45834 44324 45840
rect 43168 45552 43220 45558
rect 43168 45494 43220 45500
rect 44180 45552 44232 45558
rect 44180 45494 44232 45500
rect 42708 45076 42760 45082
rect 42708 45018 42760 45024
rect 41052 44260 41104 44266
rect 41052 44202 41104 44208
rect 41064 25974 41092 44202
rect 42800 41064 42852 41070
rect 42800 41006 42852 41012
rect 42812 39914 42840 41006
rect 42800 39908 42852 39914
rect 42800 39850 42852 39856
rect 42064 38956 42116 38962
rect 42064 38898 42116 38904
rect 42076 27606 42104 38898
rect 41420 27600 41472 27606
rect 41420 27542 41472 27548
rect 42064 27600 42116 27606
rect 42064 27542 42116 27548
rect 41432 26382 41460 27542
rect 44284 26994 44312 45834
rect 44468 45082 44496 46990
rect 45008 46096 45060 46102
rect 45008 46038 45060 46044
rect 44548 45416 44600 45422
rect 44548 45358 44600 45364
rect 44456 45076 44508 45082
rect 44456 45018 44508 45024
rect 44560 44402 44588 45358
rect 45020 44878 45048 46038
rect 45112 45626 45140 49200
rect 45376 46980 45428 46986
rect 45376 46922 45428 46928
rect 45100 45620 45152 45626
rect 45100 45562 45152 45568
rect 45100 45416 45152 45422
rect 45100 45358 45152 45364
rect 45112 45082 45140 45358
rect 45388 45082 45416 46922
rect 45756 45966 45784 49200
rect 45744 45960 45796 45966
rect 45744 45902 45796 45908
rect 45836 45960 45888 45966
rect 45836 45902 45888 45908
rect 45652 45824 45704 45830
rect 45652 45766 45704 45772
rect 45560 45620 45612 45626
rect 45560 45562 45612 45568
rect 45572 45422 45600 45562
rect 45560 45416 45612 45422
rect 45560 45358 45612 45364
rect 45100 45076 45152 45082
rect 45100 45018 45152 45024
rect 45376 45076 45428 45082
rect 45376 45018 45428 45024
rect 45008 44872 45060 44878
rect 45008 44814 45060 44820
rect 45560 44872 45612 44878
rect 45560 44814 45612 44820
rect 44548 44396 44600 44402
rect 44548 44338 44600 44344
rect 45100 40520 45152 40526
rect 45100 40462 45152 40468
rect 44272 26988 44324 26994
rect 44272 26930 44324 26936
rect 41420 26376 41472 26382
rect 41420 26318 41472 26324
rect 41052 25968 41104 25974
rect 41052 25910 41104 25916
rect 41144 25968 41196 25974
rect 41144 25910 41196 25916
rect 40316 25356 40368 25362
rect 40316 25298 40368 25304
rect 40776 25356 40828 25362
rect 40776 25298 40828 25304
rect 40224 25288 40276 25294
rect 40224 25230 40276 25236
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 40224 18420 40276 18426
rect 40224 18362 40276 18368
rect 40236 17746 40264 18362
rect 40224 17740 40276 17746
rect 40224 17682 40276 17688
rect 40040 16516 40092 16522
rect 40040 16458 40092 16464
rect 40052 16114 40080 16458
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 40328 15502 40356 25298
rect 40684 20052 40736 20058
rect 40684 19994 40736 20000
rect 40696 19446 40724 19994
rect 40684 19440 40736 19446
rect 40684 19382 40736 19388
rect 40408 17604 40460 17610
rect 40408 17546 40460 17552
rect 40316 15496 40368 15502
rect 40316 15438 40368 15444
rect 40420 12434 40448 17546
rect 40500 16040 40552 16046
rect 40500 15982 40552 15988
rect 40512 15706 40540 15982
rect 40500 15700 40552 15706
rect 40500 15642 40552 15648
rect 41064 14074 41092 25910
rect 41156 25430 41184 25910
rect 41144 25424 41196 25430
rect 41144 25366 41196 25372
rect 41432 23118 41460 26318
rect 43996 26308 44048 26314
rect 43996 26250 44048 26256
rect 41420 23112 41472 23118
rect 41420 23054 41472 23060
rect 41328 23044 41380 23050
rect 41328 22986 41380 22992
rect 41340 22438 41368 22986
rect 41432 22710 41460 23054
rect 41604 22976 41656 22982
rect 41604 22918 41656 22924
rect 41420 22704 41472 22710
rect 41420 22646 41472 22652
rect 41328 22432 41380 22438
rect 41328 22374 41380 22380
rect 41616 22030 41644 22918
rect 44008 22574 44036 26250
rect 44088 23656 44140 23662
rect 44088 23598 44140 23604
rect 42432 22568 42484 22574
rect 42432 22510 42484 22516
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 43996 22568 44048 22574
rect 43996 22510 44048 22516
rect 41604 22024 41656 22030
rect 41604 21966 41656 21972
rect 42444 21078 42472 22510
rect 42628 22234 42656 22510
rect 42616 22228 42668 22234
rect 42616 22170 42668 22176
rect 42708 22092 42760 22098
rect 42708 22034 42760 22040
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42628 21554 42656 21966
rect 42720 21622 42748 22034
rect 42800 21956 42852 21962
rect 42800 21898 42852 21904
rect 42708 21616 42760 21622
rect 42708 21558 42760 21564
rect 42616 21548 42668 21554
rect 42616 21490 42668 21496
rect 42432 21072 42484 21078
rect 42432 21014 42484 21020
rect 42524 21004 42576 21010
rect 42524 20946 42576 20952
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 41420 19168 41472 19174
rect 41420 19110 41472 19116
rect 41340 18902 41368 19110
rect 41328 18896 41380 18902
rect 41328 18838 41380 18844
rect 41432 18834 41460 19110
rect 41420 18828 41472 18834
rect 41420 18770 41472 18776
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41052 14068 41104 14074
rect 41052 14010 41104 14016
rect 40420 12406 40540 12434
rect 39488 4276 39540 4282
rect 39488 4218 39540 4224
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 39224 3738 39252 4082
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 39212 3732 39264 3738
rect 39212 3674 39264 3680
rect 39408 3670 39436 4014
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 39500 3534 39528 4218
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39488 3528 39540 3534
rect 39488 3470 39540 3476
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39500 3058 39528 3334
rect 39488 3052 39540 3058
rect 39488 2994 39540 3000
rect 39776 2774 39804 3538
rect 39868 3194 39896 4082
rect 40040 4004 40092 4010
rect 40040 3946 40092 3952
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 39960 3194 39988 3470
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39948 3188 40000 3194
rect 39948 3130 40000 3136
rect 40052 2854 40080 3946
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 40328 3126 40356 3470
rect 40316 3120 40368 3126
rect 40316 3062 40368 3068
rect 40130 2952 40186 2961
rect 40130 2887 40186 2896
rect 40144 2854 40172 2887
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 39684 2746 39804 2774
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 39028 2304 39080 2310
rect 39028 2246 39080 2252
rect 39316 800 39344 2314
rect 39684 1850 39712 2746
rect 40512 2582 40540 12406
rect 41064 10674 41092 14010
rect 41052 10668 41104 10674
rect 41052 10610 41104 10616
rect 41248 5778 41276 18702
rect 41880 16040 41932 16046
rect 41880 15982 41932 15988
rect 41892 8294 41920 15982
rect 42536 12434 42564 20946
rect 42628 20942 42656 21490
rect 42616 20936 42668 20942
rect 42616 20878 42668 20884
rect 42628 20534 42656 20878
rect 42616 20528 42668 20534
rect 42616 20470 42668 20476
rect 42352 12406 42564 12434
rect 41880 8288 41932 8294
rect 41880 8230 41932 8236
rect 41236 5772 41288 5778
rect 41236 5714 41288 5720
rect 41236 4208 41288 4214
rect 41236 4150 41288 4156
rect 41052 4140 41104 4146
rect 41052 4082 41104 4088
rect 41064 3942 41092 4082
rect 41144 4072 41196 4078
rect 41144 4014 41196 4020
rect 41052 3936 41104 3942
rect 41052 3878 41104 3884
rect 41156 3466 41184 4014
rect 41248 3777 41276 4150
rect 41420 4140 41472 4146
rect 41420 4082 41472 4088
rect 41432 3942 41460 4082
rect 41328 3936 41380 3942
rect 41328 3878 41380 3884
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41234 3768 41290 3777
rect 41234 3703 41290 3712
rect 41340 3602 41368 3878
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 41144 3460 41196 3466
rect 41144 3402 41196 3408
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 40500 2576 40552 2582
rect 40500 2518 40552 2524
rect 41340 2514 41368 3402
rect 42352 3398 42380 12406
rect 42720 9586 42748 21558
rect 42812 21486 42840 21898
rect 44100 21690 44128 23598
rect 44088 21684 44140 21690
rect 44088 21626 44140 21632
rect 42800 21480 42852 21486
rect 42800 21422 42852 21428
rect 43260 21412 43312 21418
rect 43260 21354 43312 21360
rect 43168 20528 43220 20534
rect 43168 20470 43220 20476
rect 43180 20262 43208 20470
rect 43168 20256 43220 20262
rect 43168 20198 43220 20204
rect 43180 19378 43208 20198
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 43272 5234 43300 21354
rect 43904 19372 43956 19378
rect 43904 19314 43956 19320
rect 43916 15502 43944 19314
rect 45112 16574 45140 40462
rect 45572 38418 45600 44814
rect 45560 38412 45612 38418
rect 45560 38354 45612 38360
rect 45560 31204 45612 31210
rect 45560 31146 45612 31152
rect 45192 26376 45244 26382
rect 45192 26318 45244 26324
rect 45204 23730 45232 26318
rect 45572 25906 45600 31146
rect 45664 25974 45692 45766
rect 45848 45554 45876 45902
rect 46400 45626 46428 49200
rect 46846 47696 46902 47705
rect 46846 47631 46902 47640
rect 46754 47016 46810 47025
rect 46754 46951 46810 46960
rect 46664 46504 46716 46510
rect 46664 46446 46716 46452
rect 46480 45892 46532 45898
rect 46480 45834 46532 45840
rect 46388 45620 46440 45626
rect 46388 45562 46440 45568
rect 45756 45526 45876 45554
rect 45756 44402 45784 45526
rect 46388 45348 46440 45354
rect 46388 45290 46440 45296
rect 46204 44872 46256 44878
rect 46204 44814 46256 44820
rect 45744 44396 45796 44402
rect 45744 44338 45796 44344
rect 46112 40384 46164 40390
rect 46112 40326 46164 40332
rect 45928 40112 45980 40118
rect 45928 40054 45980 40060
rect 45836 38956 45888 38962
rect 45836 38898 45888 38904
rect 45848 38350 45876 38898
rect 45836 38344 45888 38350
rect 45836 38286 45888 38292
rect 45848 37874 45876 38286
rect 45836 37868 45888 37874
rect 45836 37810 45888 37816
rect 45848 37262 45876 37810
rect 45836 37256 45888 37262
rect 45836 37198 45888 37204
rect 45848 36786 45876 37198
rect 45836 36780 45888 36786
rect 45836 36722 45888 36728
rect 45836 34128 45888 34134
rect 45836 34070 45888 34076
rect 45652 25968 45704 25974
rect 45652 25910 45704 25916
rect 45560 25900 45612 25906
rect 45560 25842 45612 25848
rect 45572 24970 45600 25842
rect 45744 25356 45796 25362
rect 45744 25298 45796 25304
rect 45652 25152 45704 25158
rect 45652 25094 45704 25100
rect 45480 24942 45600 24970
rect 45192 23724 45244 23730
rect 45192 23666 45244 23672
rect 45480 23338 45508 24942
rect 45480 23310 45600 23338
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45480 21146 45508 21966
rect 45468 21140 45520 21146
rect 45468 21082 45520 21088
rect 45468 20460 45520 20466
rect 45468 20402 45520 20408
rect 45480 19990 45508 20402
rect 45572 20058 45600 23310
rect 45664 22574 45692 25094
rect 45652 22568 45704 22574
rect 45652 22510 45704 22516
rect 45652 21956 45704 21962
rect 45652 21898 45704 21904
rect 45664 21690 45692 21898
rect 45652 21684 45704 21690
rect 45652 21626 45704 21632
rect 45756 21554 45784 25298
rect 45744 21548 45796 21554
rect 45744 21490 45796 21496
rect 45744 20392 45796 20398
rect 45744 20334 45796 20340
rect 45560 20052 45612 20058
rect 45560 19994 45612 20000
rect 45468 19984 45520 19990
rect 45468 19926 45520 19932
rect 45480 19514 45508 19926
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45468 19508 45520 19514
rect 45468 19450 45520 19456
rect 45572 19446 45600 19790
rect 45560 19440 45612 19446
rect 45560 19382 45612 19388
rect 45572 18766 45600 19382
rect 45756 19378 45784 20334
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 45560 18760 45612 18766
rect 45560 18702 45612 18708
rect 45756 18714 45784 19314
rect 45848 18834 45876 34070
rect 45940 20602 45968 40054
rect 46124 40050 46152 40326
rect 46112 40044 46164 40050
rect 46112 39986 46164 39992
rect 46110 39536 46166 39545
rect 46110 39471 46166 39480
rect 46020 38412 46072 38418
rect 46020 38354 46072 38360
rect 46032 31210 46060 38354
rect 46020 31204 46072 31210
rect 46020 31146 46072 31152
rect 46124 31090 46152 39471
rect 46216 37806 46244 44814
rect 46296 42696 46348 42702
rect 46296 42638 46348 42644
rect 46308 42226 46336 42638
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46400 41138 46428 45290
rect 46492 44538 46520 45834
rect 46676 45558 46704 46446
rect 46664 45552 46716 45558
rect 46664 45494 46716 45500
rect 46480 44532 46532 44538
rect 46480 44474 46532 44480
rect 46572 44396 46624 44402
rect 46572 44338 46624 44344
rect 46664 44396 46716 44402
rect 46664 44338 46716 44344
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46388 41132 46440 41138
rect 46388 41074 46440 41080
rect 46296 38344 46348 38350
rect 46296 38286 46348 38292
rect 46204 37800 46256 37806
rect 46204 37742 46256 37748
rect 46216 36174 46244 37742
rect 46308 37466 46336 38286
rect 46296 37460 46348 37466
rect 46296 37402 46348 37408
rect 46400 36854 46428 41074
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46492 39506 46520 39782
rect 46480 39500 46532 39506
rect 46480 39442 46532 39448
rect 46584 37194 46612 44338
rect 46676 38894 46704 44338
rect 46664 38888 46716 38894
rect 46664 38830 46716 38836
rect 46572 37188 46624 37194
rect 46572 37130 46624 37136
rect 46388 36848 46440 36854
rect 46388 36790 46440 36796
rect 46204 36168 46256 36174
rect 46204 36110 46256 36116
rect 46296 32904 46348 32910
rect 46296 32846 46348 32852
rect 46308 32026 46336 32846
rect 46296 32020 46348 32026
rect 46296 31962 46348 31968
rect 46202 31376 46258 31385
rect 46202 31311 46258 31320
rect 46032 31062 46152 31090
rect 46032 24970 46060 31062
rect 46112 28688 46164 28694
rect 46112 28630 46164 28636
rect 46124 25158 46152 28630
rect 46216 25945 46244 31311
rect 46296 28552 46348 28558
rect 46296 28494 46348 28500
rect 46202 25936 46258 25945
rect 46202 25871 46258 25880
rect 46308 25294 46336 28494
rect 46296 25288 46348 25294
rect 46296 25230 46348 25236
rect 46112 25152 46164 25158
rect 46112 25094 46164 25100
rect 46032 24942 46152 24970
rect 46020 24812 46072 24818
rect 46020 24754 46072 24760
rect 46032 22710 46060 24754
rect 46020 22704 46072 22710
rect 46020 22646 46072 22652
rect 46124 21978 46152 24942
rect 46204 24744 46256 24750
rect 46204 24686 46256 24692
rect 46216 23225 46244 24686
rect 46202 23216 46258 23225
rect 46308 23202 46336 25230
rect 46400 23338 46428 36790
rect 46584 28082 46612 37130
rect 46676 32502 46704 38830
rect 46664 32496 46716 32502
rect 46664 32438 46716 32444
rect 46572 28076 46624 28082
rect 46572 28018 46624 28024
rect 46768 26234 46796 46951
rect 46860 46510 46888 47631
rect 46848 46504 46900 46510
rect 46848 46446 46900 46452
rect 47044 46034 47072 49200
rect 47688 47054 47716 49200
rect 48332 47122 48360 49200
rect 48320 47116 48372 47122
rect 48320 47058 48372 47064
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 47952 46912 48004 46918
rect 47952 46854 48004 46860
rect 47860 46572 47912 46578
rect 47860 46514 47912 46520
rect 47768 46436 47820 46442
rect 47768 46378 47820 46384
rect 47032 46028 47084 46034
rect 47032 45970 47084 45976
rect 46848 45824 46900 45830
rect 46848 45766 46900 45772
rect 46860 45490 46888 45766
rect 46848 45484 46900 45490
rect 46848 45426 46900 45432
rect 47124 45416 47176 45422
rect 47124 45358 47176 45364
rect 47032 44940 47084 44946
rect 47032 44882 47084 44888
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 46952 43858 46980 44134
rect 46940 43852 46992 43858
rect 46940 43794 46992 43800
rect 47044 43314 47072 44882
rect 47032 43308 47084 43314
rect 47032 43250 47084 43256
rect 47136 42158 47164 45358
rect 47308 45280 47360 45286
rect 47308 45222 47360 45228
rect 46940 42152 46992 42158
rect 46940 42094 46992 42100
rect 47124 42152 47176 42158
rect 47124 42094 47176 42100
rect 46846 40896 46902 40905
rect 46846 40831 46902 40840
rect 46860 40526 46888 40831
rect 46848 40520 46900 40526
rect 46848 40462 46900 40468
rect 46848 32428 46900 32434
rect 46848 32370 46900 32376
rect 46860 32065 46888 32370
rect 46846 32056 46902 32065
rect 46846 31991 46902 32000
rect 46952 31090 46980 42094
rect 47124 34944 47176 34950
rect 47124 34886 47176 34892
rect 47136 34066 47164 34886
rect 47216 34400 47268 34406
rect 47216 34342 47268 34348
rect 47124 34060 47176 34066
rect 47124 34002 47176 34008
rect 47228 33930 47256 34342
rect 47216 33924 47268 33930
rect 47216 33866 47268 33872
rect 47216 32428 47268 32434
rect 47216 32370 47268 32376
rect 46952 31062 47164 31090
rect 46846 30016 46902 30025
rect 46846 29951 46902 29960
rect 46860 29306 46888 29951
rect 46940 29708 46992 29714
rect 46940 29650 46992 29656
rect 46848 29300 46900 29306
rect 46848 29242 46900 29248
rect 46952 28626 46980 29650
rect 46940 28620 46992 28626
rect 46940 28562 46992 28568
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47044 27538 47072 27814
rect 47032 27532 47084 27538
rect 47032 27474 47084 27480
rect 46846 26616 46902 26625
rect 46846 26551 46902 26560
rect 46860 26314 46888 26551
rect 46848 26308 46900 26314
rect 46848 26250 46900 26256
rect 46676 26206 46796 26234
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 46480 24608 46532 24614
rect 46480 24550 46532 24556
rect 46492 24274 46520 24550
rect 46480 24268 46532 24274
rect 46480 24210 46532 24216
rect 46572 23656 46624 23662
rect 46572 23598 46624 23604
rect 46400 23310 46520 23338
rect 46308 23174 46428 23202
rect 46202 23151 46258 23160
rect 46296 23112 46348 23118
rect 46296 23054 46348 23060
rect 46202 22536 46258 22545
rect 46202 22471 46258 22480
rect 46032 21950 46152 21978
rect 46032 20618 46060 21950
rect 46110 21856 46166 21865
rect 46110 21791 46166 21800
rect 46124 21486 46152 21791
rect 46216 21554 46244 22471
rect 46308 22234 46336 23054
rect 46296 22228 46348 22234
rect 46296 22170 46348 22176
rect 46400 22114 46428 23174
rect 46308 22086 46428 22114
rect 46204 21548 46256 21554
rect 46204 21490 46256 21496
rect 46112 21480 46164 21486
rect 46112 21422 46164 21428
rect 45928 20596 45980 20602
rect 46032 20590 46152 20618
rect 45928 20538 45980 20544
rect 46020 20460 46072 20466
rect 46020 20402 46072 20408
rect 45928 19780 45980 19786
rect 45928 19722 45980 19728
rect 45940 19514 45968 19722
rect 45928 19508 45980 19514
rect 45928 19450 45980 19456
rect 45836 18828 45888 18834
rect 45836 18770 45888 18776
rect 45940 18766 45968 19450
rect 46032 18970 46060 20402
rect 46124 19990 46152 20590
rect 46112 19984 46164 19990
rect 46112 19926 46164 19932
rect 46204 19848 46256 19854
rect 46204 19790 46256 19796
rect 46112 19712 46164 19718
rect 46112 19654 46164 19660
rect 46124 19378 46152 19654
rect 46112 19372 46164 19378
rect 46112 19314 46164 19320
rect 46216 19310 46244 19790
rect 46204 19304 46256 19310
rect 46124 19252 46204 19258
rect 46124 19246 46256 19252
rect 46124 19230 46244 19246
rect 46020 18964 46072 18970
rect 46020 18906 46072 18912
rect 46020 18828 46072 18834
rect 46020 18770 46072 18776
rect 45928 18760 45980 18766
rect 45468 17672 45520 17678
rect 45468 17614 45520 17620
rect 45480 17270 45508 17614
rect 45468 17264 45520 17270
rect 45468 17206 45520 17212
rect 45020 16546 45140 16574
rect 44088 16040 44140 16046
rect 44088 15982 44140 15988
rect 44100 15706 44128 15982
rect 44088 15700 44140 15706
rect 44088 15642 44140 15648
rect 43536 15496 43588 15502
rect 43536 15438 43588 15444
rect 43904 15496 43956 15502
rect 43904 15438 43956 15444
rect 43548 14414 43576 15438
rect 43720 14952 43772 14958
rect 43720 14894 43772 14900
rect 43732 14618 43760 14894
rect 43720 14612 43772 14618
rect 43720 14554 43772 14560
rect 43536 14408 43588 14414
rect 43536 14350 43588 14356
rect 43548 13870 43576 14350
rect 43536 13864 43588 13870
rect 43536 13806 43588 13812
rect 43260 5228 43312 5234
rect 43260 5170 43312 5176
rect 42432 4616 42484 4622
rect 42432 4558 42484 4564
rect 42340 3392 42392 3398
rect 42340 3334 42392 3340
rect 42444 3058 42472 4558
rect 43076 4480 43128 4486
rect 43076 4422 43128 4428
rect 43088 4214 43116 4422
rect 43076 4208 43128 4214
rect 43076 4150 43128 4156
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 39684 1822 39988 1850
rect 39960 800 39988 1822
rect 40604 800 40632 2314
rect 41248 800 41276 2382
rect 42536 800 42564 3606
rect 42984 3460 43036 3466
rect 42984 3402 43036 3408
rect 42616 3392 42668 3398
rect 42616 3334 42668 3340
rect 42628 3126 42656 3334
rect 42616 3120 42668 3126
rect 42616 3062 42668 3068
rect 42996 2990 43024 3402
rect 42984 2984 43036 2990
rect 42984 2926 43036 2932
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 43180 800 43208 2926
rect 43272 2922 43300 5170
rect 43812 4616 43864 4622
rect 43812 4558 43864 4564
rect 43260 2916 43312 2922
rect 43260 2858 43312 2864
rect 43824 800 43852 4558
rect 45020 4146 45048 16546
rect 45480 16182 45508 17206
rect 45572 16574 45600 18702
rect 45756 18686 45876 18714
rect 45928 18702 45980 18708
rect 45744 17196 45796 17202
rect 45744 17138 45796 17144
rect 45572 16546 45692 16574
rect 45468 16176 45520 16182
rect 45468 16118 45520 16124
rect 45468 16040 45520 16046
rect 45468 15982 45520 15988
rect 45100 14952 45152 14958
rect 45100 14894 45152 14900
rect 45008 4140 45060 4146
rect 45008 4082 45060 4088
rect 45112 800 45140 14894
rect 45376 9512 45428 9518
rect 45376 9454 45428 9460
rect 45192 4616 45244 4622
rect 45192 4558 45244 4564
rect 45204 3058 45232 4558
rect 45388 3534 45416 9454
rect 45480 3942 45508 15982
rect 45560 12640 45612 12646
rect 45560 12582 45612 12588
rect 45572 12238 45600 12582
rect 45560 12232 45612 12238
rect 45560 12174 45612 12180
rect 45560 8288 45612 8294
rect 45558 8256 45560 8265
rect 45612 8256 45614 8265
rect 45558 8191 45614 8200
rect 45664 5370 45692 16546
rect 45756 15706 45784 17138
rect 45744 15700 45796 15706
rect 45744 15642 45796 15648
rect 45848 13954 45876 18686
rect 46032 16574 46060 18770
rect 45756 13938 45876 13954
rect 45744 13932 45876 13938
rect 45796 13926 45876 13932
rect 45940 16546 46060 16574
rect 45744 13874 45796 13880
rect 45836 13864 45888 13870
rect 45836 13806 45888 13812
rect 45848 12918 45876 13806
rect 45836 12912 45888 12918
rect 45836 12854 45888 12860
rect 45836 12776 45888 12782
rect 45940 12730 45968 16546
rect 46124 14362 46152 19230
rect 46216 19181 46244 19230
rect 46204 17128 46256 17134
rect 46204 17070 46256 17076
rect 46216 16046 46244 17070
rect 46204 16040 46256 16046
rect 46204 15982 46256 15988
rect 46308 15434 46336 22086
rect 46492 21434 46520 23310
rect 46584 22778 46612 23598
rect 46572 22772 46624 22778
rect 46572 22714 46624 22720
rect 46676 22098 46704 26206
rect 46846 25256 46902 25265
rect 46846 25191 46902 25200
rect 46756 24676 46808 24682
rect 46756 24618 46808 24624
rect 46768 23905 46796 24618
rect 46754 23896 46810 23905
rect 46754 23831 46810 23840
rect 46860 23662 46888 25191
rect 47136 24818 47164 31062
rect 47124 24812 47176 24818
rect 47124 24754 47176 24760
rect 46848 23656 46900 23662
rect 46848 23598 46900 23604
rect 47136 23050 47164 24754
rect 47124 23044 47176 23050
rect 47124 22986 47176 22992
rect 46664 22092 46716 22098
rect 46664 22034 46716 22040
rect 46664 21480 46716 21486
rect 46492 21406 46612 21434
rect 46664 21422 46716 21428
rect 46480 21344 46532 21350
rect 46480 21286 46532 21292
rect 46492 21010 46520 21286
rect 46480 21004 46532 21010
rect 46480 20946 46532 20952
rect 46480 20256 46532 20262
rect 46480 20198 46532 20204
rect 46492 19922 46520 20198
rect 46480 19916 46532 19922
rect 46480 19858 46532 19864
rect 46386 18456 46442 18465
rect 46386 18391 46442 18400
rect 46400 18290 46428 18391
rect 46388 18284 46440 18290
rect 46388 18226 46440 18232
rect 46584 16794 46612 21406
rect 46676 17814 46704 21422
rect 47136 18290 47164 22986
rect 47124 18284 47176 18290
rect 47124 18226 47176 18232
rect 46848 18080 46900 18086
rect 46848 18022 46900 18028
rect 47032 18080 47084 18086
rect 47032 18022 47084 18028
rect 46664 17808 46716 17814
rect 46664 17750 46716 17756
rect 46572 16788 46624 16794
rect 46572 16730 46624 16736
rect 46388 16176 46440 16182
rect 46388 16118 46440 16124
rect 46400 15570 46428 16118
rect 46860 16028 46888 18022
rect 47044 16658 47072 18022
rect 47032 16652 47084 16658
rect 47032 16594 47084 16600
rect 47124 16108 47176 16114
rect 47124 16050 47176 16056
rect 46940 16040 46992 16046
rect 46860 16000 46940 16028
rect 46940 15982 46992 15988
rect 46664 15972 46716 15978
rect 46664 15914 46716 15920
rect 46388 15564 46440 15570
rect 46388 15506 46440 15512
rect 46676 15502 46704 15914
rect 46848 15904 46900 15910
rect 46848 15846 46900 15852
rect 46860 15745 46888 15846
rect 46846 15736 46902 15745
rect 47136 15706 47164 16050
rect 46846 15671 46902 15680
rect 47124 15700 47176 15706
rect 47124 15642 47176 15648
rect 46664 15496 46716 15502
rect 46664 15438 46716 15444
rect 47032 15496 47084 15502
rect 47032 15438 47084 15444
rect 46296 15428 46348 15434
rect 46296 15370 46348 15376
rect 46388 15020 46440 15026
rect 46388 14962 46440 14968
rect 46124 14334 46244 14362
rect 46400 14346 46428 14962
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 14414 46520 14758
rect 46676 14414 46704 15438
rect 47044 15162 47072 15438
rect 47032 15156 47084 15162
rect 47032 15098 47084 15104
rect 46756 15020 46808 15026
rect 46756 14962 46808 14968
rect 46768 14482 46796 14962
rect 46848 14952 46900 14958
rect 46848 14894 46900 14900
rect 46756 14476 46808 14482
rect 46756 14418 46808 14424
rect 46480 14408 46532 14414
rect 46480 14350 46532 14356
rect 46664 14408 46716 14414
rect 46664 14350 46716 14356
rect 46112 14272 46164 14278
rect 46112 14214 46164 14220
rect 46124 13938 46152 14214
rect 46020 13932 46072 13938
rect 46020 13874 46072 13880
rect 46112 13932 46164 13938
rect 46112 13874 46164 13880
rect 45888 12724 45968 12730
rect 45836 12718 45968 12724
rect 45744 12708 45796 12714
rect 45848 12702 45968 12718
rect 45744 12650 45796 12656
rect 45756 12238 45784 12650
rect 46032 12442 46060 13874
rect 46124 13326 46152 13874
rect 46112 13320 46164 13326
rect 46112 13262 46164 13268
rect 46020 12436 46072 12442
rect 46020 12378 46072 12384
rect 45744 12232 45796 12238
rect 45744 12174 45796 12180
rect 45652 5364 45704 5370
rect 45652 5306 45704 5312
rect 45664 4282 45692 5306
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 45468 3936 45520 3942
rect 45468 3878 45520 3884
rect 45560 3936 45612 3942
rect 45560 3878 45612 3884
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45376 3528 45428 3534
rect 45376 3470 45428 3476
rect 45480 3398 45508 3538
rect 45572 3466 45600 3878
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 45664 3534 45692 3606
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 45560 3460 45612 3466
rect 45560 3402 45612 3408
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45388 3126 45416 3334
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45756 2582 45784 12174
rect 46112 11824 46164 11830
rect 46112 11766 46164 11772
rect 46020 11688 46072 11694
rect 46020 11630 46072 11636
rect 46032 5302 46060 11630
rect 46124 9450 46152 11766
rect 46112 9444 46164 9450
rect 46112 9386 46164 9392
rect 46216 7954 46244 14334
rect 46388 14340 46440 14346
rect 46388 14282 46440 14288
rect 46400 13938 46428 14282
rect 46768 14074 46796 14418
rect 46860 14414 46888 14894
rect 46848 14408 46900 14414
rect 46848 14350 46900 14356
rect 46756 14068 46808 14074
rect 46756 14010 46808 14016
rect 46860 13954 46888 14350
rect 46768 13938 46888 13954
rect 46388 13932 46440 13938
rect 46388 13874 46440 13880
rect 46756 13932 46888 13938
rect 46808 13926 46888 13932
rect 46756 13874 46808 13880
rect 46296 12164 46348 12170
rect 46296 12106 46348 12112
rect 46308 11694 46336 12106
rect 46296 11688 46348 11694
rect 46296 11630 46348 11636
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46204 7948 46256 7954
rect 46204 7890 46256 7896
rect 46204 6248 46256 6254
rect 46202 6216 46204 6225
rect 46256 6216 46258 6225
rect 46202 6151 46258 6160
rect 46204 5636 46256 5642
rect 46204 5578 46256 5584
rect 46020 5296 46072 5302
rect 46020 5238 46072 5244
rect 45928 5024 45980 5030
rect 45928 4966 45980 4972
rect 45940 4690 45968 4966
rect 45928 4684 45980 4690
rect 45928 4626 45980 4632
rect 45928 4276 45980 4282
rect 45928 4218 45980 4224
rect 45940 4078 45968 4218
rect 46032 4214 46060 5238
rect 46020 4208 46072 4214
rect 46020 4150 46072 4156
rect 45836 4072 45888 4078
rect 45836 4014 45888 4020
rect 45928 4072 45980 4078
rect 45928 4014 45980 4020
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45848 2446 45876 4014
rect 46020 2508 46072 2514
rect 46020 2450 46072 2456
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45480 82 45508 2382
rect 45558 96 45614 105
rect 45480 54 45558 82
rect 45558 31 45614 40
rect 45714 0 45826 800
rect 46032 785 46060 2450
rect 46216 2378 46244 5578
rect 46296 3528 46348 3534
rect 46296 3470 46348 3476
rect 46308 3398 46336 3470
rect 46296 3392 46348 3398
rect 46296 3334 46348 3340
rect 46400 3194 46428 13874
rect 46480 13864 46532 13870
rect 46480 13806 46532 13812
rect 46492 12306 46520 13806
rect 46664 13320 46716 13326
rect 46664 13262 46716 13268
rect 46676 12986 46704 13262
rect 46664 12980 46716 12986
rect 46664 12922 46716 12928
rect 46480 12300 46532 12306
rect 46480 12242 46532 12248
rect 46768 6322 46796 13874
rect 46940 13320 46992 13326
rect 46940 13262 46992 13268
rect 46952 12374 46980 13262
rect 47228 12434 47256 32370
rect 47320 19786 47348 45222
rect 47676 44804 47728 44810
rect 47676 44746 47728 44752
rect 47688 44538 47716 44746
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47584 44260 47636 44266
rect 47584 44202 47636 44208
rect 47596 40050 47624 44202
rect 47780 43314 47808 46378
rect 47872 46345 47900 46514
rect 47858 46336 47914 46345
rect 47858 46271 47914 46280
rect 47768 43308 47820 43314
rect 47768 43250 47820 43256
rect 47676 42628 47728 42634
rect 47676 42570 47728 42576
rect 47688 42362 47716 42570
rect 47676 42356 47728 42362
rect 47676 42298 47728 42304
rect 47768 41676 47820 41682
rect 47768 41618 47820 41624
rect 47780 41138 47808 41618
rect 47768 41132 47820 41138
rect 47768 41074 47820 41080
rect 47676 40520 47728 40526
rect 47676 40462 47728 40468
rect 47584 40044 47636 40050
rect 47584 39986 47636 39992
rect 47688 39574 47716 40462
rect 47676 39568 47728 39574
rect 47676 39510 47728 39516
rect 47860 38956 47912 38962
rect 47860 38898 47912 38904
rect 47872 38865 47900 38898
rect 47858 38856 47914 38865
rect 47858 38791 47914 38800
rect 47676 38276 47728 38282
rect 47676 38218 47728 38224
rect 47688 38010 47716 38218
rect 47676 38004 47728 38010
rect 47676 37946 47728 37952
rect 47492 37868 47544 37874
rect 47492 37810 47544 37816
rect 47400 29640 47452 29646
rect 47400 29582 47452 29588
rect 47412 29345 47440 29582
rect 47398 29336 47454 29345
rect 47398 29271 47454 29280
rect 47400 22500 47452 22506
rect 47400 22442 47452 22448
rect 47308 19780 47360 19786
rect 47308 19722 47360 19728
rect 47412 13274 47440 22442
rect 47504 21554 47532 37810
rect 47768 33516 47820 33522
rect 47768 33458 47820 33464
rect 47780 33425 47808 33458
rect 47766 33416 47822 33425
rect 47766 33351 47822 33360
rect 47860 33312 47912 33318
rect 47860 33254 47912 33260
rect 47676 32836 47728 32842
rect 47676 32778 47728 32784
rect 47688 32570 47716 32778
rect 47676 32564 47728 32570
rect 47676 32506 47728 32512
rect 47584 28076 47636 28082
rect 47584 28018 47636 28024
rect 47596 23730 47624 28018
rect 47676 27872 47728 27878
rect 47676 27814 47728 27820
rect 47688 27402 47716 27814
rect 47676 27396 47728 27402
rect 47676 27338 47728 27344
rect 47872 26586 47900 33254
rect 47860 26580 47912 26586
rect 47860 26522 47912 26528
rect 47768 25696 47820 25702
rect 47768 25638 47820 25644
rect 47780 24342 47808 25638
rect 47768 24336 47820 24342
rect 47768 24278 47820 24284
rect 47584 23724 47636 23730
rect 47584 23666 47636 23672
rect 47964 23594 47992 46854
rect 48044 46368 48096 46374
rect 48044 46310 48096 46316
rect 47952 23588 48004 23594
rect 47952 23530 48004 23536
rect 47676 23520 47728 23526
rect 47676 23462 47728 23468
rect 47688 23186 47716 23462
rect 47676 23180 47728 23186
rect 47676 23122 47728 23128
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47492 21548 47544 21554
rect 47492 21490 47544 21496
rect 47492 18284 47544 18290
rect 47492 18226 47544 18232
rect 47504 16574 47532 18226
rect 47596 17202 47624 22578
rect 47860 22568 47912 22574
rect 47860 22510 47912 22516
rect 47768 19168 47820 19174
rect 47768 19110 47820 19116
rect 47780 18834 47808 19110
rect 47768 18828 47820 18834
rect 47768 18770 47820 18776
rect 47676 18692 47728 18698
rect 47676 18634 47728 18640
rect 47688 18426 47716 18634
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47872 17678 47900 22510
rect 48056 17746 48084 46310
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48226 44976 48282 44985
rect 48136 44940 48188 44946
rect 48226 44911 48282 44920
rect 48136 44882 48188 44888
rect 48240 43858 48268 44911
rect 48228 43852 48280 43858
rect 48228 43794 48280 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 42265 48176 42570
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 48136 41608 48188 41614
rect 48134 41576 48136 41585
rect 48188 41576 48190 41585
rect 48134 41511 48190 41520
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48148 39506 48176 40151
rect 48136 39500 48188 39506
rect 48136 39442 48188 39448
rect 48136 38276 48188 38282
rect 48136 38218 48188 38224
rect 48148 38185 48176 38218
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48136 35080 48188 35086
rect 48136 35022 48188 35028
rect 48148 34785 48176 35022
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 48136 34604 48188 34610
rect 48136 34546 48188 34552
rect 48148 34105 48176 34546
rect 48134 34096 48190 34105
rect 48134 34031 48190 34040
rect 48136 32836 48188 32842
rect 48136 32778 48188 32784
rect 48148 32745 48176 32778
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48148 27538 48176 27911
rect 48136 27532 48188 27538
rect 48136 27474 48188 27480
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 25362 48176 25871
rect 48136 25356 48188 25362
rect 48136 25298 48188 25304
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48228 23044 48280 23050
rect 48228 22986 48280 22992
rect 48134 21176 48190 21185
rect 48134 21111 48190 21120
rect 48148 21010 48176 21111
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 48044 17740 48096 17746
rect 48044 17682 48096 17688
rect 47860 17672 47912 17678
rect 47860 17614 47912 17620
rect 48044 17604 48096 17610
rect 48044 17546 48096 17552
rect 47584 17196 47636 17202
rect 47584 17138 47636 17144
rect 47860 17196 47912 17202
rect 47860 17138 47912 17144
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47504 16546 47624 16574
rect 47412 13258 47532 13274
rect 47412 13252 47544 13258
rect 47412 13246 47492 13252
rect 47492 13194 47544 13200
rect 47044 12406 47256 12434
rect 46940 12368 46992 12374
rect 46940 12310 46992 12316
rect 46846 9616 46902 9625
rect 46846 9551 46848 9560
rect 46900 9551 46902 9560
rect 46848 9522 46900 9528
rect 46756 6316 46808 6322
rect 46756 6258 46808 6264
rect 46940 4684 46992 4690
rect 46940 4626 46992 4632
rect 46952 4049 46980 4626
rect 46938 4040 46994 4049
rect 46938 3975 46994 3984
rect 47044 3738 47072 12406
rect 47308 8968 47360 8974
rect 47308 8910 47360 8916
rect 47400 8968 47452 8974
rect 47400 8910 47452 8916
rect 47320 7585 47348 8910
rect 47412 7954 47440 8910
rect 47400 7948 47452 7954
rect 47400 7890 47452 7896
rect 47306 7576 47362 7585
rect 47306 7511 47362 7520
rect 47124 7200 47176 7206
rect 47124 7142 47176 7148
rect 47136 6866 47164 7142
rect 47124 6860 47176 6866
rect 47124 6802 47176 6808
rect 47504 4758 47532 13194
rect 47492 4752 47544 4758
rect 47492 4694 47544 4700
rect 47032 3732 47084 3738
rect 47032 3674 47084 3680
rect 47596 3670 47624 16546
rect 47688 16522 47716 16934
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47676 16108 47728 16114
rect 47676 16050 47728 16056
rect 47688 15502 47716 16050
rect 47676 15496 47728 15502
rect 47676 15438 47728 15444
rect 47768 15020 47820 15026
rect 47768 14962 47820 14968
rect 47780 14618 47808 14962
rect 47768 14612 47820 14618
rect 47768 14554 47820 14560
rect 47676 11076 47728 11082
rect 47676 11018 47728 11024
rect 47688 10810 47716 11018
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47872 9586 47900 17138
rect 48056 16574 48084 17546
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 47964 16546 48084 16574
rect 47860 9580 47912 9586
rect 47860 9522 47912 9528
rect 47766 8936 47822 8945
rect 47766 8871 47822 8880
rect 47780 8566 47808 8871
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 47964 7954 47992 16546
rect 48240 16425 48268 22986
rect 48226 16416 48282 16425
rect 48226 16351 48282 16360
rect 48044 16040 48096 16046
rect 48044 15982 48096 15988
rect 48056 15502 48084 15982
rect 48044 15496 48096 15502
rect 48044 15438 48096 15444
rect 48044 15360 48096 15366
rect 48044 15302 48096 15308
rect 47952 7948 48004 7954
rect 47952 7890 48004 7896
rect 47964 6474 47992 7890
rect 48056 6866 48084 15302
rect 48134 12336 48190 12345
rect 48134 12271 48136 12280
rect 48188 12271 48190 12280
rect 48136 12242 48188 12248
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 48136 7404 48188 7410
rect 48136 7346 48188 7352
rect 48148 6905 48176 7346
rect 48134 6896 48190 6905
rect 48044 6860 48096 6866
rect 48134 6831 48190 6840
rect 48044 6802 48096 6808
rect 47872 6446 47992 6474
rect 47872 5778 47900 6446
rect 47952 6112 48004 6118
rect 47952 6054 48004 6060
rect 47860 5772 47912 5778
rect 47780 5732 47860 5760
rect 47780 3942 47808 5732
rect 47860 5714 47912 5720
rect 47964 5302 47992 6054
rect 47952 5296 48004 5302
rect 47952 5238 48004 5244
rect 48056 5234 48084 6802
rect 48136 6316 48188 6322
rect 48136 6258 48188 6264
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 48044 5228 48096 5234
rect 48044 5170 48096 5176
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47584 3664 47636 3670
rect 47584 3606 47636 3612
rect 47766 3496 47822 3505
rect 47766 3431 47822 3440
rect 46388 3188 46440 3194
rect 46388 3130 46440 3136
rect 47780 3126 47808 3431
rect 47768 3120 47820 3126
rect 47768 3062 47820 3068
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 46388 2372 46440 2378
rect 46388 2314 46440 2320
rect 46400 800 46428 2314
rect 47044 800 47072 2450
rect 47688 800 47716 2926
rect 47872 1465 47900 5170
rect 48148 4185 48176 6258
rect 48134 4176 48190 4185
rect 48134 4111 48190 4120
rect 48320 4140 48372 4146
rect 48320 4082 48372 4088
rect 47858 1456 47914 1465
rect 47858 1391 47914 1400
rect 48332 800 48360 4082
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 48976 800 49004 3402
rect 46018 776 46074 785
rect 46018 711 46074 720
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 47640 1454 47696
rect 3698 46960 3754 47016
rect 1398 42880 1454 42936
rect 1398 40160 1454 40216
rect 1398 33396 1400 33416
rect 1400 33396 1452 33416
rect 1452 33396 1454 33416
rect 1398 33360 1454 33396
rect 1582 35400 1638 35456
rect 1306 32680 1362 32736
rect 1398 25236 1400 25256
rect 1400 25236 1452 25256
rect 1452 25236 1454 25256
rect 1398 25200 1454 25236
rect 1858 41520 1914 41576
rect 2778 46280 2834 46336
rect 3422 44920 3478 44976
rect 1858 32000 1914 32056
rect 1858 23160 1914 23216
rect 1398 17720 1454 17776
rect 1398 12280 1454 12336
rect 2778 36760 2834 36816
rect 2226 19080 2282 19136
rect 1950 16360 2006 16416
rect 2778 15000 2834 15056
rect 2778 10240 2834 10296
rect 3514 43560 3570 43616
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3790 39480 3846 39536
rect 3974 31320 4030 31376
rect 3974 28600 4030 28656
rect 3974 19760 4030 19816
rect 3882 18400 3938 18456
rect 3974 17076 3976 17096
rect 3976 17076 4028 17096
rect 4028 17076 4030 17096
rect 3974 17040 4030 17076
rect 3974 13676 3976 13696
rect 3976 13676 4028 13696
rect 4028 13676 4030 13696
rect 3974 13640 4030 13676
rect 3514 7520 3570 7576
rect 3422 6840 3478 6896
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3882 3984 3938 4040
rect 3422 3440 3478 3496
rect 3238 1400 3294 1456
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13082 25744 13138 25800
rect 19430 46960 19486 47016
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 21086 32836 21142 32872
rect 21086 32816 21088 32836
rect 21088 32816 21140 32836
rect 21140 32816 21142 32836
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19614 25916 19616 25936
rect 19616 25916 19668 25936
rect 19668 25916 19670 25936
rect 19614 25880 19670 25916
rect 19706 25220 19762 25256
rect 19706 25200 19708 25220
rect 19708 25200 19760 25220
rect 19760 25200 19762 25220
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 16854 3712 16910 3768
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19338 2896 19394 2952
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20166 3732 20222 3768
rect 20166 3712 20168 3732
rect 20168 3712 20220 3732
rect 20220 3712 20222 3732
rect 20442 2896 20498 2952
rect 22742 32716 22744 32736
rect 22744 32716 22796 32736
rect 22796 32716 22798 32736
rect 22742 32680 22798 32716
rect 22006 28484 22062 28520
rect 22006 28464 22008 28484
rect 22008 28464 22060 28484
rect 22060 28464 22062 28484
rect 24950 32836 25006 32872
rect 24950 32816 24952 32836
rect 24952 32816 25004 32836
rect 25004 32816 25006 32836
rect 27986 32680 28042 32736
rect 24306 26288 24362 26344
rect 23662 17856 23718 17912
rect 22006 3884 22008 3904
rect 22008 3884 22060 3904
rect 22060 3884 22062 3904
rect 22006 3848 22062 3884
rect 23754 2796 23756 2816
rect 23756 2796 23808 2816
rect 23808 2796 23810 2816
rect 23754 2760 23810 2796
rect 25134 25200 25190 25256
rect 24858 3848 24914 3904
rect 24950 2760 25006 2816
rect 25778 25744 25834 25800
rect 28262 32680 28318 32736
rect 28446 26288 28502 26344
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 30010 23568 30066 23624
rect 30746 24012 30748 24032
rect 30748 24012 30800 24032
rect 30800 24012 30802 24032
rect 30746 23976 30802 24012
rect 32126 26424 32182 26480
rect 32678 26288 32734 26344
rect 32862 23568 32918 23624
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 37830 26444 37886 26480
rect 37830 26424 37832 26444
rect 37832 26424 37884 26444
rect 37884 26424 37886 26444
rect 37738 23976 37794 24032
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38934 3732 38990 3768
rect 38934 3712 38936 3732
rect 38936 3712 38988 3732
rect 38988 3712 38990 3732
rect 38382 2896 38438 2952
rect 40130 2896 40186 2952
rect 41234 3712 41290 3768
rect 46846 47640 46902 47696
rect 46754 46960 46810 47016
rect 46110 39480 46166 39536
rect 46202 31320 46258 31376
rect 46202 25880 46258 25936
rect 46202 23160 46258 23216
rect 46846 40840 46902 40896
rect 46846 32000 46902 32056
rect 46846 29960 46902 30016
rect 46846 26560 46902 26616
rect 46202 22480 46258 22536
rect 46110 21800 46166 21856
rect 45558 8236 45560 8256
rect 45560 8236 45612 8256
rect 45612 8236 45614 8256
rect 45558 8200 45614 8236
rect 46846 25200 46902 25256
rect 46754 23840 46810 23896
rect 46386 18400 46442 18456
rect 46846 15680 46902 15736
rect 46202 6196 46204 6216
rect 46204 6196 46256 6216
rect 46256 6196 46258 6216
rect 46202 6160 46258 6196
rect 2870 720 2926 776
rect 45558 40 45614 96
rect 47858 46280 47914 46336
rect 47858 38800 47914 38856
rect 47398 29280 47454 29336
rect 47766 33360 47822 33416
rect 48134 45600 48190 45656
rect 48226 44920 48282 44976
rect 48134 42200 48190 42256
rect 48134 41556 48136 41576
rect 48136 41556 48188 41576
rect 48188 41556 48190 41576
rect 48134 41520 48190 41556
rect 48134 40160 48190 40216
rect 48134 38120 48190 38176
rect 48134 34720 48190 34776
rect 48134 34040 48190 34096
rect 48134 32680 48190 32736
rect 48134 27920 48190 27976
rect 48134 25880 48190 25936
rect 48134 24520 48190 24576
rect 48134 21120 48190 21176
rect 48134 19080 48190 19136
rect 46846 9580 46902 9616
rect 46846 9560 46848 9580
rect 46848 9560 46900 9580
rect 46900 9560 46902 9580
rect 46938 3984 46994 4040
rect 47306 7520 47362 7576
rect 48134 17040 48190 17096
rect 47766 8880 47822 8936
rect 48226 16360 48282 16416
rect 48134 12300 48190 12336
rect 48134 12280 48136 12300
rect 48136 12280 48188 12300
rect 48188 12280 48190 12300
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 6840 48190 6896
rect 47766 3440 47822 3496
rect 48134 4120 48190 4176
rect 47858 1400 47914 1456
rect 46018 720 46074 776
<< metal3 >>
rect 0 49588 800 49828
rect 0 48908 800 49148
rect 49200 48908 50000 49148
rect 0 48228 800 48468
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 46841 47698 46907 47701
rect 49200 47698 50000 47788
rect 46841 47696 50000 47698
rect 46841 47640 46846 47696
rect 46902 47640 50000 47696
rect 46841 47638 50000 47640
rect 46841 47635 46907 47638
rect 49200 47548 50000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3693 47018 3759 47021
rect 0 47016 3759 47018
rect 0 46960 3698 47016
rect 3754 46960 3759 47016
rect 0 46958 3759 46960
rect 0 46868 800 46958
rect 3693 46955 3759 46958
rect 19425 47018 19491 47021
rect 20110 47018 20116 47020
rect 19425 47016 20116 47018
rect 19425 46960 19430 47016
rect 19486 46960 20116 47016
rect 19425 46958 20116 46960
rect 19425 46955 19491 46958
rect 20110 46956 20116 46958
rect 20180 46956 20186 47020
rect 46749 47018 46815 47021
rect 49200 47018 50000 47108
rect 46749 47016 50000 47018
rect 46749 46960 46754 47016
rect 46810 46960 50000 47016
rect 46749 46958 50000 46960
rect 46749 46955 46815 46958
rect 49200 46868 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46428
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46188 800 46278
rect 2773 46275 2839 46278
rect 47853 46338 47919 46341
rect 49200 46338 50000 46428
rect 47853 46336 50000 46338
rect 47853 46280 47858 46336
rect 47914 46280 50000 46336
rect 47853 46278 50000 46280
rect 47853 46275 47919 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 49200 46188 50000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 48129 45658 48195 45661
rect 49200 45658 50000 45748
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45508 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 3417 44978 3483 44981
rect 0 44976 3483 44978
rect 0 44920 3422 44976
rect 3478 44920 3483 44976
rect 0 44918 3483 44920
rect 0 44828 800 44918
rect 3417 44915 3483 44918
rect 48221 44978 48287 44981
rect 49200 44978 50000 45068
rect 48221 44976 50000 44978
rect 48221 44920 48226 44976
rect 48282 44920 50000 44976
rect 48221 44918 50000 44920
rect 48221 44915 48287 44918
rect 49200 44828 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 49200 44148 50000 44388
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 3509 43618 3575 43621
rect 0 43616 3575 43618
rect 0 43560 3514 43616
rect 3570 43560 3575 43616
rect 0 43558 3575 43560
rect 0 43468 800 43558
rect 3509 43555 3575 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 49200 43468 50000 43708
rect 0 42938 800 43028
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42788 800 42878
rect 1393 42875 1459 42878
rect 49200 42788 50000 43028
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42108 800 42348
rect 48129 42258 48195 42261
rect 49200 42258 50000 42348
rect 48129 42256 50000 42258
rect 48129 42200 48134 42256
rect 48190 42200 50000 42256
rect 48129 42198 50000 42200
rect 48129 42195 48195 42198
rect 49200 42108 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41428 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40748 800 40988
rect 46841 40898 46907 40901
rect 49200 40898 50000 40988
rect 46841 40896 50000 40898
rect 46841 40840 46846 40896
rect 46902 40840 50000 40896
rect 46841 40838 50000 40840
rect 46841 40835 46907 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 49200 40748 50000 40838
rect 0 40218 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40068 800 40158
rect 1393 40155 1459 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40308
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40068 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39628
rect 3785 39538 3851 39541
rect 0 39536 3851 39538
rect 0 39480 3790 39536
rect 3846 39480 3851 39536
rect 0 39478 3851 39480
rect 0 39388 800 39478
rect 3785 39475 3851 39478
rect 46105 39538 46171 39541
rect 49200 39538 50000 39628
rect 46105 39536 50000 39538
rect 46105 39480 46110 39536
rect 46166 39480 50000 39536
rect 46105 39478 50000 39480
rect 46105 39475 46171 39478
rect 49200 39388 50000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38708 800 38948
rect 47853 38858 47919 38861
rect 49200 38858 50000 38948
rect 47853 38856 50000 38858
rect 47853 38800 47858 38856
rect 47914 38800 50000 38856
rect 47853 38798 50000 38800
rect 47853 38795 47919 38798
rect 49200 38708 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 49200 37348 50000 37588
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36908
rect 2773 36818 2839 36821
rect 0 36816 2839 36818
rect 0 36760 2778 36816
rect 2834 36760 2839 36816
rect 0 36758 2839 36760
rect 0 36668 800 36758
rect 2773 36755 2839 36758
rect 49200 36668 50000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 35988 800 36228
rect 49200 35988 50000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35458 800 35548
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35308 800 35398
rect 1577 35395 1643 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 48129 34778 48195 34781
rect 49200 34778 50000 34868
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34628 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 48129 34098 48195 34101
rect 49200 34098 50000 34188
rect 48129 34096 50000 34098
rect 48129 34040 48134 34096
rect 48190 34040 50000 34096
rect 48129 34038 50000 34040
rect 48129 34035 48195 34038
rect 49200 33948 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 0 33418 800 33508
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33268 800 33358
rect 1393 33355 1459 33358
rect 47761 33418 47827 33421
rect 49200 33418 50000 33508
rect 47761 33416 50000 33418
rect 47761 33360 47766 33416
rect 47822 33360 50000 33416
rect 47761 33358 50000 33360
rect 47761 33355 47827 33358
rect 49200 33268 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 21081 32874 21147 32877
rect 24945 32874 25011 32877
rect 21081 32872 25011 32874
rect 0 32738 800 32828
rect 21081 32816 21086 32872
rect 21142 32816 24950 32872
rect 25006 32816 25011 32872
rect 21081 32814 25011 32816
rect 21081 32811 21147 32814
rect 24945 32811 25011 32814
rect 1301 32738 1367 32741
rect 0 32736 1367 32738
rect 0 32680 1306 32736
rect 1362 32680 1367 32736
rect 0 32678 1367 32680
rect 0 32588 800 32678
rect 1301 32675 1367 32678
rect 22737 32738 22803 32741
rect 27981 32738 28047 32741
rect 28257 32738 28323 32741
rect 22737 32736 28323 32738
rect 22737 32680 22742 32736
rect 22798 32680 27986 32736
rect 28042 32680 28262 32736
rect 28318 32680 28323 32736
rect 22737 32678 28323 32680
rect 22737 32675 22803 32678
rect 27981 32675 28047 32678
rect 28257 32675 28323 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 49200 32588 50000 32678
rect 0 32058 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 46841 32058 46907 32061
rect 49200 32058 50000 32148
rect 46841 32056 50000 32058
rect 46841 32000 46846 32056
rect 46902 32000 50000 32056
rect 46841 31998 50000 32000
rect 46841 31995 46907 31998
rect 49200 31908 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31468
rect 3969 31378 4035 31381
rect 0 31376 4035 31378
rect 0 31320 3974 31376
rect 4030 31320 4035 31376
rect 0 31318 4035 31320
rect 0 31228 800 31318
rect 3969 31315 4035 31318
rect 46197 31378 46263 31381
rect 49200 31378 50000 31468
rect 46197 31376 50000 31378
rect 46197 31320 46202 31376
rect 46258 31320 50000 31376
rect 46197 31318 50000 31320
rect 46197 31315 46263 31318
rect 49200 31228 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 46841 30018 46907 30021
rect 49200 30018 50000 30108
rect 46841 30016 50000 30018
rect 46841 29960 46846 30016
rect 46902 29960 50000 30016
rect 46841 29958 50000 29960
rect 46841 29955 46907 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 49200 29868 50000 29958
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 47393 29338 47459 29341
rect 49200 29338 50000 29428
rect 47393 29336 50000 29338
rect 47393 29280 47398 29336
rect 47454 29280 50000 29336
rect 47393 29278 50000 29280
rect 47393 29275 47459 29278
rect 49200 29188 50000 29278
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28658 800 28748
rect 3969 28658 4035 28661
rect 49200 28658 50000 28748
rect 0 28656 4035 28658
rect 0 28600 3974 28656
rect 4030 28600 4035 28656
rect 0 28598 4035 28600
rect 0 28508 800 28598
rect 3969 28595 4035 28598
rect 45510 28598 50000 28658
rect 22001 28522 22067 28525
rect 45510 28522 45570 28598
rect 22001 28520 45570 28522
rect 22001 28464 22006 28520
rect 22062 28464 45570 28520
rect 49200 28508 50000 28598
rect 22001 28462 45570 28464
rect 22001 28459 22067 28462
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27148 800 27388
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 49200 27148 50000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 46841 26618 46907 26621
rect 49200 26618 50000 26708
rect 46841 26616 50000 26618
rect 46841 26560 46846 26616
rect 46902 26560 50000 26616
rect 46841 26558 50000 26560
rect 46841 26555 46907 26558
rect 32121 26482 32187 26485
rect 37825 26482 37891 26485
rect 32121 26480 37891 26482
rect 32121 26424 32126 26480
rect 32182 26424 37830 26480
rect 37886 26424 37891 26480
rect 49200 26468 50000 26558
rect 32121 26422 37891 26424
rect 32121 26419 32187 26422
rect 37825 26419 37891 26422
rect 24301 26346 24367 26349
rect 28441 26346 28507 26349
rect 32673 26346 32739 26349
rect 24301 26344 32739 26346
rect 24301 26288 24306 26344
rect 24362 26288 28446 26344
rect 28502 26288 32678 26344
rect 32734 26288 32739 26344
rect 24301 26286 32739 26288
rect 24301 26283 24367 26286
rect 28441 26283 28507 26286
rect 32673 26283 32739 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 19609 25938 19675 25941
rect 46197 25938 46263 25941
rect 19609 25936 46263 25938
rect 19609 25880 19614 25936
rect 19670 25880 46202 25936
rect 46258 25880 46263 25936
rect 19609 25878 46263 25880
rect 19609 25875 19675 25878
rect 46197 25875 46263 25878
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 13077 25802 13143 25805
rect 25773 25802 25839 25805
rect 13077 25800 25839 25802
rect 13077 25744 13082 25800
rect 13138 25744 25778 25800
rect 25834 25744 25839 25800
rect 49200 25788 50000 25878
rect 13077 25742 25839 25744
rect 13077 25739 13143 25742
rect 25773 25739 25839 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 19701 25258 19767 25261
rect 25129 25258 25195 25261
rect 19701 25256 25195 25258
rect 19701 25200 19706 25256
rect 19762 25200 25134 25256
rect 25190 25200 25195 25256
rect 19701 25198 25195 25200
rect 19701 25195 19767 25198
rect 25129 25195 25195 25198
rect 46841 25258 46907 25261
rect 49200 25258 50000 25348
rect 46841 25256 50000 25258
rect 46841 25200 46846 25256
rect 46902 25200 50000 25256
rect 46841 25198 50000 25200
rect 46841 25195 46907 25198
rect 49200 25108 50000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 0 24428 800 24668
rect 48129 24578 48195 24581
rect 49200 24578 50000 24668
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 49200 24428 50000 24518
rect 30741 24034 30807 24037
rect 37733 24034 37799 24037
rect 30741 24032 37799 24034
rect 0 23748 800 23988
rect 30741 23976 30746 24032
rect 30802 23976 37738 24032
rect 37794 23976 37799 24032
rect 30741 23974 37799 23976
rect 30741 23971 30807 23974
rect 37733 23971 37799 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 46749 23898 46815 23901
rect 49200 23898 50000 23988
rect 46749 23896 50000 23898
rect 46749 23840 46754 23896
rect 46810 23840 50000 23896
rect 46749 23838 50000 23840
rect 46749 23835 46815 23838
rect 49200 23748 50000 23838
rect 30005 23626 30071 23629
rect 32857 23626 32923 23629
rect 30005 23624 32923 23626
rect 30005 23568 30010 23624
rect 30066 23568 32862 23624
rect 32918 23568 32923 23624
rect 30005 23566 32923 23568
rect 30005 23563 30071 23566
rect 32857 23563 32923 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23308
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23068 800 23158
rect 1853 23155 1919 23158
rect 46197 23218 46263 23221
rect 49200 23218 50000 23308
rect 46197 23216 50000 23218
rect 46197 23160 46202 23216
rect 46258 23160 50000 23216
rect 46197 23158 50000 23160
rect 46197 23155 46263 23158
rect 49200 23068 50000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22388 800 22628
rect 46197 22538 46263 22541
rect 49200 22538 50000 22628
rect 46197 22536 50000 22538
rect 46197 22480 46202 22536
rect 46258 22480 50000 22536
rect 46197 22478 50000 22480
rect 46197 22475 46263 22478
rect 49200 22388 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21708 800 21948
rect 46105 21858 46171 21861
rect 49200 21858 50000 21948
rect 46105 21856 50000 21858
rect 46105 21800 46110 21856
rect 46166 21800 50000 21856
rect 46105 21798 50000 21800
rect 46105 21795 46171 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 48129 21178 48195 21181
rect 49200 21178 50000 21268
rect 48129 21176 50000 21178
rect 48129 21120 48134 21176
rect 48190 21120 50000 21176
rect 48129 21118 50000 21120
rect 48129 21115 48195 21118
rect 49200 21028 50000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19668 800 19758
rect 3969 19755 4035 19758
rect 49200 19668 50000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 19138 800 19228
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 18988 800 19078
rect 2221 19075 2287 19078
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3877 18458 3943 18461
rect 0 18456 3943 18458
rect 0 18400 3882 18456
rect 3938 18400 3943 18456
rect 0 18398 3943 18400
rect 0 18308 800 18398
rect 3877 18395 3943 18398
rect 46381 18458 46447 18461
rect 49200 18458 50000 18548
rect 46381 18456 50000 18458
rect 46381 18400 46386 18456
rect 46442 18400 50000 18456
rect 46381 18398 50000 18400
rect 46381 18395 46447 18398
rect 49200 18308 50000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 20110 17852 20116 17916
rect 20180 17914 20186 17916
rect 23657 17914 23723 17917
rect 20180 17912 23723 17914
rect 20180 17856 23662 17912
rect 23718 17856 23723 17912
rect 20180 17854 23723 17856
rect 20180 17852 20186 17854
rect 23657 17851 23723 17854
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 49200 17628 50000 17868
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 17098 800 17188
rect 3969 17098 4035 17101
rect 0 17096 4035 17098
rect 0 17040 3974 17096
rect 4030 17040 4035 17096
rect 0 17038 4035 17040
rect 0 16948 800 17038
rect 3969 17035 4035 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1945 16418 2011 16421
rect 0 16416 2011 16418
rect 0 16360 1950 16416
rect 2006 16360 2011 16416
rect 0 16358 2011 16360
rect 0 16268 800 16358
rect 1945 16355 2011 16358
rect 48221 16418 48287 16421
rect 49200 16418 50000 16508
rect 48221 16416 50000 16418
rect 48221 16360 48226 16416
rect 48282 16360 50000 16416
rect 48221 16358 50000 16360
rect 48221 16355 48287 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 49200 16268 50000 16358
rect 0 15588 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 46841 15738 46907 15741
rect 49200 15738 50000 15828
rect 46841 15736 50000 15738
rect 46841 15680 46846 15736
rect 46902 15680 50000 15736
rect 46841 15678 50000 15680
rect 46841 15675 46907 15678
rect 49200 15588 50000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 49200 14908 50000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 49200 14228 50000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13548 800 13638
rect 3969 13635 4035 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 49200 12868 50000 13108
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12428
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12188 800 12278
rect 1393 12275 1459 12278
rect 48129 12338 48195 12341
rect 49200 12338 50000 12428
rect 48129 12336 50000 12338
rect 48129 12280 48134 12336
rect 48190 12280 50000 12336
rect 48129 12278 50000 12280
rect 48129 12275 48195 12278
rect 49200 12188 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10148 800 10238
rect 2773 10235 2839 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9468 800 9708
rect 46841 9618 46907 9621
rect 49200 9618 50000 9708
rect 46841 9616 50000 9618
rect 46841 9560 46846 9616
rect 46902 9560 50000 9616
rect 46841 9558 50000 9560
rect 46841 9555 46907 9558
rect 49200 9468 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8788 800 9028
rect 47761 8938 47827 8941
rect 49200 8938 50000 9028
rect 47761 8936 50000 8938
rect 47761 8880 47766 8936
rect 47822 8880 50000 8936
rect 47761 8878 50000 8880
rect 47761 8875 47827 8878
rect 49200 8788 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8108 800 8348
rect 45553 8258 45619 8261
rect 49200 8258 50000 8348
rect 45553 8256 50000 8258
rect 45553 8200 45558 8256
rect 45614 8200 50000 8256
rect 45553 8198 50000 8200
rect 45553 8195 45619 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 3509 7578 3575 7581
rect 0 7576 3575 7578
rect 0 7520 3514 7576
rect 3570 7520 3575 7576
rect 0 7518 3575 7520
rect 0 7428 800 7518
rect 3509 7515 3575 7518
rect 47301 7578 47367 7581
rect 49200 7578 50000 7668
rect 47301 7576 50000 7578
rect 47301 7520 47306 7576
rect 47362 7520 50000 7576
rect 47301 7518 50000 7520
rect 47301 7515 47367 7518
rect 49200 7428 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 3417 6898 3483 6901
rect 0 6896 3483 6898
rect 0 6840 3422 6896
rect 3478 6840 3483 6896
rect 0 6838 3483 6840
rect 0 6748 800 6838
rect 3417 6835 3483 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6068 800 6308
rect 46197 6218 46263 6221
rect 49200 6218 50000 6308
rect 46197 6216 50000 6218
rect 46197 6160 46202 6216
rect 46258 6160 50000 6216
rect 46197 6158 50000 6160
rect 46197 6155 46263 6158
rect 49200 6068 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5388 800 5628
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 0 4708 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 49200 4708 50000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4028 800 4268
rect 48129 4178 48195 4181
rect 49200 4178 50000 4268
rect 48129 4176 50000 4178
rect 48129 4120 48134 4176
rect 48190 4120 50000 4176
rect 48129 4118 50000 4120
rect 48129 4115 48195 4118
rect 3877 4042 3943 4045
rect 46933 4042 46999 4045
rect 3877 4040 46999 4042
rect 3877 3984 3882 4040
rect 3938 3984 46938 4040
rect 46994 3984 46999 4040
rect 49200 4028 50000 4118
rect 3877 3982 46999 3984
rect 3877 3979 3943 3982
rect 46933 3979 46999 3982
rect 22001 3906 22067 3909
rect 24853 3906 24919 3909
rect 22001 3904 24919 3906
rect 22001 3848 22006 3904
rect 22062 3848 24858 3904
rect 24914 3848 24919 3904
rect 22001 3846 24919 3848
rect 22001 3843 22067 3846
rect 24853 3843 24919 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 16849 3770 16915 3773
rect 20161 3770 20227 3773
rect 16849 3768 20227 3770
rect 16849 3712 16854 3768
rect 16910 3712 20166 3768
rect 20222 3712 20227 3768
rect 16849 3710 20227 3712
rect 16849 3707 16915 3710
rect 20161 3707 20227 3710
rect 38929 3770 38995 3773
rect 41229 3770 41295 3773
rect 38929 3768 41295 3770
rect 38929 3712 38934 3768
rect 38990 3712 41234 3768
rect 41290 3712 41295 3768
rect 38929 3710 41295 3712
rect 38929 3707 38995 3710
rect 41229 3707 41295 3710
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 47761 3498 47827 3501
rect 49200 3498 50000 3588
rect 47761 3496 50000 3498
rect 47761 3440 47766 3496
rect 47822 3440 50000 3496
rect 47761 3438 50000 3440
rect 47761 3435 47827 3438
rect 49200 3348 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 19333 2954 19399 2957
rect 20437 2954 20503 2957
rect 19333 2952 20503 2954
rect 0 2668 800 2908
rect 19333 2896 19338 2952
rect 19394 2896 20442 2952
rect 20498 2896 20503 2952
rect 19333 2894 20503 2896
rect 19333 2891 19399 2894
rect 20437 2891 20503 2894
rect 38377 2954 38443 2957
rect 40125 2954 40191 2957
rect 38377 2952 40191 2954
rect 38377 2896 38382 2952
rect 38438 2896 40130 2952
rect 40186 2896 40191 2952
rect 38377 2894 40191 2896
rect 38377 2891 38443 2894
rect 40125 2891 40191 2894
rect 23749 2818 23815 2821
rect 24945 2818 25011 2821
rect 23749 2816 25011 2818
rect 23749 2760 23754 2816
rect 23810 2760 24950 2816
rect 25006 2760 25011 2816
rect 23749 2758 25011 2760
rect 23749 2755 23815 2758
rect 24945 2755 25011 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3233 1458 3299 1461
rect 0 1456 3299 1458
rect 0 1400 3238 1456
rect 3294 1400 3299 1456
rect 0 1398 3299 1400
rect 0 1308 800 1398
rect 3233 1395 3299 1398
rect 47853 1458 47919 1461
rect 49200 1458 50000 1548
rect 47853 1456 50000 1458
rect 47853 1400 47858 1456
rect 47914 1400 50000 1456
rect 47853 1398 50000 1400
rect 47853 1395 47919 1398
rect 49200 1308 50000 1398
rect 0 778 800 868
rect 2865 778 2931 781
rect 0 776 2931 778
rect 0 720 2870 776
rect 2926 720 2931 776
rect 0 718 2931 720
rect 0 628 800 718
rect 2865 715 2931 718
rect 46013 778 46079 781
rect 49200 778 50000 868
rect 46013 776 50000 778
rect 46013 720 46018 776
rect 46074 720 50000 776
rect 46013 718 50000 720
rect 46013 715 46079 718
rect 49200 628 50000 718
rect 45553 98 45619 101
rect 49200 98 50000 188
rect 45553 96 50000 98
rect 45553 40 45558 96
rect 45614 40 50000 96
rect 45553 38 50000 40
rect 45553 35 45619 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 20116 46956 20180 47020
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 20116 17852 20180 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 20115 47020 20181 47021
rect 20115 46956 20116 47020
rect 20180 46956 20181 47020
rect 20115 46955 20181 46956
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20118 17917 20178 46955
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 20115 17916 20181 17917
rect 20115 17852 20116 17916
rect 20180 17852 20181 17916
rect 20115 17851 20181 17852
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 27968 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 30452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_200 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1644511149
transform 1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_242
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1644511149
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1644511149
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1644511149
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1644511149
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1644511149
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_116
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1644511149
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_158
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1644511149
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1644511149
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_246
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_314
timestamp 1644511149
transform 1 0 29992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1644511149
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1644511149
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_414
timestamp 1644511149
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1644511149
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_88
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_107
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1644511149
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1644511149
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_231
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_238
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1644511149
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1644511149
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_399
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_405
timestamp 1644511149
transform 1 0 38364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_409
timestamp 1644511149
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_458
timestamp 1644511149
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_465
timestamp 1644511149
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_21
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1644511149
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1644511149
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_76
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_88
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_92
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_132
timestamp 1644511149
transform 1 0 13248 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1644511149
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp 1644511149
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_196
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_268
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_413
timestamp 1644511149
transform 1 0 39100 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_432
timestamp 1644511149
transform 1 0 40848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp 1644511149
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1644511149
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_185
timestamp 1644511149
transform 1 0 18124 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1644511149
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1644511149
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1644511149
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_242
timestamp 1644511149
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1644511149
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_451
timestamp 1644511149
transform 1 0 42596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_463
timestamp 1644511149
transform 1 0 43700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_468
timestamp 1644511149
transform 1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_481
timestamp 1644511149
transform 1 0 45356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_506
timestamp 1644511149
transform 1 0 47656 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_514
timestamp 1644511149
transform 1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_203
timestamp 1644511149
transform 1 0 19780 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1644511149
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_242
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_254
timestamp 1644511149
transform 1 0 24472 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_266
timestamp 1644511149
transform 1 0 25576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1644511149
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1644511149
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_479
timestamp 1644511149
transform 1 0 45172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_483
timestamp 1644511149
transform 1 0 45540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_512
timestamp 1644511149
transform 1 0 48208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1644511149
transform 1 0 46092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1644511149
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_512
timestamp 1644511149
transform 1 0 48208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_497
timestamp 1644511149
transform 1 0 46828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_512
timestamp 1644511149
transform 1 0 48208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_199
timestamp 1644511149
transform 1 0 19412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_211
timestamp 1644511149
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_500
timestamp 1644511149
transform 1 0 47104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_218
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp 1644511149
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1644511149
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_483
timestamp 1644511149
transform 1 0 45540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_487
timestamp 1644511149
transform 1 0 45908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1644511149
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_479
timestamp 1644511149
transform 1 0 45172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_488
timestamp 1644511149
transform 1 0 46000 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1644511149
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_217
timestamp 1644511149
transform 1 0 21068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1644511149
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1644511149
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_505
timestamp 1644511149
transform 1 0 47564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_200
timestamp 1644511149
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1644511149
transform 1 0 20608 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_481
timestamp 1644511149
transform 1 0 45356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_490
timestamp 1644511149
transform 1 0 46184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_14
timestamp 1644511149
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1644511149
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_204
timestamp 1644511149
transform 1 0 19872 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1644511149
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1644511149
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_226
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1644511149
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1644511149
transform 1 0 32292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1644511149
transform 1 0 33396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_464
timestamp 1644511149
transform 1 0 43792 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_495
timestamp 1644511149
transform 1 0 46644 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_504
timestamp 1644511149
transform 1 0 47472 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_246
timestamp 1644511149
transform 1 0 23736 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_258
timestamp 1644511149
transform 1 0 24840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_284
timestamp 1644511149
transform 1 0 27232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_308
timestamp 1644511149
transform 1 0 29440 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_320
timestamp 1644511149
transform 1 0 30544 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_482
timestamp 1644511149
transform 1 0 45448 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_490
timestamp 1644511149
transform 1 0 46184 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_494
timestamp 1644511149
transform 1 0 46552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1644511149
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_155
timestamp 1644511149
transform 1 0 15364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1644511149
transform 1 0 16468 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_171
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1644511149
transform 1 0 20056 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_230
timestamp 1644511149
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_267
timestamp 1644511149
transform 1 0 25668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_293
timestamp 1644511149
transform 1 0 28060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1644511149
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_330
timestamp 1644511149
transform 1 0 31464 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_342
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1644511149
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1644511149
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_430
timestamp 1644511149
transform 1 0 40664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_442
timestamp 1644511149
transform 1 0 41768 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_454
timestamp 1644511149
transform 1 0 42872 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_462
timestamp 1644511149
transform 1 0 43608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_468
timestamp 1644511149
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_483
timestamp 1644511149
transform 1 0 45540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_487
timestamp 1644511149
transform 1 0 45908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_504
timestamp 1644511149
transform 1 0 47472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_511
timestamp 1644511149
transform 1 0 48116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1644511149
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_153
timestamp 1644511149
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1644511149
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1644511149
transform 1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1644511149
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_262
timestamp 1644511149
transform 1 0 25208 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_268
timestamp 1644511149
transform 1 0 25760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1644511149
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_444
timestamp 1644511149
transform 1 0 41952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_486
timestamp 1644511149
transform 1 0 45816 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_510
timestamp 1644511149
transform 1 0 48024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_208
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_240
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_266
timestamp 1644511149
transform 1 0 25576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_275
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_284
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_296
timestamp 1644511149
transform 1 0 28336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1644511149
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1644511149
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_183
timestamp 1644511149
transform 1 0 17940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_228
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_240
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_256
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1644511149
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1644511149
transform 1 0 27416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1644511149
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1644511149
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1644511149
transform 1 0 15456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_168
timestamp 1644511149
transform 1 0 16560 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_232
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1644511149
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1644511149
transform 1 0 25944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_296
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_434
timestamp 1644511149
transform 1 0 41032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_446
timestamp 1644511149
transform 1 0 42136 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_458
timestamp 1644511149
transform 1 0 43240 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_470
timestamp 1644511149
transform 1 0 44344 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_146
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_228
timestamp 1644511149
transform 1 0 22080 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1644511149
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_266
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_269
timestamp 1644511149
transform 1 0 25852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_489
timestamp 1644511149
transform 1 0 46092 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_493
timestamp 1644511149
transform 1 0 46460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1644511149
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1644511149
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1644511149
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_152
timestamp 1644511149
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_216
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_228
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_235
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1644511149
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_256
timestamp 1644511149
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_268
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_322
timestamp 1644511149
transform 1 0 30728 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_334
timestamp 1644511149
transform 1 0 31832 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_346
timestamp 1644511149
transform 1 0 32936 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_486
timestamp 1644511149
transform 1 0 45816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_490
timestamp 1644511149
transform 1 0 46184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1644511149
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_92
timestamp 1644511149
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1644511149
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_156
timestamp 1644511149
transform 1 0 15456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1644511149
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_290
timestamp 1644511149
transform 1 0 27784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_302
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_314
timestamp 1644511149
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_452
timestamp 1644511149
transform 1 0 42688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_464
timestamp 1644511149
transform 1 0 43792 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_476
timestamp 1644511149
transform 1 0 44896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_482
timestamp 1644511149
transform 1 0 45448 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 1644511149
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1644511149
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_144
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_173
timestamp 1644511149
transform 1 0 17020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_218
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_224
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_230
timestamp 1644511149
transform 1 0 22264 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_242
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_259
timestamp 1644511149
transform 1 0 24932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_268
timestamp 1644511149
transform 1 0 25760 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_280
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_288
timestamp 1644511149
transform 1 0 27600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_295
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_317
timestamp 1644511149
transform 1 0 30268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_481
timestamp 1644511149
transform 1 0 45356 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1644511149
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1644511149
transform 1 0 8004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1644511149
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1644511149
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_191
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1644511149
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp 1644511149
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_255
timestamp 1644511149
transform 1 0 24564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_288
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_300
timestamp 1644511149
transform 1 0 28704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_459
timestamp 1644511149
transform 1 0 43332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_471
timestamp 1644511149
transform 1 0 44436 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_479
timestamp 1644511149
transform 1 0 45172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_495
timestamp 1644511149
transform 1 0 46644 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1644511149
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1644511149
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_146
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_225
timestamp 1644511149
transform 1 0 21804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_257
timestamp 1644511149
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_278
timestamp 1644511149
transform 1 0 26680 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_286
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_296
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_324
timestamp 1644511149
transform 1 0 30912 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1644511149
transform 1 0 42780 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_465
timestamp 1644511149
transform 1 0 43884 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_473
timestamp 1644511149
transform 1 0 44620 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_483
timestamp 1644511149
transform 1 0 45540 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1644511149
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1644511149
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_119
timestamp 1644511149
transform 1 0 12052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_133
timestamp 1644511149
transform 1 0 13340 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 1644511149
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1644511149
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_248
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_260
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1644511149
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_307
timestamp 1644511149
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_311
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_364
timestamp 1644511149
transform 1 0 34592 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_372
timestamp 1644511149
transform 1 0 35328 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_377
timestamp 1644511149
transform 1 0 35788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1644511149
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_430
timestamp 1644511149
transform 1 0 40664 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_442
timestamp 1644511149
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_479
timestamp 1644511149
transform 1 0 45172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_486
timestamp 1644511149
transform 1 0 45816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1644511149
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_508
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_106
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_114
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_152
timestamp 1644511149
transform 1 0 15088 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_168
timestamp 1644511149
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_179
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1644511149
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1644511149
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_271
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_275
timestamp 1644511149
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 1644511149
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_316
timestamp 1644511149
transform 1 0 30176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_328
timestamp 1644511149
transform 1 0 31280 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_340
timestamp 1644511149
transform 1 0 32384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_346
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_356
timestamp 1644511149
transform 1 0 33856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_385
timestamp 1644511149
transform 1 0 36524 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_397
timestamp 1644511149
transform 1 0 37628 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_409
timestamp 1644511149
transform 1 0 38732 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_440
timestamp 1644511149
transform 1 0 41584 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_456
timestamp 1644511149
transform 1 0 43056 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_468
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_481
timestamp 1644511149
transform 1 0 45356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_503
timestamp 1644511149
transform 1 0 47380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_510
timestamp 1644511149
transform 1 0 48024 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_78
timestamp 1644511149
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_103
timestamp 1644511149
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_133
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_141
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_145
timestamp 1644511149
transform 1 0 14444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_157
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1644511149
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_244
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_256
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_268
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_272
timestamp 1644511149
transform 1 0 26128 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_285
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_297
timestamp 1644511149
transform 1 0 28428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_309
timestamp 1644511149
transform 1 0 29532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1644511149
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_357
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_374
timestamp 1644511149
transform 1 0 35512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1644511149
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1644511149
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_396
timestamp 1644511149
transform 1 0 37536 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_408
timestamp 1644511149
transform 1 0 38640 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_420
timestamp 1644511149
transform 1 0 39744 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_432
timestamp 1644511149
transform 1 0 40848 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1644511149
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_470
timestamp 1644511149
transform 1 0 44344 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_478
timestamp 1644511149
transform 1 0 45080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1644511149
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1644511149
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_117
timestamp 1644511149
transform 1 0 11868 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_125
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_131
timestamp 1644511149
transform 1 0 13156 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_200
timestamp 1644511149
transform 1 0 19504 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_225
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_293
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1644511149
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_320
timestamp 1644511149
transform 1 0 30544 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_341
timestamp 1644511149
transform 1 0 32476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_349
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1644511149
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_374
timestamp 1644511149
transform 1 0 35512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_386
timestamp 1644511149
transform 1 0 36616 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_407
timestamp 1644511149
transform 1 0 38548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_437
timestamp 1644511149
transform 1 0 41308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_442
timestamp 1644511149
transform 1 0 41768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_452
timestamp 1644511149
transform 1 0 42688 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_464
timestamp 1644511149
transform 1 0 43792 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1644511149
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1644511149
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_117
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_126
timestamp 1644511149
transform 1 0 12696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_172
timestamp 1644511149
transform 1 0 16928 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_209
timestamp 1644511149
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_233
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_254
timestamp 1644511149
transform 1 0 24472 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_272
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_284
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_296
timestamp 1644511149
transform 1 0 28336 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_308
timestamp 1644511149
transform 1 0 29440 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_346
timestamp 1644511149
transform 1 0 32936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_358
timestamp 1644511149
transform 1 0 34040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_362
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_367
timestamp 1644511149
transform 1 0 34868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_378
timestamp 1644511149
transform 1 0 35880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_382
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_401
timestamp 1644511149
transform 1 0 37996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_408
timestamp 1644511149
transform 1 0 38640 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_420
timestamp 1644511149
transform 1 0 39744 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_432
timestamp 1644511149
transform 1 0 40848 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1644511149
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_88
timestamp 1644511149
transform 1 0 9200 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1644511149
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1644511149
transform 1 0 17664 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_204
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_230
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_276
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_283
timestamp 1644511149
transform 1 0 27140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1644511149
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_315
timestamp 1644511149
transform 1 0 30084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1644511149
transform 1 0 31188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_334
timestamp 1644511149
transform 1 0 31832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1644511149
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_349
timestamp 1644511149
transform 1 0 33212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1644511149
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_382
timestamp 1644511149
transform 1 0 36248 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_393
timestamp 1644511149
transform 1 0 37260 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_402
timestamp 1644511149
transform 1 0 38088 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1644511149
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_90
timestamp 1644511149
transform 1 0 9384 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_98
timestamp 1644511149
transform 1 0 10120 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1644511149
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_124
timestamp 1644511149
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_131
timestamp 1644511149
transform 1 0 13156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1644511149
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_209
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_215
timestamp 1644511149
transform 1 0 20884 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1644511149
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_240
timestamp 1644511149
transform 1 0 23184 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1644511149
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_255
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_321
timestamp 1644511149
transform 1 0 30636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1644511149
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_344
timestamp 1644511149
transform 1 0 32752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_353
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_365
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_397
timestamp 1644511149
transform 1 0 37628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_409
timestamp 1644511149
transform 1 0 38732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_421
timestamp 1644511149
transform 1 0 39836 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_433
timestamp 1644511149
transform 1 0 40940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1644511149
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_489
timestamp 1644511149
transform 1 0 46092 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_74
timestamp 1644511149
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1644511149
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_95
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_147
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_155
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_179
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_205
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_218
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_224
timestamp 1644511149
transform 1 0 21712 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1644511149
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_267
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_275
timestamp 1644511149
transform 1 0 26404 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_284
timestamp 1644511149
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_317
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_329
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_344
timestamp 1644511149
transform 1 0 32752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_352
timestamp 1644511149
transform 1 0 33488 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_359
timestamp 1644511149
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_373
timestamp 1644511149
transform 1 0 35420 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_385
timestamp 1644511149
transform 1 0 36524 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_391
timestamp 1644511149
transform 1 0 37076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_399
timestamp 1644511149
transform 1 0 37812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_412
timestamp 1644511149
transform 1 0 39008 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_63
timestamp 1644511149
transform 1 0 6900 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_88
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_100
timestamp 1644511149
transform 1 0 10304 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_116
timestamp 1644511149
transform 1 0 11776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_120
timestamp 1644511149
transform 1 0 12144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_124
timestamp 1644511149
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1644511149
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_136
timestamp 1644511149
transform 1 0 13616 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1644511149
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_151
timestamp 1644511149
transform 1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_234
timestamp 1644511149
transform 1 0 22632 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_238
timestamp 1644511149
transform 1 0 23000 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_290
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_299
timestamp 1644511149
transform 1 0 28612 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_303
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_319
timestamp 1644511149
transform 1 0 30452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_346
timestamp 1644511149
transform 1 0 32936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_350
timestamp 1644511149
transform 1 0 33304 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1644511149
transform 1 0 33764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_359
timestamp 1644511149
transform 1 0 34132 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_380
timestamp 1644511149
transform 1 0 36064 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_412
timestamp 1644511149
transform 1 0 39008 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_424
timestamp 1644511149
transform 1 0 40112 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_437
timestamp 1644511149
transform 1 0 41308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_445
timestamp 1644511149
transform 1 0 42044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_496
timestamp 1644511149
transform 1 0 46736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1644511149
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_69
timestamp 1644511149
transform 1 0 7452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1644511149
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_90
timestamp 1644511149
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_99
timestamp 1644511149
transform 1 0 10212 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_105
timestamp 1644511149
transform 1 0 10764 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_112
timestamp 1644511149
transform 1 0 11408 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_123
timestamp 1644511149
transform 1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1644511149
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_218
timestamp 1644511149
transform 1 0 21160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1644511149
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_337
timestamp 1644511149
transform 1 0 32108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_350
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_371
timestamp 1644511149
transform 1 0 35236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_383
timestamp 1644511149
transform 1 0 36340 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_395
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1644511149
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_429
timestamp 1644511149
transform 1 0 40572 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_437
timestamp 1644511149
transform 1 0 41308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_449
timestamp 1644511149
transform 1 0 42412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_461
timestamp 1644511149
transform 1 0 43516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_473
timestamp 1644511149
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_515
timestamp 1644511149
transform 1 0 48484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_82
timestamp 1644511149
transform 1 0 8648 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_92
timestamp 1644511149
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_96
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1644511149
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_153
timestamp 1644511149
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1644511149
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1644511149
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_209
timestamp 1644511149
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1644511149
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_284
timestamp 1644511149
transform 1 0 27232 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_288
timestamp 1644511149
transform 1 0 27600 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_311
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_319
timestamp 1644511149
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1644511149
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_358
timestamp 1644511149
transform 1 0 34040 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_364
timestamp 1644511149
transform 1 0 34592 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_368
timestamp 1644511149
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_380
timestamp 1644511149
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_410
timestamp 1644511149
transform 1 0 38824 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_422
timestamp 1644511149
transform 1 0 39928 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_434
timestamp 1644511149
transform 1 0 41032 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1644511149
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_69
timestamp 1644511149
transform 1 0 7452 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_94
timestamp 1644511149
transform 1 0 9752 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_113
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_125
timestamp 1644511149
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_129
timestamp 1644511149
transform 1 0 12972 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_200
timestamp 1644511149
transform 1 0 19504 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_224
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_261
timestamp 1644511149
transform 1 0 25116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_288
timestamp 1644511149
transform 1 0 27600 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_300
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_343
timestamp 1644511149
transform 1 0 32660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_351
timestamp 1644511149
transform 1 0 33396 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_400
timestamp 1644511149
transform 1 0 37904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_407
timestamp 1644511149
transform 1 0 38548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_73
timestamp 1644511149
transform 1 0 7820 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_95
timestamp 1644511149
transform 1 0 9844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 1644511149
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_117
timestamp 1644511149
transform 1 0 11868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1644511149
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_210
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1644511149
transform 1 0 23644 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_256
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_301
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_309
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_315
timestamp 1644511149
transform 1 0 30084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_323
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1644511149
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_347
timestamp 1644511149
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_354
timestamp 1644511149
transform 1 0 33672 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_366
timestamp 1644511149
transform 1 0 34776 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_374
timestamp 1644511149
transform 1 0 35512 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1644511149
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_403
timestamp 1644511149
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_415
timestamp 1644511149
transform 1 0 39284 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_427
timestamp 1644511149
transform 1 0 40388 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_439
timestamp 1644511149
transform 1 0 41492 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_500
timestamp 1644511149
transform 1 0 47104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1644511149
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_128
timestamp 1644511149
transform 1 0 12880 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_167
timestamp 1644511149
transform 1 0 16468 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_173
timestamp 1644511149
transform 1 0 17020 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1644511149
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1644511149
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_240
timestamp 1644511149
transform 1 0 23184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_244
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_257
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_286
timestamp 1644511149
transform 1 0 27416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_291
timestamp 1644511149
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_314
timestamp 1644511149
transform 1 0 29992 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_326
timestamp 1644511149
transform 1 0 31096 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_341
timestamp 1644511149
transform 1 0 32476 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_348
timestamp 1644511149
transform 1 0 33120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_352
timestamp 1644511149
transform 1 0 33488 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_369
timestamp 1644511149
transform 1 0 35052 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_373
timestamp 1644511149
transform 1 0 35420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_386
timestamp 1644511149
transform 1 0 36616 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_398
timestamp 1644511149
transform 1 0 37720 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_411
timestamp 1644511149
transform 1 0 38916 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_73
timestamp 1644511149
transform 1 0 7820 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_78
timestamp 1644511149
transform 1 0 8280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_82
timestamp 1644511149
transform 1 0 8648 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_89
timestamp 1644511149
transform 1 0 9292 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_120
timestamp 1644511149
transform 1 0 12144 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_128
timestamp 1644511149
transform 1 0 12880 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_150
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1644511149
transform 1 0 17572 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1644511149
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_215
timestamp 1644511149
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_229
timestamp 1644511149
transform 1 0 22172 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_254
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_264
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_288
timestamp 1644511149
transform 1 0 27600 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_301
timestamp 1644511149
transform 1 0 28796 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_309
timestamp 1644511149
transform 1 0 29532 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1644511149
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_363
timestamp 1644511149
transform 1 0 34500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_370
timestamp 1644511149
transform 1 0 35144 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1644511149
transform 1 0 36616 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_401
timestamp 1644511149
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_408
timestamp 1644511149
transform 1 0 38640 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_420
timestamp 1644511149
transform 1 0 39744 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_432
timestamp 1644511149
transform 1 0 40848 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_444
timestamp 1644511149
transform 1 0 41952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1644511149
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_105
timestamp 1644511149
transform 1 0 10764 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_111
timestamp 1644511149
transform 1 0 11316 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_115
timestamp 1644511149
transform 1 0 11684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_126
timestamp 1644511149
transform 1 0 12696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_134
timestamp 1644511149
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_159
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_163
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_171
timestamp 1644511149
transform 1 0 16836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_181
timestamp 1644511149
transform 1 0 17756 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_200
timestamp 1644511149
transform 1 0 19504 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_212
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_224
timestamp 1644511149
transform 1 0 21712 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_235
timestamp 1644511149
transform 1 0 22724 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_259
timestamp 1644511149
transform 1 0 24932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_266
timestamp 1644511149
transform 1 0 25576 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_274
timestamp 1644511149
transform 1 0 26312 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_279
timestamp 1644511149
transform 1 0 26772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_325
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_341
timestamp 1644511149
transform 1 0 32476 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_349
timestamp 1644511149
transform 1 0 33212 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_355
timestamp 1644511149
transform 1 0 33764 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_373
timestamp 1644511149
transform 1 0 35420 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_382
timestamp 1644511149
transform 1 0 36248 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_392
timestamp 1644511149
transform 1 0 37168 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_416
timestamp 1644511149
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_98
timestamp 1644511149
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1644511149
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_150
timestamp 1644511149
transform 1 0 14904 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_179
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_191
timestamp 1644511149
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_203
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_215
timestamp 1644511149
transform 1 0 20884 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_234
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_243
timestamp 1644511149
transform 1 0 23460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_247
timestamp 1644511149
transform 1 0 23828 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1644511149
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1644511149
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_302
timestamp 1644511149
transform 1 0 28888 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_320
timestamp 1644511149
transform 1 0 30544 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_331
timestamp 1644511149
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_340
timestamp 1644511149
transform 1 0 32384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_372
timestamp 1644511149
transform 1 0 35328 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_400
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_409
timestamp 1644511149
transform 1 0 38732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_421
timestamp 1644511149
transform 1 0 39836 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_433
timestamp 1644511149
transform 1 0 40940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_445
timestamp 1644511149
transform 1 0 42044 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_116
timestamp 1644511149
transform 1 0 11776 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_124
timestamp 1644511149
transform 1 0 12512 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_130
timestamp 1644511149
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1644511149
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_144
timestamp 1644511149
transform 1 0 14352 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_152
timestamp 1644511149
transform 1 0 15088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_166
timestamp 1644511149
transform 1 0 16376 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_185
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_200
timestamp 1644511149
transform 1 0 19504 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_230
timestamp 1644511149
transform 1 0 22264 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1644511149
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_268
timestamp 1644511149
transform 1 0 25760 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_278
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_312
timestamp 1644511149
transform 1 0 29808 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_320
timestamp 1644511149
transform 1 0 30544 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_328
timestamp 1644511149
transform 1 0 31280 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_336
timestamp 1644511149
transform 1 0 32016 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_342
timestamp 1644511149
transform 1 0 32568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_349
timestamp 1644511149
transform 1 0 33212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_359
timestamp 1644511149
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_383
timestamp 1644511149
transform 1 0 36340 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_392
timestamp 1644511149
transform 1 0 37168 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_404
timestamp 1644511149
transform 1 0 38272 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1644511149
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_14
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_26
timestamp 1644511149
transform 1 0 3496 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_38
timestamp 1644511149
transform 1 0 4600 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1644511149
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_96
timestamp 1644511149
transform 1 0 9936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_100
timestamp 1644511149
transform 1 0 10304 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1644511149
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_116
timestamp 1644511149
transform 1 0 11776 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1644511149
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_176
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_202
timestamp 1644511149
transform 1 0 19688 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1644511149
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_234
timestamp 1644511149
transform 1 0 22632 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_246
timestamp 1644511149
transform 1 0 23736 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_254
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1644511149
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_287
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_309
timestamp 1644511149
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_321
timestamp 1644511149
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1644511149
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_358
timestamp 1644511149
transform 1 0 34040 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_370
timestamp 1644511149
transform 1 0 35144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_382
timestamp 1644511149
transform 1 0 36248 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_396
timestamp 1644511149
transform 1 0 37536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_408
timestamp 1644511149
transform 1 0 38640 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_420
timestamp 1644511149
transform 1 0 39744 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_432
timestamp 1644511149
transform 1 0 40848 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1644511149
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1644511149
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_146
timestamp 1644511149
transform 1 0 14536 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_152
timestamp 1644511149
transform 1 0 15088 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_173
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_185
timestamp 1644511149
transform 1 0 18124 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1644511149
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_281
timestamp 1644511149
transform 1 0 26956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_341
timestamp 1644511149
transform 1 0 32476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_353
timestamp 1644511149
transform 1 0 33580 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_397
timestamp 1644511149
transform 1 0 37628 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_409
timestamp 1644511149
transform 1 0 38732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_417
timestamp 1644511149
transform 1 0 39468 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_507
timestamp 1644511149
transform 1 0 47748 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_515
timestamp 1644511149
transform 1 0 48484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_32
timestamp 1644511149
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_44
timestamp 1644511149
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_117
timestamp 1644511149
transform 1 0 11868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_132
timestamp 1644511149
transform 1 0 13248 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_144
timestamp 1644511149
transform 1 0 14352 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_150
timestamp 1644511149
transform 1 0 14904 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1644511149
transform 1 0 16928 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1644511149
transform 1 0 18032 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_244
timestamp 1644511149
transform 1 0 23552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_267
timestamp 1644511149
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_304
timestamp 1644511149
transform 1 0 29072 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_312
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1644511149
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_371
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_375
timestamp 1644511149
transform 1 0 35604 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_396
timestamp 1644511149
transform 1 0 37536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_408
timestamp 1644511149
transform 1 0 38640 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_420
timestamp 1644511149
transform 1 0 39744 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_432
timestamp 1644511149
transform 1 0 40848 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_444
timestamp 1644511149
transform 1 0 41952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1644511149
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1644511149
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_126
timestamp 1644511149
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1644511149
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_218
timestamp 1644511149
transform 1 0 21160 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_222
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_232
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_240
timestamp 1644511149
transform 1 0 23184 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_262
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_269
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_281
timestamp 1644511149
transform 1 0 26956 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1644511149
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_319
timestamp 1644511149
transform 1 0 30452 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_329
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_336
timestamp 1644511149
transform 1 0 32016 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_342
timestamp 1644511149
transform 1 0 32568 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_347
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1644511149
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1644511149
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_373
timestamp 1644511149
transform 1 0 35420 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1644511149
transform 1 0 36524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_397
timestamp 1644511149
transform 1 0 37628 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_409
timestamp 1644511149
transform 1 0 38732 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_417
timestamp 1644511149
transform 1 0 39468 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1644511149
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1644511149
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1644511149
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_197
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_201
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_213
timestamp 1644511149
transform 1 0 20700 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_236
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_240
timestamp 1644511149
transform 1 0 23184 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_244
timestamp 1644511149
transform 1 0 23552 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_268
timestamp 1644511149
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_289
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_321
timestamp 1644511149
transform 1 0 30636 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_344
timestamp 1644511149
transform 1 0 32752 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_356
timestamp 1644511149
transform 1 0 33856 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_368
timestamp 1644511149
transform 1 0 34960 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_380
timestamp 1644511149
transform 1 0 36064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_231
timestamp 1644511149
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_262
timestamp 1644511149
transform 1 0 25208 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_286
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_313
timestamp 1644511149
transform 1 0 29900 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_334
timestamp 1644511149
transform 1 0 31832 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_346
timestamp 1644511149
transform 1 0 32936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_358
timestamp 1644511149
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_497
timestamp 1644511149
transform 1 0 46828 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_312
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_321
timestamp 1644511149
transform 1 0 30636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1644511149
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_512
timestamp 1644511149
transform 1 0 48208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1644511149
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_28
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_40
timestamp 1644511149
transform 1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_494
timestamp 1644511149
transform 1 0 46552 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_502
timestamp 1644511149
transform 1 0 47288 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1644511149
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_494
timestamp 1644511149
transform 1 0 46552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_502
timestamp 1644511149
transform 1 0 47288 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_507
timestamp 1644511149
transform 1 0 47748 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_481
timestamp 1644511149
transform 1 0 45356 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_496
timestamp 1644511149
transform 1 0 46736 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_487
timestamp 1644511149
transform 1 0 45908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_481
timestamp 1644511149
transform 1 0 45356 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_494
timestamp 1644511149
transform 1 0 46552 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_502
timestamp 1644511149
transform 1 0 47288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_292
timestamp 1644511149
transform 1 0 27968 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1644511149
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_490
timestamp 1644511149
transform 1 0 46184 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_496
timestamp 1644511149
transform 1 0 46736 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_500
timestamp 1644511149
transform 1 0 47104 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_507
timestamp 1644511149
transform 1 0 47748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_515
timestamp 1644511149
transform 1 0 48484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_9
timestamp 1644511149
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_13
timestamp 1644511149
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_25
timestamp 1644511149
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_37
timestamp 1644511149
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1644511149
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_302
timestamp 1644511149
transform 1 0 28888 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_314
timestamp 1644511149
transform 1 0 29992 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_326
timestamp 1644511149
transform 1 0 31096 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_334
timestamp 1644511149
transform 1 0 31832 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_498
timestamp 1644511149
transform 1 0 46920 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_288
timestamp 1644511149
transform 1 0 27600 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_300
timestamp 1644511149
transform 1 0 28704 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1644511149
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1644511149
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_9
timestamp 1644511149
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_21
timestamp 1644511149
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_33
timestamp 1644511149
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1644511149
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_483
timestamp 1644511149
transform 1 0 45540 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_487
timestamp 1644511149
transform 1 0 45908 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_476
timestamp 1644511149
transform 1 0 44896 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_482
timestamp 1644511149
transform 1 0 45448 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_486
timestamp 1644511149
transform 1 0 45816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_14
timestamp 1644511149
transform 1 0 2392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1644511149
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_456
timestamp 1644511149
transform 1 0 43056 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_468
timestamp 1644511149
transform 1 0 44160 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_472
timestamp 1644511149
transform 1 0 44528 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1644511149
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_440
timestamp 1644511149
transform 1 0 41584 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_452
timestamp 1644511149
transform 1 0 42688 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_459
timestamp 1644511149
transform 1 0 43332 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_463
timestamp 1644511149
transform 1 0 43700 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_468
timestamp 1644511149
transform 1 0 44160 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_493
timestamp 1644511149
transform 1 0 46460 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_509
timestamp 1644511149
transform 1 0 47932 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_515
timestamp 1644511149
transform 1 0 48484 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1644511149
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_33
timestamp 1644511149
transform 1 0 4140 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_37
timestamp 1644511149
transform 1 0 4508 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_45
timestamp 1644511149
transform 1 0 5244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_57
timestamp 1644511149
transform 1 0 6348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_69
timestamp 1644511149
transform 1 0 7452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1644511149
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_117
timestamp 1644511149
transform 1 0 11868 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_130
timestamp 1644511149
transform 1 0 13064 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1644511149
transform 1 0 15456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1644511149
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_188
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1644511149
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_200
timestamp 1644511149
transform 1 0 19504 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_212
timestamp 1644511149
transform 1 0 20608 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_234
timestamp 1644511149
transform 1 0 22632 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_246
timestamp 1644511149
transform 1 0 23736 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1644511149
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_283
timestamp 1644511149
transform 1 0 27140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_336
timestamp 1644511149
transform 1 0 32016 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_348
timestamp 1644511149
transform 1 0 33120 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1644511149
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_406
timestamp 1644511149
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1644511149
transform 1 0 39560 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_7
timestamp 1644511149
transform 1 0 1748 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_19
timestamp 1644511149
transform 1 0 2852 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_218
timestamp 1644511149
transform 1 0 21160 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_228
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_240
timestamp 1644511149
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_252
timestamp 1644511149
transform 1 0 24288 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1644511149
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_315
timestamp 1644511149
transform 1 0 30084 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_327
timestamp 1644511149
transform 1 0 31188 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_358
timestamp 1644511149
transform 1 0 34040 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_370
timestamp 1644511149
transform 1 0 35144 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_382
timestamp 1644511149
transform 1 0 36248 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_390
timestamp 1644511149
transform 1 0 36984 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_401
timestamp 1644511149
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_423
timestamp 1644511149
transform 1 0 40020 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_431
timestamp 1644511149
transform 1 0 40756 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_437
timestamp 1644511149
transform 1 0 41308 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_444
timestamp 1644511149
transform 1 0 41952 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_470
timestamp 1644511149
transform 1 0 44344 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_478
timestamp 1644511149
transform 1 0 45080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1644511149
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1644511149
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_45
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_91
timestamp 1644511149
transform 1 0 9476 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_103
timestamp 1644511149
transform 1 0 10580 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_149
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_161
timestamp 1644511149
transform 1 0 15916 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_216
timestamp 1644511149
transform 1 0 20976 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_259
timestamp 1644511149
transform 1 0 24932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_266
timestamp 1644511149
transform 1 0 25576 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1644511149
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_315
timestamp 1644511149
transform 1 0 30084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_332
timestamp 1644511149
transform 1 0 31648 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1644511149
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1644511149
transform 1 0 40572 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_441
timestamp 1644511149
transform 1 0 41676 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_447
timestamp 1644511149
transform 1 0 42228 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1644511149
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_472
timestamp 1644511149
transform 1 0 44528 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1644511149
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_505
timestamp 1644511149
transform 1 0 47564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_511
timestamp 1644511149
transform 1 0 48116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_515
timestamp 1644511149
transform 1 0 48484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36616 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36616 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0620_
timestamp 1644511149
transform 1 0 31280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0621_
timestamp 1644511149
transform 1 0 32108 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0622_
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0623_
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0624_
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0625_
timestamp 1644511149
transform 1 0 30544 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0627_
timestamp 1644511149
transform 1 0 23000 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0628_
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0629_
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0630_
timestamp 1644511149
transform 1 0 23368 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0632_
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1644511149
transform 1 0 23000 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0636_
timestamp 1644511149
transform 1 0 10120 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0637_
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1644511149
transform 1 0 19412 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0640_
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 1644511149
transform 1 0 18124 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0642_
timestamp 1644511149
transform 1 0 18400 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0643_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0644_
timestamp 1644511149
transform 1 0 14628 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0646_
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0649_
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0650_
timestamp 1644511149
transform 1 0 17112 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0652_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1644511149
transform 1 0 15824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0656_
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0661_
timestamp 1644511149
transform 1 0 15364 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1644511149
transform 1 0 15456 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 1644511149
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0665_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0666_
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1644511149
transform 1 0 10672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0671_
timestamp 1644511149
transform 1 0 8924 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1644511149
transform 1 0 9844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0673_
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0674_
timestamp 1644511149
transform 1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0675_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0676_
timestamp 1644511149
transform 1 0 9016 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0677_
timestamp 1644511149
transform 1 0 8740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1644511149
transform 1 0 11408 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0682_
timestamp 1644511149
transform 1 0 9384 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0683_
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0685_
timestamp 1644511149
transform 1 0 7176 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0686_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0689_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 9752 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1644511149
transform 1 0 9568 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1644511149
transform 1 0 12144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0693_
timestamp 1644511149
transform 1 0 16652 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0694_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0695_
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0696_
timestamp 1644511149
transform 1 0 10856 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0699_
timestamp 1644511149
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0700_
timestamp 1644511149
transform 1 0 9568 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0702_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1644511149
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0707_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1644511149
transform 1 0 12328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0709_
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0710_
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _0711_
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0712_
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0713_
timestamp 1644511149
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1644511149
transform 1 0 11592 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0715_
timestamp 1644511149
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0717_
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0718_
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0720_
timestamp 1644511149
transform 1 0 12144 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0722_
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0723_
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0724_
timestamp 1644511149
transform 1 0 11500 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0725_
timestamp 1644511149
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0727_
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0728_
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1644511149
transform 1 0 16744 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0732_
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0733_
timestamp 1644511149
transform 1 0 17664 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1644511149
transform 1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0736_
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0737_
timestamp 1644511149
transform 1 0 17204 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0738_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 1644511149
transform 1 0 16928 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0742_
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0743_
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0744_
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0745_
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0746_
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0747_
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0749_
timestamp 1644511149
transform 1 0 20424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0750_
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1644511149
transform 1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1644511149
transform 1 0 20792 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0754_
timestamp 1644511149
transform 1 0 21160 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0757_
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_1  _0758_
timestamp 1644511149
transform 1 0 20424 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0759_
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0760_
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0762_
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0764_
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0765_
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0768_
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1644511149
transform 1 0 19872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1644511149
transform 1 0 19596 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1644511149
transform 1 0 20424 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0775_
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0776_
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1644511149
transform 1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0778_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1644511149
transform 1 0 24196 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0780_
timestamp 1644511149
transform 1 0 23552 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0782_
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0783_
timestamp 1644511149
transform 1 0 23552 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1644511149
transform 1 0 22448 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0787_
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0788_
timestamp 1644511149
transform 1 0 22356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0789_
timestamp 1644511149
transform 1 0 22172 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0790_
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0793_
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0794_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0795_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0797_
timestamp 1644511149
transform 1 0 22816 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0798_
timestamp 1644511149
transform 1 0 22080 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0800_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0801_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0802_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1644511149
transform 1 0 21988 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1644511149
transform 1 0 21620 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0805_
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0806_
timestamp 1644511149
transform 1 0 24840 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0807_
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1644511149
transform 1 0 27508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0809_
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0810_
timestamp 1644511149
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0811_
timestamp 1644511149
transform 1 0 25668 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0812_
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0813_
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0817_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0818_
timestamp 1644511149
transform 1 0 30084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0819_
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0820_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0822_
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0823_
timestamp 1644511149
transform 1 0 24472 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0825_
timestamp 1644511149
transform 1 0 22724 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0826_
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0827_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0828_
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0829_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0830_
timestamp 1644511149
transform 1 0 30544 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0831_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0833_
timestamp 1644511149
transform 1 0 25668 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0834_
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1644511149
transform 1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0839_
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1644511149
transform 1 0 26772 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0842_
timestamp 1644511149
transform 1 0 27600 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1644511149
transform 1 0 27140 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0844_
timestamp 1644511149
transform 1 0 27784 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0845_
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0846_
timestamp 1644511149
transform 1 0 25300 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0847_
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0849_
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0852_
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0853_
timestamp 1644511149
transform 1 0 31280 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0854_
timestamp 1644511149
transform 1 0 30820 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0855_
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1644511149
transform 1 0 28152 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0858_
timestamp 1644511149
transform 1 0 27968 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0859_
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0860_
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0861_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0862_
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0863_
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0864_
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0865_
timestamp 1644511149
transform 1 0 33396 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0866_
timestamp 1644511149
transform 1 0 34868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1644511149
transform 1 0 34408 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0868_
timestamp 1644511149
transform 1 0 32752 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 33396 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 1644511149
transform 1 0 32292 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33580 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0872_
timestamp 1644511149
transform 1 0 38088 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0873_
timestamp 1644511149
transform 1 0 38456 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0875_
timestamp 1644511149
transform 1 0 32384 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0876_
timestamp 1644511149
transform 1 0 30912 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0877_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0879_
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0880_
timestamp 1644511149
transform 1 0 30452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0881_
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0882_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0883_
timestamp 1644511149
transform 1 0 30268 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0884_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28888 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0885_
timestamp 1644511149
transform 1 0 29624 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0886_
timestamp 1644511149
transform 1 0 33120 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0888_
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0889_
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0890_
timestamp 1644511149
transform 1 0 33120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1644511149
transform 1 0 33856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0893_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0894_
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0895_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1644511149
transform 1 0 31924 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1644511149
transform 1 0 33396 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1644511149
transform 1 0 31096 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0899_
timestamp 1644511149
transform 1 0 32108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0900_
timestamp 1644511149
transform 1 0 29716 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _0901_
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0904_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0905_
timestamp 1644511149
transform 1 0 28428 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0906_
timestamp 1644511149
transform 1 0 27876 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0907_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0908_
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0909_
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1644511149
transform 1 0 30360 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0912_
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0913_
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1644511149
transform 1 0 36708 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1644511149
transform 1 0 35880 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0916_
timestamp 1644511149
transform 1 0 35144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 1644511149
transform 1 0 35604 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0920_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1644511149
transform 1 0 38272 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0922_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1644511149
transform 1 0 36064 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0924_
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 1644511149
transform 1 0 35696 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp 1644511149
transform 1 0 35696 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1644511149
transform 1 0 36340 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0929_
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0930_
timestamp 1644511149
transform 1 0 36708 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0931_
timestamp 1644511149
transform 1 0 38548 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0932_
timestamp 1644511149
transform 1 0 37444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0933_
timestamp 1644511149
transform 1 0 35236 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1644511149
transform 1 0 34684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1644511149
transform 1 0 35880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0938_
timestamp 1644511149
transform 1 0 35880 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0939_
timestamp 1644511149
transform 1 0 37628 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0940_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0941_
timestamp 1644511149
transform 1 0 23828 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1644511149
transform 1 0 22448 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0944_
timestamp 1644511149
transform 1 0 41400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0945_
timestamp 1644511149
transform 1 0 42780 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 43884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1644511149
transform 1 0 43516 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 45264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0957_
timestamp 1644511149
transform 1 0 41676 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1644511149
transform 1 0 12052 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0963_
timestamp 1644511149
transform 1 0 41952 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1644511149
transform 1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0969_
timestamp 1644511149
transform 1 0 40756 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40112 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 31188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1644511149
transform 1 0 40388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 45540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0976_
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 14904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0982_
timestamp 1644511149
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 8004 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 7544 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0988_
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1644511149
transform 1 0 12420 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0994_
timestamp 1644511149
transform 1 0 40204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp 1644511149
transform 1 0 41308 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1000_
timestamp 1644511149
transform 1 0 44988 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _1001_
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1007_
timestamp 1644511149
transform 1 0 45632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1644511149
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1013_
timestamp 1644511149
transform 1 0 45080 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 46460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 27324 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1019_
timestamp 1644511149
transform 1 0 45724 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 4968 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1025_
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 46644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1031_
timestamp 1644511149
transform 1 0 41400 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1032_
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 9016 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1644511149
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 8096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1038_
timestamp 1644511149
transform 1 0 19596 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 19320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42136 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 43056 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1050_
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1644511149
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1056_
timestamp 1644511149
transform 1 0 10304 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1644511149
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1644511149
transform 1 0 41308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1063_
timestamp 1644511149
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1064_
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _1066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1644511149
transform 1 0 45448 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1644511149
transform 1 0 45172 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1644511149
transform 1 0 45632 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1071_
timestamp 1644511149
transform 1 0 46276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1644511149
transform 1 0 47840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1644511149
transform 1 0 25944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1644511149
transform 1 0 25392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1076_
timestamp 1644511149
transform 1 0 27784 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46368 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1080_
timestamp 1644511149
transform 1 0 46552 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1081_
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1644511149
transform 1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45540 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45816 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1085_
timestamp 1644511149
transform 1 0 45540 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1086_
timestamp 1644511149
transform 1 0 46368 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45540 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1088_
timestamp 1644511149
transform 1 0 47012 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1089_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1090_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 1644511149
transform 1 0 45632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45908 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1093_
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1095_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1096_
timestamp 1644511149
transform 1 0 26036 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1099_
timestamp 1644511149
transform 1 0 26772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _1100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1101_
timestamp 1644511149
transform 1 0 26036 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1102_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1103_
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1644511149
transform 1 0 45540 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45448 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1106_
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1107_
timestamp 1644511149
transform 1 0 44804 0 -1 40256
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1108_
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1644511149
transform 1 0 35512 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1112_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform 1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1644511149
transform 1 0 33672 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1644511149
transform 1 0 34684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1124_
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1644511149
transform 1 0 32936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 31096 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1130_
timestamp 1644511149
transform 1 0 26128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1644511149
transform 1 0 27232 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1644511149
transform 1 0 28336 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1644511149
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1136_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1644511149
transform 1 0 26496 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1644511149
transform 1 0 25576 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1644511149
transform 1 0 25576 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1142_
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1644511149
transform 1 0 21528 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1644511149
transform 1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1147_
timestamp 1644511149
transform 1 0 20516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1148_
timestamp 1644511149
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1149_
timestamp 1644511149
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1150_
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1151_
timestamp 1644511149
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1152_
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1154_
timestamp 1644511149
transform 1 0 19136 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1155_
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1156_
timestamp 1644511149
transform 1 0 16928 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1157_
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1158_
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1159_
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1160_
timestamp 1644511149
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1161_
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1162_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1163_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1165_
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1644511149
transform 1 0 10304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1169_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1170_
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1171_
timestamp 1644511149
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1172_
timestamp 1644511149
transform 1 0 6532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1173_
timestamp 1644511149
transform 1 0 10396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1174_
timestamp 1644511149
transform 1 0 7912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1175_
timestamp 1644511149
transform 1 0 11776 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1644511149
transform 1 0 10028 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1177_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1178_
timestamp 1644511149
transform 1 0 12696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1644511149
transform 1 0 14628 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1180_
timestamp 1644511149
transform 1 0 14260 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1181_
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1182_
timestamp 1644511149
transform 1 0 18124 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36708 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1644511149
transform 1 0 37536 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1644511149
transform 1 0 36064 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1644511149
transform 1 0 32660 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1644511149
transform 1 0 29992 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1644511149
transform 1 0 32200 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1644511149
transform 1 0 34224 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1644511149
transform 1 0 33488 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1644511149
transform 1 0 32200 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1644511149
transform 1 0 24840 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1644511149
transform 1 0 25300 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1644511149
transform 1 0 25668 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1644511149
transform 1 0 23920 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1644511149
transform 1 0 24564 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1644511149
transform 1 0 20424 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1644511149
transform 1 0 20056 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1218_
timestamp 1644511149
transform 1 0 22448 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1219_
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1220_
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1222_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1225_
timestamp 1644511149
transform 1 0 16652 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1226_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1229_
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1230_
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1232_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1233_
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1235_
timestamp 1644511149
transform 1 0 9936 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1644511149
transform 1 0 7544 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1238_
timestamp 1644511149
transform 1 0 7268 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1241_
timestamp 1644511149
transform 1 0 9660 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1242_
timestamp 1644511149
transform 1 0 11684 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1243_
timestamp 1644511149
transform 1 0 12880 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1248_
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1249_
timestamp 1644511149
transform 1 0 18400 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1250__81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1251__82
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1252__83
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1253__84
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1254__85
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1255__86
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1256__87
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1257__88
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1258__89
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1259__90
timestamp 1644511149
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1260__91
timestamp 1644511149
transform 1 0 47748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1261__92
timestamp 1644511149
transform 1 0 1840 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1262__93
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1263__94
timestamp 1644511149
transform 1 0 4232 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1264__95
timestamp 1644511149
transform 1 0 1472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1265__96
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1266__97
timestamp 1644511149
transform 1 0 45540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1267__98
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1268__99
timestamp 1644511149
transform 1 0 45632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1269__100
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1270__101
timestamp 1644511149
transform 1 0 38088 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1271__102
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1272__103
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1273__104
timestamp 1644511149
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1274__105
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1275__106
timestamp 1644511149
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1276__107
timestamp 1644511149
transform 1 0 47472 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1277__108
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1278__109
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1279__110
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1280__111
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1281__112
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1282__113
timestamp 1644511149
transform 1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1283__114
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1284__115
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1285__116
timestamp 1644511149
transform 1 0 42780 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1286__117
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1287__118
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1288__119
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1289__120
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1290__121
timestamp 1644511149
transform 1 0 45632 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1291__122
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1292__123
timestamp 1644511149
transform 1 0 47472 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1293__124
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1294__125
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1295__126
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1296__127
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1297__128
timestamp 1644511149
transform 1 0 47472 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1298__129
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1299__130
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1300__131
timestamp 1644511149
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1301__132
timestamp 1644511149
transform 1 0 45080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1302__133
timestamp 1644511149
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1303__134
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1304__135
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41216 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1309_
timestamp 1644511149
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1310_
timestamp 1644511149
transform 1 0 45724 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1311_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1312_
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1313_
timestamp 1644511149
transform 1 0 38732 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1314_
timestamp 1644511149
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1315_
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1316_
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1317_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1318_
timestamp 1644511149
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1319_
timestamp 1644511149
transform 1 0 20700 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1320_
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1321_
timestamp 1644511149
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1322_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1323_
timestamp 1644511149
transform 1 0 25208 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1324_
timestamp 1644511149
transform 1 0 46276 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1325_
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1326_
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1327_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1328_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1329_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1330_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1331_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1332_
timestamp 1644511149
transform 1 0 46276 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1333_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1334_
timestamp 1644511149
transform 1 0 38088 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1335_
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1336_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1337_
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1338_
timestamp 1644511149
transform 1 0 45448 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1339_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1340_
timestamp 1644511149
transform 1 0 19412 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1341_
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1342_
timestamp 1644511149
transform 1 0 30360 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1343_
timestamp 1644511149
transform 1 0 19504 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1344_
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1345_
timestamp 1644511149
transform 1 0 40020 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1346_
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1347_
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1348_
timestamp 1644511149
transform 1 0 16560 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1349_
timestamp 1644511149
transform 1 0 9200 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1350_
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1351_
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1352_
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1353_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1354_
timestamp 1644511149
transform 1 0 15640 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1355_
timestamp 1644511149
transform 1 0 8832 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1356_
timestamp 1644511149
transform 1 0 12696 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1357_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1358_
timestamp 1644511149
transform 1 0 9568 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1359_
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1360_
timestamp 1644511149
transform 1 0 7912 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1361_
timestamp 1644511149
transform 1 0 8740 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1362_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1363_
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1364_
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1365_
timestamp 1644511149
transform 1 0 20148 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1366_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1367_
timestamp 1644511149
transform 1 0 12972 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1368_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1369_
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1370_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1371_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1372_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1373_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1374_
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1375_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1376_
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1377_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1378_
timestamp 1644511149
transform 1 0 41216 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1379_
timestamp 1644511149
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1380_
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1381_
timestamp 1644511149
transform 1 0 42596 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1382_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1383_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1384_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1385_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1386_
timestamp 1644511149
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1387_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1388_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1389_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1390_
timestamp 1644511149
transform 1 0 45172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1391_
timestamp 1644511149
transform 1 0 19228 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1392_
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1393_
timestamp 1644511149
transform 1 0 45172 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1394_
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1395_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1396_
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1397_
timestamp 1644511149
transform 1 0 45172 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1398_
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1399_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1400_
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 33396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 33580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 47932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1644511149
transform 1 0 29716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 47932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1644511149
transform 1 0 46184 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 47288 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1644511149
transform 1 0 47656 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1644511149
transform 1 0 35512 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1644511149
transform 1 0 47748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1644511149
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1644511149
transform 1 0 9108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 44896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1644511149
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1644511149
transform 1 0 17020 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1644511149
transform 1 0 47656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 40204 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 30728 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 43792 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1644511149
transform 1 0 26496 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 46184 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 46184 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 46828 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 24380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 47932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 47932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.bypass1._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.bypass2._0_
timestamp 1644511149
transform 1 0 41308 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_1  instrumented_adder.control1._0_
timestamp 1644511149
transform 1 0 38456 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.control2._0_
timestamp 1644511149
transform 1 0 39560 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[0\]._0_
timestamp 1644511149
transform 1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[1\]._0_
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[2\]._0_
timestamp 1644511149
transform 1 0 39192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.control_inverters\[3\]._0_
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[0\]._0_
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[1\]._0_
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[2\]._0_
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[3\]._0_
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[4\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[5\]._0_
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[6\]._0_
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[7\]._0_
timestamp 1644511149
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[8\]._0_
timestamp 1644511149
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[9\]._0_
timestamp 1644511149
transform 1 0 18216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[10\]._0_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[11\]._0_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[12\]._0_
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[13\]._0_
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[14\]._0_
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[15\]._0_
timestamp 1644511149
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[16\]._0_
timestamp 1644511149
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[17\]._0_
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[18\]._0_
timestamp 1644511149
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[19\]._0_
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[20\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[21\]._0_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[22\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[23\]._0_
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[24\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[25\]._0_
timestamp 1644511149
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[26\]._0_
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[27\]._0_
timestamp 1644511149
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[28\]._0_
timestamp 1644511149
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[29\]._0_
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  instrumented_adder.inverters\[30\]._0_
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[0\]._0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 28152 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ext_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 47012 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 29348 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ext_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[0\]._0_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[1\]._0_
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[2\]._0_
timestamp 1644511149
transform 1 0 2116 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[3\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[4\]._0_
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  instrumented_adder.tristate_ring_inputs\[5\]._0_
timestamp 1644511149
transform 1 0 45908 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[6\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_ring_inputs\[7\]._0_
timestamp 1644511149
transform 1 0 42872 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[0\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[1\]._0_
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[2\]._0_
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[3\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[4\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[5\]._0_
timestamp 1644511149
transform 1 0 45172 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[6\]._0_
timestamp 1644511149
transform 1 0 46276 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  instrumented_adder.tristate_sum_outputs\[7\]._0_
timestamp 1644511149
transform 1 0 26036 0 1 40256
box -38 -48 1970 592
<< labels >>
rlabel metal3 s 49200 38708 50000 38948 6 active
port 0 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[0]
port 1 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[10]
port 2 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[11]
port 3 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 la1_data_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 33948 50000 34188 6 la1_data_in[13]
port 5 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[14]
port 6 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[15]
port 7 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 la1_data_in[16]
port 8 nsew signal input
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_in[17]
port 9 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la1_data_in[18]
port 10 nsew signal input
rlabel metal3 s 49200 4028 50000 4268 6 la1_data_in[19]
port 11 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[1]
port 12 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 la1_data_in[20]
port 13 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_data_in[21]
port 14 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_data_in[22]
port 15 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 628 50000 868 6 la1_data_in[24]
port 17 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_data_in[25]
port 18 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[26]
port 19 nsew signal input
rlabel metal3 s 49200 46188 50000 46428 6 la1_data_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 29188 50000 29428 6 la1_data_in[28]
port 21 nsew signal input
rlabel metal3 s 49200 23068 50000 23308 6 la1_data_in[29]
port 22 nsew signal input
rlabel metal2 s 5142 0 5254 800 6 la1_data_in[2]
port 23 nsew signal input
rlabel metal3 s 49200 7428 50000 7668 6 la1_data_in[30]
port 24 nsew signal input
rlabel metal2 s 1922 49200 2034 50000 6 la1_data_in[31]
port 25 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[3]
port 26 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[4]
port 27 nsew signal input
rlabel metal3 s 49200 33268 50000 33508 6 la1_data_in[5]
port 28 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_data_in[6]
port 29 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 la1_data_in[7]
port 30 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[8]
port 31 nsew signal input
rlabel metal2 s 35410 0 35522 800 6 la1_data_in[9]
port 32 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[0]
port 33 nsew signal bidirectional
rlabel metal2 s 32190 49200 32302 50000 6 la1_data_out[10]
port 34 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la1_data_out[11]
port 35 nsew signal bidirectional
rlabel metal3 s 49200 38028 50000 38268 6 la1_data_out[12]
port 36 nsew signal bidirectional
rlabel metal3 s 49200 27828 50000 28068 6 la1_data_out[13]
port 37 nsew signal bidirectional
rlabel metal2 s 21242 49200 21354 50000 6 la1_data_out[14]
port 38 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[15]
port 39 nsew signal bidirectional
rlabel metal2 s 25106 49200 25218 50000 6 la1_data_out[16]
port 40 nsew signal bidirectional
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_out[17]
port 41 nsew signal bidirectional
rlabel metal2 s 25750 49200 25862 50000 6 la1_data_out[18]
port 42 nsew signal bidirectional
rlabel metal3 s 49200 16268 50000 16508 6 la1_data_out[19]
port 43 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 la1_data_out[1]
port 44 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 la1_data_out[20]
port 45 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 la1_data_out[21]
port 46 nsew signal bidirectional
rlabel metal2 s 3854 49200 3966 50000 6 la1_data_out[22]
port 47 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[23]
port 48 nsew signal bidirectional
rlabel metal2 s 43138 0 43250 800 6 la1_data_out[24]
port 49 nsew signal bidirectional
rlabel metal2 s 47002 49200 47114 50000 6 la1_data_out[25]
port 50 nsew signal bidirectional
rlabel metal3 s 49200 47548 50000 47788 6 la1_data_out[26]
port 51 nsew signal bidirectional
rlabel metal3 s 49200 21028 50000 21268 6 la1_data_out[27]
port 52 nsew signal bidirectional
rlabel metal3 s 49200 41428 50000 41668 6 la1_data_out[28]
port 53 nsew signal bidirectional
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_out[29]
port 54 nsew signal bidirectional
rlabel metal2 s 45070 0 45182 800 6 la1_data_out[2]
port 55 nsew signal bidirectional
rlabel metal2 s 7718 0 7830 800 6 la1_data_out[30]
port 56 nsew signal bidirectional
rlabel metal2 s 42494 49200 42606 50000 6 la1_data_out[31]
port 57 nsew signal bidirectional
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[3]
port 58 nsew signal bidirectional
rlabel metal3 s 49200 25788 50000 26028 6 la1_data_out[4]
port 59 nsew signal bidirectional
rlabel metal2 s 3854 0 3966 800 6 la1_data_out[5]
port 60 nsew signal bidirectional
rlabel metal3 s 49200 39388 50000 39628 6 la1_data_out[6]
port 61 nsew signal bidirectional
rlabel metal2 s 27038 49200 27150 50000 6 la1_data_out[7]
port 62 nsew signal bidirectional
rlabel metal2 s 39918 49200 40030 50000 6 la1_data_out[8]
port 63 nsew signal bidirectional
rlabel metal3 s 49200 12188 50000 12428 6 la1_data_out[9]
port 64 nsew signal bidirectional
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[0]
port 65 nsew signal input
rlabel metal3 s 49200 19668 50000 19908 6 la1_oenb[10]
port 66 nsew signal input
rlabel metal3 s 49200 13548 50000 13788 6 la1_oenb[11]
port 67 nsew signal input
rlabel metal3 s 49200 27148 50000 27388 6 la1_oenb[12]
port 68 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[13]
port 69 nsew signal input
rlabel metal3 s 49200 43468 50000 43708 6 la1_oenb[14]
port 70 nsew signal input
rlabel metal2 s 19310 49200 19422 50000 6 la1_oenb[15]
port 71 nsew signal input
rlabel metal2 s 24462 49200 24574 50000 6 la1_oenb[16]
port 72 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[17]
port 73 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[18]
port 74 nsew signal input
rlabel metal3 s 49200 4708 50000 4948 6 la1_oenb[19]
port 75 nsew signal input
rlabel metal3 s 49200 48228 50000 48468 6 la1_oenb[1]
port 76 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[20]
port 77 nsew signal input
rlabel metal2 s 22530 49200 22642 50000 6 la1_oenb[21]
port 78 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[22]
port 79 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_oenb[23]
port 80 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la1_oenb[24]
port 81 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la1_oenb[25]
port 82 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_oenb[26]
port 83 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la1_oenb[27]
port 84 nsew signal input
rlabel metal3 s 0 8108 800 8348 6 la1_oenb[28]
port 85 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 la1_oenb[29]
port 86 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[2]
port 87 nsew signal input
rlabel metal3 s 49200 30548 50000 30788 6 la1_oenb[30]
port 88 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 la1_oenb[31]
port 89 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_oenb[3]
port 90 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_oenb[4]
port 91 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_oenb[5]
port 92 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[6]
port 93 nsew signal input
rlabel metal3 s 49200 42788 50000 43028 6 la1_oenb[7]
port 94 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la1_oenb[8]
port 95 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_oenb[9]
port 96 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 la2_data_in[0]
port 97 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la2_data_in[10]
port 98 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_data_in[11]
port 99 nsew signal input
rlabel metal2 s 43782 49200 43894 50000 6 la2_data_in[12]
port 100 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la2_data_in[13]
port 101 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la2_data_in[14]
port 102 nsew signal input
rlabel metal2 s 47646 49200 47758 50000 6 la2_data_in[15]
port 103 nsew signal input
rlabel metal3 s 49200 -52 50000 188 6 la2_data_in[16]
port 104 nsew signal input
rlabel metal3 s 49200 31908 50000 32148 6 la2_data_in[17]
port 105 nsew signal input
rlabel metal2 s 9006 49200 9118 50000 6 la2_data_in[18]
port 106 nsew signal input
rlabel metal3 s 49200 1308 50000 1548 6 la2_data_in[19]
port 107 nsew signal input
rlabel metal3 s 49200 21708 50000 21948 6 la2_data_in[1]
port 108 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la2_data_in[20]
port 109 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la2_data_in[21]
port 110 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la2_data_in[22]
port 111 nsew signal input
rlabel metal2 s 45714 49200 45826 50000 6 la2_data_in[23]
port 112 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la2_data_in[24]
port 113 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la2_data_in[25]
port 114 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 la2_data_in[26]
port 115 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la2_data_in[27]
port 116 nsew signal input
rlabel metal2 s 13514 49200 13626 50000 6 la2_data_in[28]
port 117 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la2_data_in[29]
port 118 nsew signal input
rlabel metal3 s 0 12188 800 12428 6 la2_data_in[2]
port 119 nsew signal input
rlabel metal3 s 49200 3348 50000 3588 6 la2_data_in[30]
port 120 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la2_data_in[31]
port 121 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 la2_data_in[3]
port 122 nsew signal input
rlabel metal2 s 30902 49200 31014 50000 6 la2_data_in[4]
port 123 nsew signal input
rlabel metal2 s 44426 49200 44538 50000 6 la2_data_in[5]
port 124 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la2_data_in[6]
port 125 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la2_data_in[7]
port 126 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 la2_data_in[8]
port 127 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la2_data_in[9]
port 128 nsew signal input
rlabel metal3 s 49200 26468 50000 26708 6 la2_data_out[0]
port 129 nsew signal bidirectional
rlabel metal3 s 49200 31228 50000 31468 6 la2_data_out[10]
port 130 nsew signal bidirectional
rlabel metal2 s -10 49200 102 50000 6 la2_data_out[11]
port 131 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la2_data_out[12]
port 132 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[13]
port 133 nsew signal bidirectional
rlabel metal3 s 0 43468 800 43708 6 la2_data_out[14]
port 134 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la2_data_out[15]
port 135 nsew signal bidirectional
rlabel metal2 s 15446 49200 15558 50000 6 la2_data_out[16]
port 136 nsew signal bidirectional
rlabel metal2 s 17378 49200 17490 50000 6 la2_data_out[17]
port 137 nsew signal bidirectional
rlabel metal3 s 0 16948 800 17188 6 la2_data_out[18]
port 138 nsew signal bidirectional
rlabel metal2 s 8362 49200 8474 50000 6 la2_data_out[19]
port 139 nsew signal bidirectional
rlabel metal3 s 49200 46868 50000 47108 6 la2_data_out[1]
port 140 nsew signal bidirectional
rlabel metal3 s 0 13548 800 13788 6 la2_data_out[20]
port 141 nsew signal bidirectional
rlabel metal2 s 18666 0 18778 800 6 la2_data_out[21]
port 142 nsew signal bidirectional
rlabel metal3 s 49200 29868 50000 30108 6 la2_data_out[22]
port 143 nsew signal bidirectional
rlabel metal3 s 0 28508 800 28748 6 la2_data_out[23]
port 144 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[24]
port 145 nsew signal bidirectional
rlabel metal2 s 41206 49200 41318 50000 6 la2_data_out[25]
port 146 nsew signal bidirectional
rlabel metal2 s 19310 0 19422 800 6 la2_data_out[26]
port 147 nsew signal bidirectional
rlabel metal2 s 37986 49200 38098 50000 6 la2_data_out[27]
port 148 nsew signal bidirectional
rlabel metal3 s 49200 28508 50000 28748 6 la2_data_out[28]
port 149 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la2_data_out[29]
port 150 nsew signal bidirectional
rlabel metal3 s 0 1308 800 1548 6 la2_data_out[2]
port 151 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la2_data_out[30]
port 152 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la2_data_out[31]
port 153 nsew signal bidirectional
rlabel metal3 s 0 3348 800 3588 6 la2_data_out[3]
port 154 nsew signal bidirectional
rlabel metal3 s 0 6748 800 6988 6 la2_data_out[4]
port 155 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[5]
port 156 nsew signal bidirectional
rlabel metal2 s 14802 0 14914 800 6 la2_data_out[6]
port 157 nsew signal bidirectional
rlabel metal3 s 0 7428 800 7668 6 la2_data_out[7]
port 158 nsew signal bidirectional
rlabel metal3 s 49200 8108 50000 8348 6 la2_data_out[8]
port 159 nsew signal bidirectional
rlabel metal3 s 49200 15588 50000 15828 6 la2_data_out[9]
port 160 nsew signal bidirectional
rlabel metal2 s 34766 49200 34878 50000 6 la2_oenb[0]
port 161 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la2_oenb[10]
port 162 nsew signal input
rlabel metal2 s 27682 49200 27794 50000 6 la2_oenb[11]
port 163 nsew signal input
rlabel metal3 s 49200 14908 50000 15148 6 la2_oenb[12]
port 164 nsew signal input
rlabel metal3 s 49200 44148 50000 44388 6 la2_oenb[13]
port 165 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la2_oenb[14]
port 166 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la2_oenb[15]
port 167 nsew signal input
rlabel metal3 s 49200 36668 50000 36908 6 la2_oenb[16]
port 168 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la2_oenb[17]
port 169 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la2_oenb[18]
port 170 nsew signal input
rlabel metal2 s 36698 0 36810 800 6 la2_oenb[19]
port 171 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la2_oenb[1]
port 172 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la2_oenb[20]
port 173 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[21]
port 174 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la2_oenb[22]
port 175 nsew signal input
rlabel metal3 s 49200 17628 50000 17868 6 la2_oenb[23]
port 176 nsew signal input
rlabel metal3 s 0 15588 800 15828 6 la2_oenb[24]
port 177 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la2_oenb[25]
port 178 nsew signal input
rlabel metal2 s 36698 49200 36810 50000 6 la2_oenb[26]
port 179 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_oenb[27]
port 180 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la2_oenb[28]
port 181 nsew signal input
rlabel metal2 s 33478 49200 33590 50000 6 la2_oenb[29]
port 182 nsew signal input
rlabel metal3 s 0 1988 800 2228 6 la2_oenb[2]
port 183 nsew signal input
rlabel metal3 s 0 27148 800 27388 6 la2_oenb[30]
port 184 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la2_oenb[31]
port 185 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 la2_oenb[3]
port 186 nsew signal input
rlabel metal2 s 49578 49200 49690 50000 6 la2_oenb[4]
port 187 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la2_oenb[5]
port 188 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la2_oenb[6]
port 189 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la2_oenb[7]
port 190 nsew signal input
rlabel metal2 s 10294 49200 10406 50000 6 la2_oenb[8]
port 191 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la2_oenb[9]
port 192 nsew signal input
rlabel metal3 s 49200 22388 50000 22628 6 la3_data_in[0]
port 193 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la3_data_in[10]
port 194 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 la3_data_in[11]
port 195 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 la3_data_in[12]
port 196 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[13]
port 197 nsew signal input
rlabel metal2 s 46358 49200 46470 50000 6 la3_data_in[14]
port 198 nsew signal input
rlabel metal3 s 49200 40748 50000 40988 6 la3_data_in[15]
port 199 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la3_data_in[16]
port 200 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la3_data_in[17]
port 201 nsew signal input
rlabel metal3 s 49200 2668 50000 2908 6 la3_data_in[18]
port 202 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la3_data_in[19]
port 203 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la3_data_in[1]
port 204 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_data_in[20]
port 205 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 la3_data_in[21]
port 206 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la3_data_in[22]
port 207 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_in[23]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la3_data_in[24]
port 209 nsew signal input
rlabel metal3 s 49200 48908 50000 49148 6 la3_data_in[25]
port 210 nsew signal input
rlabel metal3 s 49200 12868 50000 13108 6 la3_data_in[26]
port 211 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la3_data_in[27]
port 212 nsew signal input
rlabel metal2 s 48934 49200 49046 50000 6 la3_data_in[28]
port 213 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la3_data_in[29]
port 214 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la3_data_in[2]
port 215 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la3_data_in[30]
port 216 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_data_in[31]
port 217 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 la3_data_in[3]
port 218 nsew signal input
rlabel metal2 s 28326 49200 28438 50000 6 la3_data_in[4]
port 219 nsew signal input
rlabel metal3 s 49200 34628 50000 34868 6 la3_data_in[5]
port 220 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la3_data_in[6]
port 221 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la3_data_in[7]
port 222 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la3_data_in[8]
port 223 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la3_data_in[9]
port 224 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la3_data_out[0]
port 225 nsew signal bidirectional
rlabel metal3 s 49200 18988 50000 19228 6 la3_data_out[10]
port 226 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la3_data_out[11]
port 227 nsew signal bidirectional
rlabel metal2 s 43138 49200 43250 50000 6 la3_data_out[12]
port 228 nsew signal bidirectional
rlabel metal3 s 49200 45508 50000 45748 6 la3_data_out[13]
port 229 nsew signal bidirectional
rlabel metal2 s 14158 49200 14270 50000 6 la3_data_out[14]
port 230 nsew signal bidirectional
rlabel metal2 s 6430 0 6542 800 6 la3_data_out[15]
port 231 nsew signal bidirectional
rlabel metal3 s 0 628 800 868 6 la3_data_out[16]
port 232 nsew signal bidirectional
rlabel metal3 s 49200 44828 50000 45068 6 la3_data_out[17]
port 233 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 la3_data_out[18]
port 234 nsew signal bidirectional
rlabel metal3 s 49200 32588 50000 32828 6 la3_data_out[19]
port 235 nsew signal bidirectional
rlabel metal3 s 49200 10828 50000 11068 6 la3_data_out[1]
port 236 nsew signal bidirectional
rlabel metal3 s 0 16268 800 16508 6 la3_data_out[20]
port 237 nsew signal bidirectional
rlabel metal2 s 48290 49200 48402 50000 6 la3_data_out[21]
port 238 nsew signal bidirectional
rlabel metal2 s 20598 49200 20710 50000 6 la3_data_out[22]
port 239 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 la3_data_out[23]
port 240 nsew signal bidirectional
rlabel metal3 s 49200 25108 50000 25348 6 la3_data_out[24]
port 241 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 la3_data_out[25]
port 242 nsew signal bidirectional
rlabel metal3 s 49200 10148 50000 10388 6 la3_data_out[26]
port 243 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 la3_data_out[27]
port 244 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la3_data_out[28]
port 245 nsew signal bidirectional
rlabel metal2 s 7074 0 7186 800 6 la3_data_out[29]
port 246 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[2]
port 247 nsew signal bidirectional
rlabel metal3 s 49200 16948 50000 17188 6 la3_data_out[30]
port 248 nsew signal bidirectional
rlabel metal2 s 45070 49200 45182 50000 6 la3_data_out[31]
port 249 nsew signal bidirectional
rlabel metal3 s 49200 40068 50000 40308 6 la3_data_out[3]
port 250 nsew signal bidirectional
rlabel metal2 s 48934 0 49046 800 6 la3_data_out[4]
port 251 nsew signal bidirectional
rlabel metal3 s 0 14908 800 15148 6 la3_data_out[5]
port 252 nsew signal bidirectional
rlabel metal3 s 49200 24428 50000 24668 6 la3_data_out[6]
port 253 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la3_data_out[7]
port 254 nsew signal bidirectional
rlabel metal3 s 49200 42108 50000 42348 6 la3_data_out[8]
port 255 nsew signal bidirectional
rlabel metal2 s 41850 49200 41962 50000 6 la3_data_out[9]
port 256 nsew signal bidirectional
rlabel metal3 s 49200 1988 50000 2228 6 la3_oenb[0]
port 257 nsew signal input
rlabel metal2 s 40562 49200 40674 50000 6 la3_oenb[10]
port 258 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la3_oenb[11]
port 259 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[12]
port 260 nsew signal input
rlabel metal2 s 31546 0 31658 800 6 la3_oenb[13]
port 261 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 262 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la3_oenb[15]
port 263 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la3_oenb[16]
port 264 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la3_oenb[17]
port 265 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_oenb[18]
port 266 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[19]
port 267 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la3_oenb[1]
port 268 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_oenb[20]
port 269 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la3_oenb[21]
port 270 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la3_oenb[22]
port 271 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 la3_oenb[23]
port 272 nsew signal input
rlabel metal2 s 37342 49200 37454 50000 6 la3_oenb[24]
port 273 nsew signal input
rlabel metal3 s 49200 11508 50000 11748 6 la3_oenb[25]
port 274 nsew signal input
rlabel metal3 s 0 35988 800 36228 6 la3_oenb[26]
port 275 nsew signal input
rlabel metal3 s 49200 37348 50000 37588 6 la3_oenb[27]
port 276 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la3_oenb[28]
port 277 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la3_oenb[29]
port 278 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 279 nsew signal input
rlabel metal3 s 49200 35988 50000 36228 6 la3_oenb[30]
port 280 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la3_oenb[31]
port 281 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 la3_oenb[3]
port 282 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la3_oenb[4]
port 283 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la3_oenb[5]
port 284 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la3_oenb[6]
port 285 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la3_oenb[7]
port 286 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la3_oenb[8]
port 287 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_oenb[9]
port 288 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 289 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 290 nsew ground input
rlabel metal3 s 49200 23748 50000 23988 6 wb_clk_i
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
