magic
tech sky130A
magscale 1 2
timestamp 1654618827
<< obsli1 >>
rect 1104 2159 74888 73457
<< obsm1 >>
rect 198 1300 75426 73488
<< metal2 >>
rect -10 75200 102 76000
rect 634 75200 746 76000
rect 1922 75200 2034 76000
rect 2566 75200 2678 76000
rect 3210 75200 3322 76000
rect 3854 75200 3966 76000
rect 4498 75200 4610 76000
rect 5142 75200 5254 76000
rect 5786 75200 5898 76000
rect 6430 75200 6542 76000
rect 7718 75200 7830 76000
rect 8362 75200 8474 76000
rect 9006 75200 9118 76000
rect 9650 75200 9762 76000
rect 10294 75200 10406 76000
rect 10938 75200 11050 76000
rect 11582 75200 11694 76000
rect 12870 75200 12982 76000
rect 13514 75200 13626 76000
rect 14158 75200 14270 76000
rect 14802 75200 14914 76000
rect 15446 75200 15558 76000
rect 16090 75200 16202 76000
rect 16734 75200 16846 76000
rect 18022 75200 18134 76000
rect 18666 75200 18778 76000
rect 19310 75200 19422 76000
rect 19954 75200 20066 76000
rect 20598 75200 20710 76000
rect 21242 75200 21354 76000
rect 21886 75200 21998 76000
rect 23174 75200 23286 76000
rect 23818 75200 23930 76000
rect 24462 75200 24574 76000
rect 25106 75200 25218 76000
rect 25750 75200 25862 76000
rect 26394 75200 26506 76000
rect 27038 75200 27150 76000
rect 27682 75200 27794 76000
rect 28970 75200 29082 76000
rect 29614 75200 29726 76000
rect 30258 75200 30370 76000
rect 30902 75200 31014 76000
rect 31546 75200 31658 76000
rect 32190 75200 32302 76000
rect 32834 75200 32946 76000
rect 34122 75200 34234 76000
rect 34766 75200 34878 76000
rect 35410 75200 35522 76000
rect 36054 75200 36166 76000
rect 36698 75200 36810 76000
rect 37342 75200 37454 76000
rect 37986 75200 38098 76000
rect 39274 75200 39386 76000
rect 39918 75200 40030 76000
rect 40562 75200 40674 76000
rect 41206 75200 41318 76000
rect 41850 75200 41962 76000
rect 42494 75200 42606 76000
rect 43138 75200 43250 76000
rect 44426 75200 44538 76000
rect 45070 75200 45182 76000
rect 45714 75200 45826 76000
rect 46358 75200 46470 76000
rect 47002 75200 47114 76000
rect 47646 75200 47758 76000
rect 48290 75200 48402 76000
rect 49578 75200 49690 76000
rect 50222 75200 50334 76000
rect 50866 75200 50978 76000
rect 51510 75200 51622 76000
rect 52154 75200 52266 76000
rect 52798 75200 52910 76000
rect 53442 75200 53554 76000
rect 54086 75200 54198 76000
rect 55374 75200 55486 76000
rect 56018 75200 56130 76000
rect 56662 75200 56774 76000
rect 57306 75200 57418 76000
rect 57950 75200 58062 76000
rect 58594 75200 58706 76000
rect 59238 75200 59350 76000
rect 60526 75200 60638 76000
rect 61170 75200 61282 76000
rect 61814 75200 61926 76000
rect 62458 75200 62570 76000
rect 63102 75200 63214 76000
rect 63746 75200 63858 76000
rect 64390 75200 64502 76000
rect 65678 75200 65790 76000
rect 66322 75200 66434 76000
rect 66966 75200 67078 76000
rect 67610 75200 67722 76000
rect 68254 75200 68366 76000
rect 68898 75200 69010 76000
rect 69542 75200 69654 76000
rect 70830 75200 70942 76000
rect 71474 75200 71586 76000
rect 72118 75200 72230 76000
rect 72762 75200 72874 76000
rect 73406 75200 73518 76000
rect 74050 75200 74162 76000
rect 74694 75200 74806 76000
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
rect 50222 0 50334 800
rect 50866 0 50978 800
rect 51510 0 51622 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54086 0 54198 800
rect 54730 0 54842 800
rect 55374 0 55486 800
rect 56018 0 56130 800
rect 56662 0 56774 800
rect 57306 0 57418 800
rect 58594 0 58706 800
rect 59238 0 59350 800
rect 59882 0 59994 800
rect 60526 0 60638 800
rect 61170 0 61282 800
rect 61814 0 61926 800
rect 62458 0 62570 800
rect 63746 0 63858 800
rect 64390 0 64502 800
rect 65034 0 65146 800
rect 65678 0 65790 800
rect 66322 0 66434 800
rect 66966 0 67078 800
rect 67610 0 67722 800
rect 68898 0 69010 800
rect 69542 0 69654 800
rect 70186 0 70298 800
rect 70830 0 70942 800
rect 71474 0 71586 800
rect 72118 0 72230 800
rect 72762 0 72874 800
rect 73406 0 73518 800
rect 74694 0 74806 800
rect 75338 0 75450 800
<< obsm2 >>
rect 204 75144 578 75585
rect 802 75144 1866 75585
rect 2090 75144 2510 75585
rect 2734 75144 3154 75585
rect 3378 75144 3798 75585
rect 4022 75144 4442 75585
rect 4666 75144 5086 75585
rect 5310 75144 5730 75585
rect 5954 75144 6374 75585
rect 6598 75144 7662 75585
rect 7886 75144 8306 75585
rect 8530 75144 8950 75585
rect 9174 75144 9594 75585
rect 9818 75144 10238 75585
rect 10462 75144 10882 75585
rect 11106 75144 11526 75585
rect 11750 75144 12814 75585
rect 13038 75144 13458 75585
rect 13682 75144 14102 75585
rect 14326 75144 14746 75585
rect 14970 75144 15390 75585
rect 15614 75144 16034 75585
rect 16258 75144 16678 75585
rect 16902 75144 17966 75585
rect 18190 75144 18610 75585
rect 18834 75144 19254 75585
rect 19478 75144 19898 75585
rect 20122 75144 20542 75585
rect 20766 75144 21186 75585
rect 21410 75144 21830 75585
rect 22054 75144 23118 75585
rect 23342 75144 23762 75585
rect 23986 75144 24406 75585
rect 24630 75144 25050 75585
rect 25274 75144 25694 75585
rect 25918 75144 26338 75585
rect 26562 75144 26982 75585
rect 27206 75144 27626 75585
rect 27850 75144 28914 75585
rect 29138 75144 29558 75585
rect 29782 75144 30202 75585
rect 30426 75144 30846 75585
rect 31070 75144 31490 75585
rect 31714 75144 32134 75585
rect 32358 75144 32778 75585
rect 33002 75144 34066 75585
rect 34290 75144 34710 75585
rect 34934 75144 35354 75585
rect 35578 75144 35998 75585
rect 36222 75144 36642 75585
rect 36866 75144 37286 75585
rect 37510 75144 37930 75585
rect 38154 75144 39218 75585
rect 39442 75144 39862 75585
rect 40086 75144 40506 75585
rect 40730 75144 41150 75585
rect 41374 75144 41794 75585
rect 42018 75144 42438 75585
rect 42662 75144 43082 75585
rect 43306 75144 44370 75585
rect 44594 75144 45014 75585
rect 45238 75144 45658 75585
rect 45882 75144 46302 75585
rect 46526 75144 46946 75585
rect 47170 75144 47590 75585
rect 47814 75144 48234 75585
rect 48458 75144 49522 75585
rect 49746 75144 50166 75585
rect 50390 75144 50810 75585
rect 51034 75144 51454 75585
rect 51678 75144 52098 75585
rect 52322 75144 52742 75585
rect 52966 75144 53386 75585
rect 53610 75144 54030 75585
rect 54254 75144 55318 75585
rect 55542 75144 55962 75585
rect 56186 75144 56606 75585
rect 56830 75144 57250 75585
rect 57474 75144 57894 75585
rect 58118 75144 58538 75585
rect 58762 75144 59182 75585
rect 59406 75144 60470 75585
rect 60694 75144 61114 75585
rect 61338 75144 61758 75585
rect 61982 75144 62402 75585
rect 62626 75144 63046 75585
rect 63270 75144 63690 75585
rect 63914 75144 64334 75585
rect 64558 75144 65622 75585
rect 65846 75144 66266 75585
rect 66490 75144 66910 75585
rect 67134 75144 67554 75585
rect 67778 75144 68198 75585
rect 68422 75144 68842 75585
rect 69066 75144 69486 75585
rect 69710 75144 70774 75585
rect 70998 75144 71418 75585
rect 71642 75144 72062 75585
rect 72286 75144 72706 75585
rect 72930 75144 73350 75585
rect 73574 75144 73994 75585
rect 74218 75144 74638 75585
rect 74862 75144 75420 75585
rect 204 856 75420 75144
rect 204 31 578 856
rect 802 31 1222 856
rect 1446 31 1866 856
rect 2090 31 2510 856
rect 2734 31 3154 856
rect 3378 31 3798 856
rect 4022 31 4442 856
rect 4666 31 5730 856
rect 5954 31 6374 856
rect 6598 31 7018 856
rect 7242 31 7662 856
rect 7886 31 8306 856
rect 8530 31 8950 856
rect 9174 31 9594 856
rect 9818 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12170 856
rect 12394 31 12814 856
rect 13038 31 13458 856
rect 13682 31 14102 856
rect 14326 31 14746 856
rect 14970 31 16034 856
rect 16258 31 16678 856
rect 16902 31 17322 856
rect 17546 31 17966 856
rect 18190 31 18610 856
rect 18834 31 19254 856
rect 19478 31 19898 856
rect 20122 31 21186 856
rect 21410 31 21830 856
rect 22054 31 22474 856
rect 22698 31 23118 856
rect 23342 31 23762 856
rect 23986 31 24406 856
rect 24630 31 25050 856
rect 25274 31 25694 856
rect 25918 31 26982 856
rect 27206 31 27626 856
rect 27850 31 28270 856
rect 28494 31 28914 856
rect 29138 31 29558 856
rect 29782 31 30202 856
rect 30426 31 30846 856
rect 31070 31 32134 856
rect 32358 31 32778 856
rect 33002 31 33422 856
rect 33646 31 34066 856
rect 34290 31 34710 856
rect 34934 31 35354 856
rect 35578 31 35998 856
rect 36222 31 37286 856
rect 37510 31 37930 856
rect 38154 31 38574 856
rect 38798 31 39218 856
rect 39442 31 39862 856
rect 40086 31 40506 856
rect 40730 31 41150 856
rect 41374 31 42438 856
rect 42662 31 43082 856
rect 43306 31 43726 856
rect 43950 31 44370 856
rect 44594 31 45014 856
rect 45238 31 45658 856
rect 45882 31 46302 856
rect 46526 31 47590 856
rect 47814 31 48234 856
rect 48458 31 48878 856
rect 49102 31 49522 856
rect 49746 31 50166 856
rect 50390 31 50810 856
rect 51034 31 51454 856
rect 51678 31 52098 856
rect 52322 31 53386 856
rect 53610 31 54030 856
rect 54254 31 54674 856
rect 54898 31 55318 856
rect 55542 31 55962 856
rect 56186 31 56606 856
rect 56830 31 57250 856
rect 57474 31 58538 856
rect 58762 31 59182 856
rect 59406 31 59826 856
rect 60050 31 60470 856
rect 60694 31 61114 856
rect 61338 31 61758 856
rect 61982 31 62402 856
rect 62626 31 63690 856
rect 63914 31 64334 856
rect 64558 31 64978 856
rect 65202 31 65622 856
rect 65846 31 66266 856
rect 66490 31 66910 856
rect 67134 31 67554 856
rect 67778 31 68842 856
rect 69066 31 69486 856
rect 69710 31 70130 856
rect 70354 31 70774 856
rect 70998 31 71418 856
rect 71642 31 72062 856
rect 72286 31 72706 856
rect 72930 31 73350 856
rect 73574 31 74638 856
rect 74862 31 75282 856
<< metal3 >>
rect 0 75428 800 75668
rect 75200 75428 76000 75668
rect 0 74748 800 74988
rect 75200 74748 76000 74988
rect 0 74068 800 74308
rect 75200 74068 76000 74308
rect 0 73388 800 73628
rect 75200 73388 76000 73628
rect 0 72708 800 72948
rect 75200 72708 76000 72948
rect 75200 72028 76000 72268
rect 0 71348 800 71588
rect 75200 71348 76000 71588
rect 0 70668 800 70908
rect 75200 70668 76000 70908
rect 0 69988 800 70228
rect 0 69308 800 69548
rect 75200 69308 76000 69548
rect 0 68628 800 68868
rect 75200 68628 76000 68868
rect 0 67948 800 68188
rect 75200 67948 76000 68188
rect 0 67268 800 67508
rect 75200 67268 76000 67508
rect 75200 66588 76000 66828
rect 0 65908 800 66148
rect 75200 65908 76000 66148
rect 0 65228 800 65468
rect 75200 65228 76000 65468
rect 0 64548 800 64788
rect 0 63868 800 64108
rect 75200 63868 76000 64108
rect 0 63188 800 63428
rect 75200 63188 76000 63428
rect 0 62508 800 62748
rect 75200 62508 76000 62748
rect 0 61828 800 62068
rect 75200 61828 76000 62068
rect 75200 61148 76000 61388
rect 0 60468 800 60708
rect 75200 60468 76000 60708
rect 0 59788 800 60028
rect 75200 59788 76000 60028
rect 0 59108 800 59348
rect 0 58428 800 58668
rect 75200 58428 76000 58668
rect 0 57748 800 57988
rect 75200 57748 76000 57988
rect 0 57068 800 57308
rect 75200 57068 76000 57308
rect 0 56388 800 56628
rect 75200 56388 76000 56628
rect 75200 55708 76000 55948
rect 0 55028 800 55268
rect 75200 55028 76000 55268
rect 0 54348 800 54588
rect 75200 54348 76000 54588
rect 0 53668 800 53908
rect 0 52988 800 53228
rect 75200 52988 76000 53228
rect 0 52308 800 52548
rect 75200 52308 76000 52548
rect 0 51628 800 51868
rect 75200 51628 76000 51868
rect 0 50948 800 51188
rect 75200 50948 76000 51188
rect 0 50268 800 50508
rect 75200 50268 76000 50508
rect 75200 49588 76000 49828
rect 0 48908 800 49148
rect 75200 48908 76000 49148
rect 0 48228 800 48468
rect 75200 48228 76000 48468
rect 0 47548 800 47788
rect 0 46868 800 47108
rect 75200 46868 76000 47108
rect 0 46188 800 46428
rect 75200 46188 76000 46428
rect 0 45508 800 45748
rect 75200 45508 76000 45748
rect 0 44828 800 45068
rect 75200 44828 76000 45068
rect 75200 44148 76000 44388
rect 0 43468 800 43708
rect 75200 43468 76000 43708
rect 0 42788 800 43028
rect 75200 42788 76000 43028
rect 0 42108 800 42348
rect 0 41428 800 41668
rect 75200 41428 76000 41668
rect 0 40748 800 40988
rect 75200 40748 76000 40988
rect 0 40068 800 40308
rect 75200 40068 76000 40308
rect 0 39388 800 39628
rect 75200 39388 76000 39628
rect 75200 38708 76000 38948
rect 0 38028 800 38268
rect 75200 38028 76000 38268
rect 0 37348 800 37588
rect 75200 37348 76000 37588
rect 0 36668 800 36908
rect 0 35988 800 36228
rect 75200 35988 76000 36228
rect 0 35308 800 35548
rect 75200 35308 76000 35548
rect 0 34628 800 34868
rect 75200 34628 76000 34868
rect 0 33948 800 34188
rect 75200 33948 76000 34188
rect 75200 33268 76000 33508
rect 0 32588 800 32828
rect 75200 32588 76000 32828
rect 0 31908 800 32148
rect 75200 31908 76000 32148
rect 0 31228 800 31468
rect 0 30548 800 30788
rect 75200 30548 76000 30788
rect 0 29868 800 30108
rect 75200 29868 76000 30108
rect 0 29188 800 29428
rect 75200 29188 76000 29428
rect 0 28508 800 28748
rect 75200 28508 76000 28748
rect 75200 27828 76000 28068
rect 0 27148 800 27388
rect 75200 27148 76000 27388
rect 0 26468 800 26708
rect 75200 26468 76000 26708
rect 0 25788 800 26028
rect 0 25108 800 25348
rect 75200 25108 76000 25348
rect 0 24428 800 24668
rect 75200 24428 76000 24668
rect 0 23748 800 23988
rect 75200 23748 76000 23988
rect 0 23068 800 23308
rect 75200 23068 76000 23308
rect 0 22388 800 22628
rect 75200 22388 76000 22628
rect 75200 21708 76000 21948
rect 0 21028 800 21268
rect 75200 21028 76000 21268
rect 0 20348 800 20588
rect 75200 20348 76000 20588
rect 0 19668 800 19908
rect 0 18988 800 19228
rect 75200 18988 76000 19228
rect 0 18308 800 18548
rect 75200 18308 76000 18548
rect 0 17628 800 17868
rect 75200 17628 76000 17868
rect 0 16948 800 17188
rect 75200 16948 76000 17188
rect 75200 16268 76000 16508
rect 0 15588 800 15828
rect 75200 15588 76000 15828
rect 0 14908 800 15148
rect 75200 14908 76000 15148
rect 0 14228 800 14468
rect 0 13548 800 13788
rect 75200 13548 76000 13788
rect 0 12868 800 13108
rect 75200 12868 76000 13108
rect 0 12188 800 12428
rect 75200 12188 76000 12428
rect 0 11508 800 11748
rect 75200 11508 76000 11748
rect 75200 10828 76000 11068
rect 0 10148 800 10388
rect 75200 10148 76000 10388
rect 0 9468 800 9708
rect 75200 9468 76000 9708
rect 0 8788 800 9028
rect 0 8108 800 8348
rect 75200 8108 76000 8348
rect 0 7428 800 7668
rect 75200 7428 76000 7668
rect 0 6748 800 6988
rect 75200 6748 76000 6988
rect 0 6068 800 6308
rect 75200 6068 76000 6308
rect 75200 5388 76000 5628
rect 0 4708 800 4948
rect 75200 4708 76000 4948
rect 0 4028 800 4268
rect 75200 4028 76000 4268
rect 0 3348 800 3588
rect 0 2668 800 2908
rect 75200 2668 76000 2908
rect 0 1988 800 2228
rect 75200 1988 76000 2228
rect 0 1308 800 1548
rect 75200 1308 76000 1548
rect 0 628 800 868
rect 75200 628 76000 868
rect 75200 -52 76000 188
<< obsm3 >>
rect 880 75348 75120 75581
rect 800 75068 75200 75348
rect 880 74668 75120 75068
rect 800 74388 75200 74668
rect 880 73988 75120 74388
rect 800 73708 75200 73988
rect 880 73308 75120 73708
rect 800 73028 75200 73308
rect 880 72628 75120 73028
rect 800 72348 75200 72628
rect 800 71948 75120 72348
rect 800 71668 75200 71948
rect 880 71268 75120 71668
rect 800 70988 75200 71268
rect 880 70588 75120 70988
rect 800 70308 75200 70588
rect 880 69908 75200 70308
rect 800 69628 75200 69908
rect 880 69228 75120 69628
rect 800 68948 75200 69228
rect 880 68548 75120 68948
rect 800 68268 75200 68548
rect 880 67868 75120 68268
rect 800 67588 75200 67868
rect 880 67188 75120 67588
rect 800 66908 75200 67188
rect 800 66508 75120 66908
rect 800 66228 75200 66508
rect 880 65828 75120 66228
rect 800 65548 75200 65828
rect 880 65148 75120 65548
rect 800 64868 75200 65148
rect 880 64468 75200 64868
rect 800 64188 75200 64468
rect 880 63788 75120 64188
rect 800 63508 75200 63788
rect 880 63108 75120 63508
rect 800 62828 75200 63108
rect 880 62428 75120 62828
rect 800 62148 75200 62428
rect 880 61748 75120 62148
rect 800 61468 75200 61748
rect 800 61068 75120 61468
rect 800 60788 75200 61068
rect 880 60388 75120 60788
rect 800 60108 75200 60388
rect 880 59708 75120 60108
rect 800 59428 75200 59708
rect 880 59028 75200 59428
rect 800 58748 75200 59028
rect 880 58348 75120 58748
rect 800 58068 75200 58348
rect 880 57668 75120 58068
rect 800 57388 75200 57668
rect 880 56988 75120 57388
rect 800 56708 75200 56988
rect 880 56308 75120 56708
rect 800 56028 75200 56308
rect 800 55628 75120 56028
rect 800 55348 75200 55628
rect 880 54948 75120 55348
rect 800 54668 75200 54948
rect 880 54268 75120 54668
rect 800 53988 75200 54268
rect 880 53588 75200 53988
rect 800 53308 75200 53588
rect 880 52908 75120 53308
rect 800 52628 75200 52908
rect 880 52228 75120 52628
rect 800 51948 75200 52228
rect 880 51548 75120 51948
rect 800 51268 75200 51548
rect 880 50868 75120 51268
rect 800 50588 75200 50868
rect 880 50188 75120 50588
rect 800 49908 75200 50188
rect 800 49508 75120 49908
rect 800 49228 75200 49508
rect 880 48828 75120 49228
rect 800 48548 75200 48828
rect 880 48148 75120 48548
rect 800 47868 75200 48148
rect 880 47468 75200 47868
rect 800 47188 75200 47468
rect 880 46788 75120 47188
rect 800 46508 75200 46788
rect 880 46108 75120 46508
rect 800 45828 75200 46108
rect 880 45428 75120 45828
rect 800 45148 75200 45428
rect 880 44748 75120 45148
rect 800 44468 75200 44748
rect 800 44068 75120 44468
rect 800 43788 75200 44068
rect 880 43388 75120 43788
rect 800 43108 75200 43388
rect 880 42708 75120 43108
rect 800 42428 75200 42708
rect 880 42028 75200 42428
rect 800 41748 75200 42028
rect 880 41348 75120 41748
rect 800 41068 75200 41348
rect 880 40668 75120 41068
rect 800 40388 75200 40668
rect 880 39988 75120 40388
rect 800 39708 75200 39988
rect 880 39308 75120 39708
rect 800 39028 75200 39308
rect 800 38628 75120 39028
rect 800 38348 75200 38628
rect 880 37948 75120 38348
rect 800 37668 75200 37948
rect 880 37268 75120 37668
rect 800 36988 75200 37268
rect 880 36588 75200 36988
rect 800 36308 75200 36588
rect 880 35908 75120 36308
rect 800 35628 75200 35908
rect 880 35228 75120 35628
rect 800 34948 75200 35228
rect 880 34548 75120 34948
rect 800 34268 75200 34548
rect 880 33868 75120 34268
rect 800 33588 75200 33868
rect 800 33188 75120 33588
rect 800 32908 75200 33188
rect 880 32508 75120 32908
rect 800 32228 75200 32508
rect 880 31828 75120 32228
rect 800 31548 75200 31828
rect 880 31148 75200 31548
rect 800 30868 75200 31148
rect 880 30468 75120 30868
rect 800 30188 75200 30468
rect 880 29788 75120 30188
rect 800 29508 75200 29788
rect 880 29108 75120 29508
rect 800 28828 75200 29108
rect 880 28428 75120 28828
rect 800 28148 75200 28428
rect 800 27748 75120 28148
rect 800 27468 75200 27748
rect 880 27068 75120 27468
rect 800 26788 75200 27068
rect 880 26388 75120 26788
rect 800 26108 75200 26388
rect 880 25708 75200 26108
rect 800 25428 75200 25708
rect 880 25028 75120 25428
rect 800 24748 75200 25028
rect 880 24348 75120 24748
rect 800 24068 75200 24348
rect 880 23668 75120 24068
rect 800 23388 75200 23668
rect 880 22988 75120 23388
rect 800 22708 75200 22988
rect 880 22308 75120 22708
rect 800 22028 75200 22308
rect 800 21628 75120 22028
rect 800 21348 75200 21628
rect 880 20948 75120 21348
rect 800 20668 75200 20948
rect 880 20268 75120 20668
rect 800 19988 75200 20268
rect 880 19588 75200 19988
rect 800 19308 75200 19588
rect 880 18908 75120 19308
rect 800 18628 75200 18908
rect 880 18228 75120 18628
rect 800 17948 75200 18228
rect 880 17548 75120 17948
rect 800 17268 75200 17548
rect 880 16868 75120 17268
rect 800 16588 75200 16868
rect 800 16188 75120 16588
rect 800 15908 75200 16188
rect 880 15508 75120 15908
rect 800 15228 75200 15508
rect 880 14828 75120 15228
rect 800 14548 75200 14828
rect 880 14148 75200 14548
rect 800 13868 75200 14148
rect 880 13468 75120 13868
rect 800 13188 75200 13468
rect 880 12788 75120 13188
rect 800 12508 75200 12788
rect 880 12108 75120 12508
rect 800 11828 75200 12108
rect 880 11428 75120 11828
rect 800 11148 75200 11428
rect 800 10748 75120 11148
rect 800 10468 75200 10748
rect 880 10068 75120 10468
rect 800 9788 75200 10068
rect 880 9388 75120 9788
rect 800 9108 75200 9388
rect 880 8708 75200 9108
rect 800 8428 75200 8708
rect 880 8028 75120 8428
rect 800 7748 75200 8028
rect 880 7348 75120 7748
rect 800 7068 75200 7348
rect 880 6668 75120 7068
rect 800 6388 75200 6668
rect 880 5988 75120 6388
rect 800 5708 75200 5988
rect 800 5308 75120 5708
rect 800 5028 75200 5308
rect 880 4628 75120 5028
rect 800 4348 75200 4628
rect 880 3948 75120 4348
rect 800 3668 75200 3948
rect 880 3268 75200 3668
rect 800 2988 75200 3268
rect 880 2588 75120 2988
rect 800 2308 75200 2588
rect 880 1908 75120 2308
rect 800 1628 75200 1908
rect 880 1228 75120 1628
rect 800 948 75200 1228
rect 880 548 75120 948
rect 800 268 75200 548
rect 800 35 75120 268
<< metal4 >>
rect 4208 2128 4528 73488
rect 19568 2128 19888 73488
rect 34928 2128 35248 73488
rect 50288 2128 50608 73488
rect 65648 2128 65968 73488
<< labels >>
rlabel metal3 s 75200 20348 76000 20588 6 active
port 1 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 74694 0 74806 800 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 75200 60468 76000 60708 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 75200 70668 76000 70908 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 75200 40068 76000 40308 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 75200 67948 76000 68188 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 68628 800 68868 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 39918 75200 40030 76000 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 42494 75200 42606 76000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 58594 75200 58706 76000 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 0 54348 800 54588 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 67610 75200 67722 76000 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 0 75428 800 75668 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 52154 0 52266 800 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 75200 74068 76000 74308 6 io_in[28]
port 22 nsew signal input
rlabel metal3 s 75200 51628 76000 51868 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 48934 0 49046 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 0 56388 800 56628 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 44426 75200 44538 76000 6 io_in[33]
port 28 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 75200 27148 76000 27388 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 60526 75200 60638 76000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 14802 75200 14914 76000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 46358 75200 46470 76000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 47002 75200 47114 76000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 5142 75200 5254 76000 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 75200 8108 76000 8348 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 74068 800 74308 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 66966 0 67078 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 75200 16948 76000 17188 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 0 25108 800 25348 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 75200 52308 76000 52548 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal2 s 50222 75200 50334 76000 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 73388 800 73628 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 24462 75200 24574 76000 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal2 s 59882 0 59994 800 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal3 s 75200 61828 76000 62068 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 10294 75200 10406 76000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 0 52308 800 52548 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 0 70668 800 70908 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 75200 10148 76000 10388 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 35410 0 35522 800 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 634 75200 746 76000 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal3 s 75200 1988 76000 2228 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal3 s 0 74748 800 74988 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 0 47548 800 47788 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal3 s 75200 27828 76000 28068 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 0 36668 800 36908 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 45714 0 45826 800 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal2 s 66322 75200 66434 76000 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal3 s 75200 29188 76000 29428 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 70186 0 70298 800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 45070 75200 45182 76000 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 0 53668 800 53908 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 43138 75200 43250 76000 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 27148 800 27388 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 75200 68628 76000 68868 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal2 s 13514 75200 13626 76000 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal3 s 75200 -52 76000 188 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 0 69988 800 70228 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 65228 800 65468 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 0 35308 800 35548 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 30902 75200 31014 76000 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 61814 0 61926 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal2 s 74050 75200 74162 76000 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 75200 52988 76000 53228 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal2 s 2566 75200 2678 76000 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal2 s 48290 75200 48402 76000 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal3 s 0 52988 800 53228 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 0 62508 800 62748 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 75200 72708 76000 72948 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 10938 75200 11050 76000 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 39274 75200 39386 76000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal3 s 75200 38708 76000 38948 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 15588 800 15828 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal3 s 75200 4028 76000 4268 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 0 41428 800 41668 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 71474 0 71586 800 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 75200 66588 76000 66828 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 75200 22388 76000 22628 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 34122 0 34234 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 3854 75200 3966 76000 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal2 s 37986 75200 38098 76000 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 75200 55028 76000 55268 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal2 s 56018 75200 56130 76000 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 48908 800 49148 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal2 s 68898 0 69010 800 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal2 s 25750 0 25862 800 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal2 s 19954 75200 20066 76000 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 34766 75200 34878 76000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal2 s 72118 75200 72230 76000 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 27038 75200 27150 76000 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal2 s 1922 75200 2034 76000 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 15446 75200 15558 76000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 0 35988 800 36228 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 75200 12868 76000 13108 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 5786 75200 5898 76000 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 75200 7428 76000 7668 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal2 s 41850 75200 41962 76000 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 3210 75200 3322 76000 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 19310 75200 19422 76000 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 75200 12188 76000 12428 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 43138 0 43250 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal2 s 61170 0 61282 800 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 75200 16268 76000 16508 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 75200 11508 76000 11748 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 75200 28508 76000 28748 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 64390 75200 64502 76000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 68254 75200 68366 76000 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 75200 71348 76000 71588 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 75200 63188 76000 63428 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 66322 0 66434 800 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal2 s 51510 75200 51622 76000 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 57306 75200 57418 76000 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal2 s 62458 75200 62570 76000 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 73406 75200 73518 76000 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 75200 74748 76000 74988 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 75200 50948 76000 51188 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 54086 75200 54198 76000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal2 s 50222 0 50334 800 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal2 s 14158 75200 14270 76000 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 54086 0 54198 800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 34122 75200 34234 76000 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal2 s 32834 0 32946 800 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal3 s 75200 46188 76000 46428 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal3 s 75200 15588 76000 15828 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal3 s 0 21028 800 21268 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal2 s 47646 0 47758 800 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 0 63188 800 63428 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal2 s 30258 0 30370 800 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal2 s 12226 0 12338 800 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 75200 30548 76000 30788 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 32588 800 32828 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal3 s 0 69308 800 69548 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 21242 75200 21354 76000 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal3 s 0 72708 800 72948 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 75200 61148 76000 61388 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal2 s 70830 75200 70942 76000 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 75200 33268 76000 33508 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal2 s 45714 75200 45826 76000 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal3 s 0 40748 800 40988 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 75200 26468 76000 26708 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 0 30548 800 30788 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal2 s 18666 75200 18778 76000 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 41206 75200 41318 76000 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal3 s 75200 57068 76000 57308 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal2 s 32190 75200 32302 76000 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal3 s 75200 65908 76000 66148 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal3 s 75200 5388 76000 5628 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal2 s 63102 75200 63214 76000 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 0 1308 800 1548 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s 16734 75200 16846 76000 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal2 s 7718 75200 7830 76000 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 9006 75200 9118 76000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 60468 800 60708 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 29614 75200 29726 76000 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 0 59788 800 60028 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 75200 9468 76000 9708 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 34766 0 34878 800 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 75200 56388 76000 56628 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 75200 25108 76000 25348 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal2 s 72762 0 72874 800 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal2 s 30258 75200 30370 76000 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 56662 75200 56774 76000 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 0 3348 800 3588 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 55028 800 55268 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal2 s 37342 75200 37454 76000 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 3854 0 3966 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal2 s 65678 0 65790 800 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 0 57068 800 57308 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal2 s 65034 0 65146 800 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 75200 34628 76000 34868 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal2 s 16090 75200 16202 76000 6 la2_data_in[0]
port 212 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la2_data_in[10]
port 213 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la2_data_in[11]
port 214 nsew signal input
rlabel metal3 s 0 65908 800 66148 6 la2_data_in[12]
port 215 nsew signal input
rlabel metal2 s 23174 75200 23286 76000 6 la2_data_in[13]
port 216 nsew signal input
rlabel metal2 s 36054 75200 36166 76000 6 la2_data_in[14]
port 217 nsew signal input
rlabel metal3 s 75200 13548 76000 13788 6 la2_data_in[15]
port 218 nsew signal input
rlabel metal2 s 61814 75200 61926 76000 6 la2_data_in[16]
port 219 nsew signal input
rlabel metal3 s 75200 48908 76000 49148 6 la2_data_in[17]
port 220 nsew signal input
rlabel metal3 s 75200 63868 76000 64108 6 la2_data_in[18]
port 221 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la2_data_in[19]
port 222 nsew signal input
rlabel metal2 s 26394 75200 26506 76000 6 la2_data_in[1]
port 223 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 la2_data_in[20]
port 224 nsew signal input
rlabel metal2 s 62458 0 62570 800 6 la2_data_in[21]
port 225 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la2_data_in[22]
port 226 nsew signal input
rlabel metal3 s 75200 17628 76000 17868 6 la2_data_in[23]
port 227 nsew signal input
rlabel metal3 s 75200 75428 76000 75668 6 la2_data_in[24]
port 228 nsew signal input
rlabel metal2 s 45070 0 45182 800 6 la2_data_in[25]
port 229 nsew signal input
rlabel metal3 s 75200 32588 76000 32828 6 la2_data_in[26]
port 230 nsew signal input
rlabel metal3 s 75200 24428 76000 24668 6 la2_data_in[27]
port 231 nsew signal input
rlabel metal3 s 75200 50268 76000 50508 6 la2_data_in[28]
port 232 nsew signal input
rlabel metal3 s 75200 39388 76000 39628 6 la2_data_in[29]
port 233 nsew signal input
rlabel metal2 s 32834 75200 32946 76000 6 la2_data_in[2]
port 234 nsew signal input
rlabel metal3 s 75200 40748 76000 40988 6 la2_data_in[30]
port 235 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la2_data_in[31]
port 236 nsew signal input
rlabel metal2 s 63746 0 63858 800 6 la2_data_in[3]
port 237 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la2_data_in[4]
port 238 nsew signal input
rlabel metal3 s 0 50268 800 50508 6 la2_data_in[5]
port 239 nsew signal input
rlabel metal2 s 57306 0 57418 800 6 la2_data_in[6]
port 240 nsew signal input
rlabel metal3 s 75200 2668 76000 2908 6 la2_data_in[7]
port 241 nsew signal input
rlabel metal2 s 12870 75200 12982 76000 6 la2_data_in[8]
port 242 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 la2_data_in[9]
port 243 nsew signal input
rlabel metal2 s 35410 75200 35522 76000 6 la2_data_out[0]
port 244 nsew signal bidirectional
rlabel metal3 s 0 59108 800 59348 6 la2_data_out[10]
port 245 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la2_data_out[11]
port 246 nsew signal bidirectional
rlabel metal3 s 75200 43468 76000 43708 6 la2_data_out[12]
port 247 nsew signal bidirectional
rlabel metal2 s 64390 0 64502 800 6 la2_data_out[13]
port 248 nsew signal bidirectional
rlabel metal3 s 0 23068 800 23308 6 la2_data_out[14]
port 249 nsew signal bidirectional
rlabel metal2 s 12870 0 12982 800 6 la2_data_out[15]
port 250 nsew signal bidirectional
rlabel metal3 s 75200 37348 76000 37588 6 la2_data_out[16]
port 251 nsew signal bidirectional
rlabel metal3 s 0 26468 800 26708 6 la2_data_out[17]
port 252 nsew signal bidirectional
rlabel metal3 s 75200 73388 76000 73628 6 la2_data_out[18]
port 253 nsew signal bidirectional
rlabel metal3 s 75200 62508 76000 62748 6 la2_data_out[19]
port 254 nsew signal bidirectional
rlabel metal3 s 75200 59788 76000 60028 6 la2_data_out[1]
port 255 nsew signal bidirectional
rlabel metal3 s 75200 58428 76000 58668 6 la2_data_out[20]
port 256 nsew signal bidirectional
rlabel metal2 s 37342 0 37454 800 6 la2_data_out[21]
port 257 nsew signal bidirectional
rlabel metal2 s 69542 75200 69654 76000 6 la2_data_out[22]
port 258 nsew signal bidirectional
rlabel metal2 s 1922 0 2034 800 6 la2_data_out[23]
port 259 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la2_data_out[24]
port 260 nsew signal bidirectional
rlabel metal2 s 4498 75200 4610 76000 6 la2_data_out[25]
port 261 nsew signal bidirectional
rlabel metal2 s 37986 0 38098 800 6 la2_data_out[26]
port 262 nsew signal bidirectional
rlabel metal2 s 75338 0 75450 800 6 la2_data_out[27]
port 263 nsew signal bidirectional
rlabel metal2 s 74694 75200 74806 76000 6 la2_data_out[28]
port 264 nsew signal bidirectional
rlabel metal3 s 75200 6068 76000 6308 6 la2_data_out[29]
port 265 nsew signal bidirectional
rlabel metal2 s 31546 75200 31658 76000 6 la2_data_out[2]
port 266 nsew signal bidirectional
rlabel metal3 s 0 50948 800 51188 6 la2_data_out[30]
port 267 nsew signal bidirectional
rlabel metal2 s 13514 0 13626 800 6 la2_data_out[31]
port 268 nsew signal bidirectional
rlabel metal2 s 32190 0 32302 800 6 la2_data_out[3]
port 269 nsew signal bidirectional
rlabel metal2 s 65678 75200 65790 76000 6 la2_data_out[4]
port 270 nsew signal bidirectional
rlabel metal3 s 0 20348 800 20588 6 la2_data_out[5]
port 271 nsew signal bidirectional
rlabel metal2 s 27682 0 27794 800 6 la2_data_out[6]
port 272 nsew signal bidirectional
rlabel metal3 s 0 58428 800 58668 6 la2_data_out[7]
port 273 nsew signal bidirectional
rlabel metal3 s 75200 33948 76000 34188 6 la2_data_out[8]
port 274 nsew signal bidirectional
rlabel metal3 s 75200 48228 76000 48468 6 la2_data_out[9]
port 275 nsew signal bidirectional
rlabel metal2 s 56018 0 56130 800 6 la2_oenb[0]
port 276 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la2_oenb[10]
port 277 nsew signal input
rlabel metal2 s 72118 0 72230 800 6 la2_oenb[11]
port 278 nsew signal input
rlabel metal3 s 75200 45508 76000 45748 6 la2_oenb[12]
port 279 nsew signal input
rlabel metal2 s 53442 75200 53554 76000 6 la2_oenb[13]
port 280 nsew signal input
rlabel metal3 s 0 628 800 868 6 la2_oenb[14]
port 281 nsew signal input
rlabel metal2 s 55374 0 55486 800 6 la2_oenb[15]
port 282 nsew signal input
rlabel metal2 s 68898 75200 69010 76000 6 la2_oenb[16]
port 283 nsew signal input
rlabel metal3 s 75200 4708 76000 4948 6 la2_oenb[17]
port 284 nsew signal input
rlabel metal2 s 47646 75200 47758 76000 6 la2_oenb[18]
port 285 nsew signal input
rlabel metal2 s 67610 0 67722 800 6 la2_oenb[19]
port 286 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 la2_oenb[1]
port 287 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la2_oenb[20]
port 288 nsew signal input
rlabel metal3 s 75200 35308 76000 35548 6 la2_oenb[21]
port 289 nsew signal input
rlabel metal2 s -10 75200 102 76000 6 la2_oenb[22]
port 290 nsew signal input
rlabel metal3 s 75200 46868 76000 47108 6 la2_oenb[23]
port 291 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la2_oenb[24]
port 292 nsew signal input
rlabel metal2 s 69542 0 69654 800 6 la2_oenb[25]
port 293 nsew signal input
rlabel metal2 s 25106 75200 25218 76000 6 la2_oenb[26]
port 294 nsew signal input
rlabel metal2 s 66966 75200 67078 76000 6 la2_oenb[27]
port 295 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la2_oenb[28]
port 296 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la2_oenb[29]
port 297 nsew signal input
rlabel metal2 s 28970 75200 29082 76000 6 la2_oenb[2]
port 298 nsew signal input
rlabel metal3 s 75200 10828 76000 11068 6 la2_oenb[30]
port 299 nsew signal input
rlabel metal2 s 18022 75200 18134 76000 6 la2_oenb[31]
port 300 nsew signal input
rlabel metal3 s 75200 23748 76000 23988 6 la2_oenb[3]
port 301 nsew signal input
rlabel metal2 s 52154 75200 52266 76000 6 la2_oenb[4]
port 302 nsew signal input
rlabel metal2 s 36698 75200 36810 76000 6 la2_oenb[5]
port 303 nsew signal input
rlabel metal2 s 8362 75200 8474 76000 6 la2_oenb[6]
port 304 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la2_oenb[7]
port 305 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la2_oenb[8]
port 306 nsew signal input
rlabel metal3 s 75200 54348 76000 54588 6 la2_oenb[9]
port 307 nsew signal input
rlabel metal3 s 75200 49588 76000 49828 6 la3_data_in[0]
port 308 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 la3_data_in[10]
port 309 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la3_data_in[11]
port 310 nsew signal input
rlabel metal3 s 75200 21708 76000 21948 6 la3_data_in[12]
port 311 nsew signal input
rlabel metal2 s 70830 0 70942 800 6 la3_data_in[13]
port 312 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_data_in[14]
port 313 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la3_data_in[15]
port 314 nsew signal input
rlabel metal2 s 41206 0 41318 800 6 la3_data_in[16]
port 315 nsew signal input
rlabel metal2 s 59238 0 59350 800 6 la3_data_in[17]
port 316 nsew signal input
rlabel metal3 s 75200 14908 76000 15148 6 la3_data_in[18]
port 317 nsew signal input
rlabel metal2 s 11582 75200 11694 76000 6 la3_data_in[19]
port 318 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 la3_data_in[1]
port 319 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la3_data_in[20]
port 320 nsew signal input
rlabel metal2 s 27682 75200 27794 76000 6 la3_data_in[21]
port 321 nsew signal input
rlabel metal3 s 75200 42788 76000 43028 6 la3_data_in[22]
port 322 nsew signal input
rlabel metal3 s 75200 72028 76000 72268 6 la3_data_in[23]
port 323 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la3_data_in[24]
port 324 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la3_data_in[25]
port 325 nsew signal input
rlabel metal3 s 75200 29868 76000 30108 6 la3_data_in[26]
port 326 nsew signal input
rlabel metal2 s 56662 0 56774 800 6 la3_data_in[27]
port 327 nsew signal input
rlabel metal2 s 59238 75200 59350 76000 6 la3_data_in[28]
port 328 nsew signal input
rlabel metal2 s 54730 0 54842 800 6 la3_data_in[29]
port 329 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la3_data_in[2]
port 330 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_data_in[30]
port 331 nsew signal input
rlabel metal2 s 73406 0 73518 800 6 la3_data_in[31]
port 332 nsew signal input
rlabel metal3 s 75200 18308 76000 18548 6 la3_data_in[3]
port 333 nsew signal input
rlabel metal2 s 25750 75200 25862 76000 6 la3_data_in[4]
port 334 nsew signal input
rlabel metal3 s 75200 65228 76000 65468 6 la3_data_in[5]
port 335 nsew signal input
rlabel metal3 s 0 61828 800 62068 6 la3_data_in[6]
port 336 nsew signal input
rlabel metal3 s 0 67268 800 67508 6 la3_data_in[7]
port 337 nsew signal input
rlabel metal3 s 0 64548 800 64788 6 la3_data_in[8]
port 338 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la3_data_in[9]
port 339 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_out[0]
port 340 nsew signal bidirectional
rlabel metal3 s 75200 38028 76000 38268 6 la3_data_out[10]
port 341 nsew signal bidirectional
rlabel metal2 s 42494 0 42606 800 6 la3_data_out[11]
port 342 nsew signal bidirectional
rlabel metal3 s 0 12868 800 13108 6 la3_data_out[12]
port 343 nsew signal bidirectional
rlabel metal2 s 71474 75200 71586 76000 6 la3_data_out[13]
port 344 nsew signal bidirectional
rlabel metal2 s 6430 75200 6542 76000 6 la3_data_out[14]
port 345 nsew signal bidirectional
rlabel metal3 s 0 33948 800 34188 6 la3_data_out[15]
port 346 nsew signal bidirectional
rlabel metal3 s 75200 44148 76000 44388 6 la3_data_out[16]
port 347 nsew signal bidirectional
rlabel metal2 s 72762 75200 72874 76000 6 la3_data_out[17]
port 348 nsew signal bidirectional
rlabel metal3 s 0 46868 800 47108 6 la3_data_out[18]
port 349 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la3_data_out[19]
port 350 nsew signal bidirectional
rlabel metal3 s 75200 23068 76000 23308 6 la3_data_out[1]
port 351 nsew signal bidirectional
rlabel metal2 s 50866 0 50978 800 6 la3_data_out[20]
port 352 nsew signal bidirectional
rlabel metal2 s 63746 75200 63858 76000 6 la3_data_out[21]
port 353 nsew signal bidirectional
rlabel metal2 s 20598 75200 20710 76000 6 la3_data_out[22]
port 354 nsew signal bidirectional
rlabel metal2 s 23174 0 23286 800 6 la3_data_out[23]
port 355 nsew signal bidirectional
rlabel metal3 s 75200 44828 76000 45068 6 la3_data_out[24]
port 356 nsew signal bidirectional
rlabel metal2 s 60526 0 60638 800 6 la3_data_out[25]
port 357 nsew signal bidirectional
rlabel metal3 s 75200 21028 76000 21268 6 la3_data_out[26]
port 358 nsew signal bidirectional
rlabel metal3 s 0 42108 800 42348 6 la3_data_out[27]
port 359 nsew signal bidirectional
rlabel metal3 s 75200 628 76000 868 6 la3_data_out[28]
port 360 nsew signal bidirectional
rlabel metal2 s 11582 0 11694 800 6 la3_data_out[29]
port 361 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 la3_data_out[2]
port 362 nsew signal bidirectional
rlabel metal3 s 75200 31908 76000 32148 6 la3_data_out[30]
port 363 nsew signal bidirectional
rlabel metal2 s 61170 75200 61282 76000 6 la3_data_out[31]
port 364 nsew signal bidirectional
rlabel metal3 s 75200 67268 76000 67508 6 la3_data_out[3]
port 365 nsew signal bidirectional
rlabel metal3 s 75200 1308 76000 1548 6 la3_data_out[4]
port 366 nsew signal bidirectional
rlabel metal2 s 5786 0 5898 800 6 la3_data_out[5]
port 367 nsew signal bidirectional
rlabel metal3 s 75200 41428 76000 41668 6 la3_data_out[6]
port 368 nsew signal bidirectional
rlabel metal2 s 1278 0 1390 800 6 la3_data_out[7]
port 369 nsew signal bidirectional
rlabel metal3 s 75200 69308 76000 69548 6 la3_data_out[8]
port 370 nsew signal bidirectional
rlabel metal2 s 57950 75200 58062 76000 6 la3_data_out[9]
port 371 nsew signal bidirectional
rlabel metal3 s 75200 6748 76000 6988 6 la3_oenb[0]
port 372 nsew signal input
rlabel metal2 s 55374 75200 55486 76000 6 la3_oenb[10]
port 373 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la3_oenb[11]
port 374 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 la3_oenb[12]
port 375 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 la3_oenb[13]
port 376 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 377 nsew signal input
rlabel metal2 s 58594 0 58706 800 6 la3_oenb[15]
port 378 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la3_oenb[16]
port 379 nsew signal input
rlabel metal3 s 0 67948 800 68188 6 la3_oenb[17]
port 380 nsew signal input
rlabel metal2 s 21886 75200 21998 76000 6 la3_oenb[18]
port 381 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 la3_oenb[19]
port 382 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 la3_oenb[1]
port 383 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_oenb[20]
port 384 nsew signal input
rlabel metal2 s 40562 75200 40674 76000 6 la3_oenb[21]
port 385 nsew signal input
rlabel metal2 s 23818 75200 23930 76000 6 la3_oenb[22]
port 386 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la3_oenb[23]
port 387 nsew signal input
rlabel metal2 s 52798 75200 52910 76000 6 la3_oenb[24]
port 388 nsew signal input
rlabel metal3 s 75200 18988 76000 19228 6 la3_oenb[25]
port 389 nsew signal input
rlabel metal3 s 0 51628 800 51868 6 la3_oenb[26]
port 390 nsew signal input
rlabel metal3 s 75200 57748 76000 57988 6 la3_oenb[27]
port 391 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la3_oenb[28]
port 392 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la3_oenb[29]
port 393 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la3_oenb[2]
port 394 nsew signal input
rlabel metal3 s 75200 55708 76000 55948 6 la3_oenb[30]
port 395 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 la3_oenb[31]
port 396 nsew signal input
rlabel metal2 s 50866 75200 50978 76000 6 la3_oenb[3]
port 397 nsew signal input
rlabel metal2 s 49578 75200 49690 76000 6 la3_oenb[4]
port 398 nsew signal input
rlabel metal3 s 0 71348 800 71588 6 la3_oenb[5]
port 399 nsew signal input
rlabel metal2 s 9650 75200 9762 76000 6 la3_oenb[6]
port 400 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 la3_oenb[7]
port 401 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la3_oenb[8]
port 402 nsew signal input
rlabel metal3 s 0 63868 800 64108 6 la3_oenb[9]
port 403 nsew signal input
rlabel metal4 s 4208 2128 4528 73488 6 vccd1
port 404 nsew power input
rlabel metal4 s 34928 2128 35248 73488 6 vccd1
port 404 nsew power input
rlabel metal4 s 65648 2128 65968 73488 6 vccd1
port 404 nsew power input
rlabel metal4 s 19568 2128 19888 73488 6 vssd1
port 405 nsew ground input
rlabel metal4 s 50288 2128 50608 73488 6 vssd1
port 405 nsew ground input
rlabel metal3 s 75200 35988 76000 36228 6 wb_clk_i
port 406 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 76000 76000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6551782
string GDS_FILE /openlane/designs/wrapped_instrumented_adder_sklansky/runs/RUN_2022.06.07_16.18.46/results/finishing/wrapped_instrumented_adder_sklansky.magic.gds
string GDS_START 685842
<< end >>

