magic
tech sky130A
magscale 1 2
timestamp 1654608992
<< obsli1 >>
rect 1104 2159 72864 71825
<< obsm1 >>
rect 198 1300 73494 72140
<< metal2 >>
rect -10 73200 102 74000
rect 634 73200 746 74000
rect 1278 73200 1390 74000
rect 2566 73200 2678 74000
rect 3210 73200 3322 74000
rect 3854 73200 3966 74000
rect 4498 73200 4610 74000
rect 5142 73200 5254 74000
rect 5786 73200 5898 74000
rect 6430 73200 6542 74000
rect 7074 73200 7186 74000
rect 7718 73200 7830 74000
rect 9006 73200 9118 74000
rect 9650 73200 9762 74000
rect 10294 73200 10406 74000
rect 10938 73200 11050 74000
rect 11582 73200 11694 74000
rect 12226 73200 12338 74000
rect 12870 73200 12982 74000
rect 13514 73200 13626 74000
rect 14158 73200 14270 74000
rect 15446 73200 15558 74000
rect 16090 73200 16202 74000
rect 16734 73200 16846 74000
rect 17378 73200 17490 74000
rect 18022 73200 18134 74000
rect 18666 73200 18778 74000
rect 19310 73200 19422 74000
rect 19954 73200 20066 74000
rect 20598 73200 20710 74000
rect 21886 73200 21998 74000
rect 22530 73200 22642 74000
rect 23174 73200 23286 74000
rect 23818 73200 23930 74000
rect 24462 73200 24574 74000
rect 25106 73200 25218 74000
rect 25750 73200 25862 74000
rect 26394 73200 26506 74000
rect 27038 73200 27150 74000
rect 28326 73200 28438 74000
rect 28970 73200 29082 74000
rect 29614 73200 29726 74000
rect 30258 73200 30370 74000
rect 30902 73200 31014 74000
rect 31546 73200 31658 74000
rect 32190 73200 32302 74000
rect 32834 73200 32946 74000
rect 33478 73200 33590 74000
rect 34766 73200 34878 74000
rect 35410 73200 35522 74000
rect 36054 73200 36166 74000
rect 36698 73200 36810 74000
rect 37342 73200 37454 74000
rect 37986 73200 38098 74000
rect 38630 73200 38742 74000
rect 39274 73200 39386 74000
rect 39918 73200 40030 74000
rect 40562 73200 40674 74000
rect 41850 73200 41962 74000
rect 42494 73200 42606 74000
rect 43138 73200 43250 74000
rect 43782 73200 43894 74000
rect 44426 73200 44538 74000
rect 45070 73200 45182 74000
rect 45714 73200 45826 74000
rect 46358 73200 46470 74000
rect 47002 73200 47114 74000
rect 48290 73200 48402 74000
rect 48934 73200 49046 74000
rect 49578 73200 49690 74000
rect 50222 73200 50334 74000
rect 50866 73200 50978 74000
rect 51510 73200 51622 74000
rect 52154 73200 52266 74000
rect 52798 73200 52910 74000
rect 53442 73200 53554 74000
rect 54730 73200 54842 74000
rect 55374 73200 55486 74000
rect 56018 73200 56130 74000
rect 56662 73200 56774 74000
rect 57306 73200 57418 74000
rect 57950 73200 58062 74000
rect 58594 73200 58706 74000
rect 59238 73200 59350 74000
rect 59882 73200 59994 74000
rect 61170 73200 61282 74000
rect 61814 73200 61926 74000
rect 62458 73200 62570 74000
rect 63102 73200 63214 74000
rect 63746 73200 63858 74000
rect 64390 73200 64502 74000
rect 65034 73200 65146 74000
rect 65678 73200 65790 74000
rect 66322 73200 66434 74000
rect 67610 73200 67722 74000
rect 68254 73200 68366 74000
rect 68898 73200 69010 74000
rect 69542 73200 69654 74000
rect 70186 73200 70298 74000
rect 70830 73200 70942 74000
rect 71474 73200 71586 74000
rect 72118 73200 72230 74000
rect 72762 73200 72874 74000
rect 73406 73200 73518 74000
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 41850 0 41962 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
rect 50222 0 50334 800
rect 50866 0 50978 800
rect 51510 0 51622 800
rect 52798 0 52910 800
rect 53442 0 53554 800
rect 54086 0 54198 800
rect 54730 0 54842 800
rect 55374 0 55486 800
rect 56018 0 56130 800
rect 56662 0 56774 800
rect 57306 0 57418 800
rect 57950 0 58062 800
rect 59238 0 59350 800
rect 59882 0 59994 800
rect 60526 0 60638 800
rect 61170 0 61282 800
rect 61814 0 61926 800
rect 62458 0 62570 800
rect 63102 0 63214 800
rect 63746 0 63858 800
rect 64390 0 64502 800
rect 65678 0 65790 800
rect 66322 0 66434 800
rect 66966 0 67078 800
rect 67610 0 67722 800
rect 68254 0 68366 800
rect 68898 0 69010 800
rect 69542 0 69654 800
rect 70186 0 70298 800
rect 70830 0 70942 800
rect 72118 0 72230 800
rect 72762 0 72874 800
rect 73406 0 73518 800
<< obsm2 >>
rect 204 73144 578 73250
rect 802 73144 1222 73250
rect 1446 73144 2510 73250
rect 2734 73144 3154 73250
rect 3378 73144 3798 73250
rect 4022 73144 4442 73250
rect 4666 73144 5086 73250
rect 5310 73144 5730 73250
rect 5954 73144 6374 73250
rect 6598 73144 7018 73250
rect 7242 73144 7662 73250
rect 7886 73144 8950 73250
rect 9174 73144 9594 73250
rect 9818 73144 10238 73250
rect 10462 73144 10882 73250
rect 11106 73144 11526 73250
rect 11750 73144 12170 73250
rect 12394 73144 12814 73250
rect 13038 73144 13458 73250
rect 13682 73144 14102 73250
rect 14326 73144 15390 73250
rect 15614 73144 16034 73250
rect 16258 73144 16678 73250
rect 16902 73144 17322 73250
rect 17546 73144 17966 73250
rect 18190 73144 18610 73250
rect 18834 73144 19254 73250
rect 19478 73144 19898 73250
rect 20122 73144 20542 73250
rect 20766 73144 21830 73250
rect 22054 73144 22474 73250
rect 22698 73144 23118 73250
rect 23342 73144 23762 73250
rect 23986 73144 24406 73250
rect 24630 73144 25050 73250
rect 25274 73144 25694 73250
rect 25918 73144 26338 73250
rect 26562 73144 26982 73250
rect 27206 73144 28270 73250
rect 28494 73144 28914 73250
rect 29138 73144 29558 73250
rect 29782 73144 30202 73250
rect 30426 73144 30846 73250
rect 31070 73144 31490 73250
rect 31714 73144 32134 73250
rect 32358 73144 32778 73250
rect 33002 73144 33422 73250
rect 33646 73144 34710 73250
rect 34934 73144 35354 73250
rect 35578 73144 35998 73250
rect 36222 73144 36642 73250
rect 36866 73144 37286 73250
rect 37510 73144 37930 73250
rect 38154 73144 38574 73250
rect 38798 73144 39218 73250
rect 39442 73144 39862 73250
rect 40086 73144 40506 73250
rect 40730 73144 41794 73250
rect 42018 73144 42438 73250
rect 42662 73144 43082 73250
rect 43306 73144 43726 73250
rect 43950 73144 44370 73250
rect 44594 73144 45014 73250
rect 45238 73144 45658 73250
rect 45882 73144 46302 73250
rect 46526 73144 46946 73250
rect 47170 73144 48234 73250
rect 48458 73144 48878 73250
rect 49102 73144 49522 73250
rect 49746 73144 50166 73250
rect 50390 73144 50810 73250
rect 51034 73144 51454 73250
rect 51678 73144 52098 73250
rect 52322 73144 52742 73250
rect 52966 73144 53386 73250
rect 53610 73144 54674 73250
rect 54898 73144 55318 73250
rect 55542 73144 55962 73250
rect 56186 73144 56606 73250
rect 56830 73144 57250 73250
rect 57474 73144 57894 73250
rect 58118 73144 58538 73250
rect 58762 73144 59182 73250
rect 59406 73144 59826 73250
rect 60050 73144 61114 73250
rect 61338 73144 61758 73250
rect 61982 73144 62402 73250
rect 62626 73144 63046 73250
rect 63270 73144 63690 73250
rect 63914 73144 64334 73250
rect 64558 73144 64978 73250
rect 65202 73144 65622 73250
rect 65846 73144 66266 73250
rect 66490 73144 67554 73250
rect 67778 73144 68198 73250
rect 68422 73144 68842 73250
rect 69066 73144 69486 73250
rect 69710 73144 70130 73250
rect 70354 73144 70774 73250
rect 70998 73144 71418 73250
rect 71642 73144 72062 73250
rect 72286 73144 72706 73250
rect 72930 73144 73350 73250
rect 204 856 73488 73144
rect 204 31 578 856
rect 802 31 1222 856
rect 1446 31 1866 856
rect 2090 31 2510 856
rect 2734 31 3154 856
rect 3378 31 3798 856
rect 4022 31 4442 856
rect 4666 31 5086 856
rect 5310 31 5730 856
rect 5954 31 7018 856
rect 7242 31 7662 856
rect 7886 31 8306 856
rect 8530 31 8950 856
rect 9174 31 9594 856
rect 9818 31 10238 856
rect 10462 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12170 856
rect 12394 31 13458 856
rect 13682 31 14102 856
rect 14326 31 14746 856
rect 14970 31 15390 856
rect 15614 31 16034 856
rect 16258 31 16678 856
rect 16902 31 17322 856
rect 17546 31 17966 856
rect 18190 31 18610 856
rect 18834 31 19898 856
rect 20122 31 20542 856
rect 20766 31 21186 856
rect 21410 31 21830 856
rect 22054 31 22474 856
rect 22698 31 23118 856
rect 23342 31 23762 856
rect 23986 31 24406 856
rect 24630 31 25050 856
rect 25274 31 26338 856
rect 26562 31 26982 856
rect 27206 31 27626 856
rect 27850 31 28270 856
rect 28494 31 28914 856
rect 29138 31 29558 856
rect 29782 31 30202 856
rect 30426 31 30846 856
rect 31070 31 31490 856
rect 31714 31 32778 856
rect 33002 31 33422 856
rect 33646 31 34066 856
rect 34290 31 34710 856
rect 34934 31 35354 856
rect 35578 31 35998 856
rect 36222 31 36642 856
rect 36866 31 37286 856
rect 37510 31 37930 856
rect 38154 31 38574 856
rect 38798 31 39862 856
rect 40086 31 40506 856
rect 40730 31 41150 856
rect 41374 31 41794 856
rect 42018 31 42438 856
rect 42662 31 43082 856
rect 43306 31 43726 856
rect 43950 31 44370 856
rect 44594 31 45014 856
rect 45238 31 46302 856
rect 46526 31 46946 856
rect 47170 31 47590 856
rect 47814 31 48234 856
rect 48458 31 48878 856
rect 49102 31 49522 856
rect 49746 31 50166 856
rect 50390 31 50810 856
rect 51034 31 51454 856
rect 51678 31 52742 856
rect 52966 31 53386 856
rect 53610 31 54030 856
rect 54254 31 54674 856
rect 54898 31 55318 856
rect 55542 31 55962 856
rect 56186 31 56606 856
rect 56830 31 57250 856
rect 57474 31 57894 856
rect 58118 31 59182 856
rect 59406 31 59826 856
rect 60050 31 60470 856
rect 60694 31 61114 856
rect 61338 31 61758 856
rect 61982 31 62402 856
rect 62626 31 63046 856
rect 63270 31 63690 856
rect 63914 31 64334 856
rect 64558 31 65622 856
rect 65846 31 66266 856
rect 66490 31 66910 856
rect 67134 31 67554 856
rect 67778 31 68198 856
rect 68422 31 68842 856
rect 69066 31 69486 856
rect 69710 31 70130 856
rect 70354 31 70774 856
rect 70998 31 72062 856
rect 72286 31 72706 856
rect 72930 31 73350 856
<< metal3 >>
rect 0 73388 800 73628
rect 0 72708 800 72948
rect 73200 72708 74000 72948
rect 0 72028 800 72268
rect 73200 72028 74000 72268
rect 0 71348 800 71588
rect 73200 71348 74000 71588
rect 0 70668 800 70908
rect 73200 70668 74000 70908
rect 0 69988 800 70228
rect 73200 69988 74000 70228
rect 0 69308 800 69548
rect 73200 69308 74000 69548
rect 73200 68628 74000 68868
rect 0 67948 800 68188
rect 73200 67948 74000 68188
rect 0 67268 800 67508
rect 73200 67268 74000 67508
rect 0 66588 800 66828
rect 0 65908 800 66148
rect 73200 65908 74000 66148
rect 0 65228 800 65468
rect 73200 65228 74000 65468
rect 0 64548 800 64788
rect 73200 64548 74000 64788
rect 0 63868 800 64108
rect 73200 63868 74000 64108
rect 0 63188 800 63428
rect 73200 63188 74000 63428
rect 0 62508 800 62748
rect 73200 62508 74000 62748
rect 73200 61828 74000 62068
rect 0 61148 800 61388
rect 73200 61148 74000 61388
rect 0 60468 800 60708
rect 73200 60468 74000 60708
rect 0 59788 800 60028
rect 0 59108 800 59348
rect 73200 59108 74000 59348
rect 0 58428 800 58668
rect 73200 58428 74000 58668
rect 0 57748 800 57988
rect 73200 57748 74000 57988
rect 0 57068 800 57308
rect 73200 57068 74000 57308
rect 0 56388 800 56628
rect 73200 56388 74000 56628
rect 0 55708 800 55948
rect 73200 55708 74000 55948
rect 73200 55028 74000 55268
rect 0 54348 800 54588
rect 73200 54348 74000 54588
rect 0 53668 800 53908
rect 73200 53668 74000 53908
rect 0 52988 800 53228
rect 0 52308 800 52548
rect 73200 52308 74000 52548
rect 0 51628 800 51868
rect 73200 51628 74000 51868
rect 0 50948 800 51188
rect 73200 50948 74000 51188
rect 0 50268 800 50508
rect 73200 50268 74000 50508
rect 0 49588 800 49828
rect 73200 49588 74000 49828
rect 0 48908 800 49148
rect 73200 48908 74000 49148
rect 73200 48228 74000 48468
rect 0 47548 800 47788
rect 73200 47548 74000 47788
rect 0 46868 800 47108
rect 73200 46868 74000 47108
rect 0 46188 800 46428
rect 0 45508 800 45748
rect 73200 45508 74000 45748
rect 0 44828 800 45068
rect 73200 44828 74000 45068
rect 0 44148 800 44388
rect 73200 44148 74000 44388
rect 0 43468 800 43708
rect 73200 43468 74000 43708
rect 0 42788 800 43028
rect 73200 42788 74000 43028
rect 0 42108 800 42348
rect 73200 42108 74000 42348
rect 73200 41428 74000 41668
rect 0 40748 800 40988
rect 73200 40748 74000 40988
rect 0 40068 800 40308
rect 73200 40068 74000 40308
rect 0 39388 800 39628
rect 0 38708 800 38948
rect 73200 38708 74000 38948
rect 0 38028 800 38268
rect 73200 38028 74000 38268
rect 0 37348 800 37588
rect 73200 37348 74000 37588
rect 0 36668 800 36908
rect 73200 36668 74000 36908
rect 0 35988 800 36228
rect 73200 35988 74000 36228
rect 0 35308 800 35548
rect 73200 35308 74000 35548
rect 0 34628 800 34868
rect 73200 34628 74000 34868
rect 73200 33948 74000 34188
rect 0 33268 800 33508
rect 73200 33268 74000 33508
rect 0 32588 800 32828
rect 73200 32588 74000 32828
rect 0 31908 800 32148
rect 0 31228 800 31468
rect 73200 31228 74000 31468
rect 0 30548 800 30788
rect 73200 30548 74000 30788
rect 0 29868 800 30108
rect 73200 29868 74000 30108
rect 0 29188 800 29428
rect 73200 29188 74000 29428
rect 0 28508 800 28748
rect 73200 28508 74000 28748
rect 0 27828 800 28068
rect 73200 27828 74000 28068
rect 73200 27148 74000 27388
rect 0 26468 800 26708
rect 73200 26468 74000 26708
rect 0 25788 800 26028
rect 73200 25788 74000 26028
rect 0 25108 800 25348
rect 0 24428 800 24668
rect 73200 24428 74000 24668
rect 0 23748 800 23988
rect 73200 23748 74000 23988
rect 0 23068 800 23308
rect 73200 23068 74000 23308
rect 0 22388 800 22628
rect 73200 22388 74000 22628
rect 0 21708 800 21948
rect 73200 21708 74000 21948
rect 0 21028 800 21268
rect 73200 21028 74000 21268
rect 73200 20348 74000 20588
rect 0 19668 800 19908
rect 73200 19668 74000 19908
rect 0 18988 800 19228
rect 73200 18988 74000 19228
rect 0 18308 800 18548
rect 0 17628 800 17868
rect 73200 17628 74000 17868
rect 0 16948 800 17188
rect 73200 16948 74000 17188
rect 0 16268 800 16508
rect 73200 16268 74000 16508
rect 0 15588 800 15828
rect 73200 15588 74000 15828
rect 0 14908 800 15148
rect 73200 14908 74000 15148
rect 0 14228 800 14468
rect 73200 14228 74000 14468
rect 73200 13548 74000 13788
rect 0 12868 800 13108
rect 73200 12868 74000 13108
rect 0 12188 800 12428
rect 73200 12188 74000 12428
rect 0 11508 800 11748
rect 0 10828 800 11068
rect 73200 10828 74000 11068
rect 0 10148 800 10388
rect 73200 10148 74000 10388
rect 0 9468 800 9708
rect 73200 9468 74000 9708
rect 0 8788 800 9028
rect 73200 8788 74000 9028
rect 0 8108 800 8348
rect 73200 8108 74000 8348
rect 0 7428 800 7668
rect 73200 7428 74000 7668
rect 73200 6748 74000 6988
rect 0 6068 800 6308
rect 73200 6068 74000 6308
rect 0 5388 800 5628
rect 73200 5388 74000 5628
rect 0 4708 800 4948
rect 0 4028 800 4268
rect 73200 4028 74000 4268
rect 0 3348 800 3588
rect 73200 3348 74000 3588
rect 0 2668 800 2908
rect 73200 2668 74000 2908
rect 0 1988 800 2228
rect 73200 1988 74000 2228
rect 0 1308 800 1548
rect 73200 1308 74000 1548
rect 0 628 800 868
rect 73200 628 74000 868
rect 73200 -52 74000 188
<< obsm3 >>
rect 880 72628 73120 72861
rect 800 72348 73200 72628
rect 880 71948 73120 72348
rect 800 71668 73200 71948
rect 880 71268 73120 71668
rect 800 70988 73200 71268
rect 880 70588 73120 70988
rect 800 70308 73200 70588
rect 880 69908 73120 70308
rect 800 69628 73200 69908
rect 880 69228 73120 69628
rect 800 68948 73200 69228
rect 800 68548 73120 68948
rect 800 68268 73200 68548
rect 880 67868 73120 68268
rect 800 67588 73200 67868
rect 880 67188 73120 67588
rect 800 66908 73200 67188
rect 880 66508 73200 66908
rect 800 66228 73200 66508
rect 880 65828 73120 66228
rect 800 65548 73200 65828
rect 880 65148 73120 65548
rect 800 64868 73200 65148
rect 880 64468 73120 64868
rect 800 64188 73200 64468
rect 880 63788 73120 64188
rect 800 63508 73200 63788
rect 880 63108 73120 63508
rect 800 62828 73200 63108
rect 880 62428 73120 62828
rect 800 62148 73200 62428
rect 800 61748 73120 62148
rect 800 61468 73200 61748
rect 880 61068 73120 61468
rect 800 60788 73200 61068
rect 880 60388 73120 60788
rect 800 60108 73200 60388
rect 880 59708 73200 60108
rect 800 59428 73200 59708
rect 880 59028 73120 59428
rect 800 58748 73200 59028
rect 880 58348 73120 58748
rect 800 58068 73200 58348
rect 880 57668 73120 58068
rect 800 57388 73200 57668
rect 880 56988 73120 57388
rect 800 56708 73200 56988
rect 880 56308 73120 56708
rect 800 56028 73200 56308
rect 880 55628 73120 56028
rect 800 55348 73200 55628
rect 800 54948 73120 55348
rect 800 54668 73200 54948
rect 880 54268 73120 54668
rect 800 53988 73200 54268
rect 880 53588 73120 53988
rect 800 53308 73200 53588
rect 880 52908 73200 53308
rect 800 52628 73200 52908
rect 880 52228 73120 52628
rect 800 51948 73200 52228
rect 880 51548 73120 51948
rect 800 51268 73200 51548
rect 880 50868 73120 51268
rect 800 50588 73200 50868
rect 880 50188 73120 50588
rect 800 49908 73200 50188
rect 880 49508 73120 49908
rect 800 49228 73200 49508
rect 880 48828 73120 49228
rect 800 48548 73200 48828
rect 800 48148 73120 48548
rect 800 47868 73200 48148
rect 880 47468 73120 47868
rect 800 47188 73200 47468
rect 880 46788 73120 47188
rect 800 46508 73200 46788
rect 880 46108 73200 46508
rect 800 45828 73200 46108
rect 880 45428 73120 45828
rect 800 45148 73200 45428
rect 880 44748 73120 45148
rect 800 44468 73200 44748
rect 880 44068 73120 44468
rect 800 43788 73200 44068
rect 880 43388 73120 43788
rect 800 43108 73200 43388
rect 880 42708 73120 43108
rect 800 42428 73200 42708
rect 880 42028 73120 42428
rect 800 41748 73200 42028
rect 800 41348 73120 41748
rect 800 41068 73200 41348
rect 880 40668 73120 41068
rect 800 40388 73200 40668
rect 880 39988 73120 40388
rect 800 39708 73200 39988
rect 880 39308 73200 39708
rect 800 39028 73200 39308
rect 880 38628 73120 39028
rect 800 38348 73200 38628
rect 880 37948 73120 38348
rect 800 37668 73200 37948
rect 880 37268 73120 37668
rect 800 36988 73200 37268
rect 880 36588 73120 36988
rect 800 36308 73200 36588
rect 880 35908 73120 36308
rect 800 35628 73200 35908
rect 880 35228 73120 35628
rect 800 34948 73200 35228
rect 880 34548 73120 34948
rect 800 34268 73200 34548
rect 800 33868 73120 34268
rect 800 33588 73200 33868
rect 880 33188 73120 33588
rect 800 32908 73200 33188
rect 880 32508 73120 32908
rect 800 32228 73200 32508
rect 880 31828 73200 32228
rect 800 31548 73200 31828
rect 880 31148 73120 31548
rect 800 30868 73200 31148
rect 880 30468 73120 30868
rect 800 30188 73200 30468
rect 880 29788 73120 30188
rect 800 29508 73200 29788
rect 880 29108 73120 29508
rect 800 28828 73200 29108
rect 880 28428 73120 28828
rect 800 28148 73200 28428
rect 880 27748 73120 28148
rect 800 27468 73200 27748
rect 800 27068 73120 27468
rect 800 26788 73200 27068
rect 880 26388 73120 26788
rect 800 26108 73200 26388
rect 880 25708 73120 26108
rect 800 25428 73200 25708
rect 880 25028 73200 25428
rect 800 24748 73200 25028
rect 880 24348 73120 24748
rect 800 24068 73200 24348
rect 880 23668 73120 24068
rect 800 23388 73200 23668
rect 880 22988 73120 23388
rect 800 22708 73200 22988
rect 880 22308 73120 22708
rect 800 22028 73200 22308
rect 880 21628 73120 22028
rect 800 21348 73200 21628
rect 880 20948 73120 21348
rect 800 20668 73200 20948
rect 800 20268 73120 20668
rect 800 19988 73200 20268
rect 880 19588 73120 19988
rect 800 19308 73200 19588
rect 880 18908 73120 19308
rect 800 18628 73200 18908
rect 880 18228 73200 18628
rect 800 17948 73200 18228
rect 880 17548 73120 17948
rect 800 17268 73200 17548
rect 880 16868 73120 17268
rect 800 16588 73200 16868
rect 880 16188 73120 16588
rect 800 15908 73200 16188
rect 880 15508 73120 15908
rect 800 15228 73200 15508
rect 880 14828 73120 15228
rect 800 14548 73200 14828
rect 880 14148 73120 14548
rect 800 13868 73200 14148
rect 800 13468 73120 13868
rect 800 13188 73200 13468
rect 880 12788 73120 13188
rect 800 12508 73200 12788
rect 880 12108 73120 12508
rect 800 11828 73200 12108
rect 880 11428 73200 11828
rect 800 11148 73200 11428
rect 880 10748 73120 11148
rect 800 10468 73200 10748
rect 880 10068 73120 10468
rect 800 9788 73200 10068
rect 880 9388 73120 9788
rect 800 9108 73200 9388
rect 880 8708 73120 9108
rect 800 8428 73200 8708
rect 880 8028 73120 8428
rect 800 7748 73200 8028
rect 880 7348 73120 7748
rect 800 7068 73200 7348
rect 800 6668 73120 7068
rect 800 6388 73200 6668
rect 880 5988 73120 6388
rect 800 5708 73200 5988
rect 880 5308 73120 5708
rect 800 5028 73200 5308
rect 880 4628 73200 5028
rect 800 4348 73200 4628
rect 880 3948 73120 4348
rect 800 3668 73200 3948
rect 880 3268 73120 3668
rect 800 2988 73200 3268
rect 880 2588 73120 2988
rect 800 2308 73200 2588
rect 880 1908 73120 2308
rect 800 1628 73200 1908
rect 880 1228 73120 1628
rect 800 948 73200 1228
rect 880 548 73120 948
rect 800 268 73200 548
rect 800 35 73120 268
<< metal4 >>
rect 4208 2128 4528 71856
rect 19568 2128 19888 71856
rect 34928 2128 35248 71856
rect 50288 2128 50608 71856
rect 65648 2128 65968 71856
<< obsm4 >>
rect 19379 3435 19488 35597
rect 19968 3435 34848 35597
rect 35328 3435 36925 35597
<< labels >>
rlabel metal3 s 73200 19668 74000 19908 6 active
port 1 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 72762 0 72874 800 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 73200 58428 74000 58668 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 73200 68628 74000 68868 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 50222 0 50334 800 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 73200 38708 74000 38948 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 73200 65908 74000 66148 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 66588 800 66828 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 38630 73200 38742 74000 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 38708 800 38948 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 41850 73200 41962 74000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 57306 73200 57418 74000 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 0 52988 800 53228 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 65678 73200 65790 74000 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 0 73388 800 73628 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 73200 72028 74000 72268 6 io_in[28]
port 22 nsew signal input
rlabel metal3 s 73200 50268 74000 50508 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 47646 0 47758 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 0 54348 800 54588 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 43138 73200 43250 74000 6 io_in[33]
port 28 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 73200 26468 74000 26708 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 0 46868 800 47108 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 58594 73200 58706 74000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 14158 73200 14270 74000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 45070 73200 45182 74000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 45714 73200 45826 74000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 5142 73200 5254 74000 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 73200 8108 74000 8348 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 72028 800 72268 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 65678 0 65790 800 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal3 s 73200 16268 74000 16508 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal3 s 0 24428 800 24668 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 73200 50948 74000 51188 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal2 s 48934 73200 49046 74000 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 71348 800 71588 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 23818 73200 23930 74000 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal2 s 57950 0 58062 800 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal3 s 73200 60468 74000 60708 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 10294 73200 10406 74000 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 0 50948 800 51188 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 0 69308 800 69548 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal3 s 73200 9468 74000 9708 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal2 s 34766 0 34878 800 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal2 s 634 73200 746 74000 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal3 s 73200 1988 74000 2228 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal3 s 0 72708 800 72948 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal3 s 0 18988 800 19228 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal3 s 0 46188 800 46428 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal3 s 73200 27148 74000 27388 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 0 35988 800 36228 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 44426 0 44538 800 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal2 s 64390 73200 64502 74000 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal3 s 73200 28508 74000 28748 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 68254 0 68366 800 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal2 s 43782 73200 43894 74000 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 0 52308 800 52548 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 42494 73200 42606 74000 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal3 s 0 26468 800 26708 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 73200 67268 74000 67508 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal2 s 12870 73200 12982 74000 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal3 s 73200 -52 74000 188 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 0 67948 800 68188 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 0 63868 800 64108 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 0 34628 800 34868 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 0 18308 800 18548 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 30258 73200 30370 74000 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 60526 0 60638 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal2 s 72118 73200 72230 74000 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal3 s 73200 51628 74000 51868 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal2 s 2566 73200 2678 74000 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal2 s 47002 73200 47114 74000 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal3 s 0 51628 800 51868 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal3 s 0 60468 800 60708 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 73200 70668 74000 70908 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal2 s 10938 73200 11050 74000 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal2 s 37986 73200 38098 74000 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal3 s 0 1988 800 2228 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal2 s 14158 0 14270 800 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 0 56388 800 56628 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal3 s 73200 37348 74000 37588 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal3 s 0 15588 800 15828 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal3 s 0 8108 800 8348 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal3 s 73200 3348 74000 3588 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 0 40068 800 40308 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 69542 0 69654 800 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal3 s 73200 64548 74000 64788 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal3 s 73200 21708 74000 21948 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 33478 0 33590 800 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 3854 73200 3966 74000 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal2 s 37342 73200 37454 74000 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal3 s 73200 53668 74000 53908 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal2 s 54730 73200 54842 74000 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal3 s 0 47548 800 47788 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal2 s 66966 0 67078 800 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal2 s 25106 0 25218 800 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal2 s 19310 73200 19422 74000 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal2 s 33478 73200 33590 74000 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal2 s 70186 73200 70298 74000 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal2 s 26394 73200 26506 74000 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal2 s 1278 73200 1390 74000 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal2 s 15446 73200 15558 74000 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 0 35308 800 35548 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal3 s 73200 12868 74000 13108 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal2 s 5786 73200 5898 74000 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal3 s 73200 7428 74000 7668 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal2 s 40562 73200 40674 74000 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 3210 73200 3322 74000 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 18666 73200 18778 74000 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 73200 12188 74000 12428 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal2 s 59882 0 59994 800 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 73200 15588 74000 15828 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 73200 10828 74000 11068 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 73200 27828 74000 28068 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 63102 73200 63214 74000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 66322 73200 66434 74000 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 73200 69308 74000 69548 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 73200 61828 74000 62068 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 64390 0 64502 800 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal2 s 50222 73200 50334 74000 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 56018 73200 56130 74000 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal2 s 61170 73200 61282 74000 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 71474 73200 71586 74000 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 73200 72708 74000 72948 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 73200 49588 74000 49828 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 0 44148 800 44388 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 4028 800 4268 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 52798 73200 52910 74000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal2 s 48934 0 49046 800 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal2 s 13514 73200 13626 74000 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 52798 0 52910 800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 32834 73200 32946 74000 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal2 s 31546 0 31658 800 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal3 s 0 11508 800 11748 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal3 s 73200 44828 74000 45068 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal3 s 73200 14908 74000 15148 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal3 s 0 21028 800 21268 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal2 s 46358 0 46470 800 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 0 61148 800 61388 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal2 s 24462 0 24574 800 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal2 s 29614 0 29726 800 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal2 s 11582 0 11694 800 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 73200 29868 74000 30108 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 31908 800 32148 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal3 s 0 67268 800 67508 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal3 s 0 31228 800 31468 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 20598 73200 20710 74000 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal3 s 0 70668 800 70908 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 73200 59108 74000 59348 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal2 s 68898 73200 69010 74000 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 73200 32588 74000 32828 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal2 s 44426 73200 44538 74000 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal3 s 0 39388 800 39628 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 21886 0 21998 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal2 s 26394 0 26506 800 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 73200 25788 74000 26028 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 0 29868 800 30108 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal2 s 18022 73200 18134 74000 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 39918 73200 40030 74000 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal3 s 73200 55708 74000 55948 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal2 s 31546 73200 31658 74000 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal3 s 73200 63868 74000 64108 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal3 s 73200 5388 74000 5628 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal2 s 61814 73200 61926 74000 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 0 1308 800 1548 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 37342 0 37454 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s 16734 73200 16846 74000 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 9650 0 9762 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal2 s 7074 73200 7186 74000 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 9006 73200 9118 74000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 59108 800 59348 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 28970 73200 29082 74000 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 0 58428 800 58668 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 73200 8788 74000 9028 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 73200 55028 74000 55268 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 73200 24428 74000 24668 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal2 s 70830 0 70942 800 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal2 s 29614 73200 29726 74000 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 55374 73200 55486 74000 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 0 3348 800 3588 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 53668 800 53908 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal2 s 36698 73200 36810 74000 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 3854 0 3966 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 0 4708 800 4948 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal2 s 63746 0 63858 800 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 0 55708 800 55948 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal2 s 63102 0 63214 800 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 73200 33948 74000 34188 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal2 s 16090 73200 16202 74000 6 la2_data_in[0]
port 212 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la2_data_in[10]
port 213 nsew signal input
rlabel metal3 s 0 33268 800 33508 6 la2_data_in[11]
port 214 nsew signal input
rlabel metal3 s 0 64548 800 64788 6 la2_data_in[12]
port 215 nsew signal input
rlabel metal2 s 22530 73200 22642 74000 6 la2_data_in[13]
port 216 nsew signal input
rlabel metal2 s 35410 73200 35522 74000 6 la2_data_in[14]
port 217 nsew signal input
rlabel metal3 s 73200 13548 74000 13788 6 la2_data_in[15]
port 218 nsew signal input
rlabel metal2 s 59882 73200 59994 74000 6 la2_data_in[16]
port 219 nsew signal input
rlabel metal3 s 73200 47548 74000 47788 6 la2_data_in[17]
port 220 nsew signal input
rlabel metal3 s 73200 62508 74000 62748 6 la2_data_in[18]
port 221 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la2_data_in[19]
port 222 nsew signal input
rlabel metal2 s 25750 73200 25862 74000 6 la2_data_in[1]
port 223 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la2_data_in[20]
port 224 nsew signal input
rlabel metal2 s 61170 0 61282 800 6 la2_data_in[21]
port 225 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la2_data_in[22]
port 226 nsew signal input
rlabel metal3 s 73200 16948 74000 17188 6 la2_data_in[23]
port 227 nsew signal input
rlabel metal2 s 73406 73200 73518 74000 6 la2_data_in[24]
port 228 nsew signal input
rlabel metal2 s 43782 0 43894 800 6 la2_data_in[25]
port 229 nsew signal input
rlabel metal3 s 73200 31228 74000 31468 6 la2_data_in[26]
port 230 nsew signal input
rlabel metal3 s 73200 23748 74000 23988 6 la2_data_in[27]
port 231 nsew signal input
rlabel metal3 s 73200 48908 74000 49148 6 la2_data_in[28]
port 232 nsew signal input
rlabel metal3 s 73200 38028 74000 38268 6 la2_data_in[29]
port 233 nsew signal input
rlabel metal2 s 32190 73200 32302 74000 6 la2_data_in[2]
port 234 nsew signal input
rlabel metal3 s 73200 40068 74000 40308 6 la2_data_in[30]
port 235 nsew signal input
rlabel metal3 s 0 2668 800 2908 6 la2_data_in[31]
port 236 nsew signal input
rlabel metal2 s 61814 0 61926 800 6 la2_data_in[3]
port 237 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la2_data_in[4]
port 238 nsew signal input
rlabel metal3 s 0 48908 800 49148 6 la2_data_in[5]
port 239 nsew signal input
rlabel metal2 s 56018 0 56130 800 6 la2_data_in[6]
port 240 nsew signal input
rlabel metal3 s 73200 2668 74000 2908 6 la2_data_in[7]
port 241 nsew signal input
rlabel metal2 s 12226 73200 12338 74000 6 la2_data_in[8]
port 242 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la2_data_in[9]
port 243 nsew signal input
rlabel metal2 s 34766 73200 34878 74000 6 la2_data_out[0]
port 244 nsew signal bidirectional
rlabel metal3 s 0 57748 800 57988 6 la2_data_out[10]
port 245 nsew signal bidirectional
rlabel metal2 s 19954 0 20066 800 6 la2_data_out[11]
port 246 nsew signal bidirectional
rlabel metal3 s 73200 42108 74000 42348 6 la2_data_out[12]
port 247 nsew signal bidirectional
rlabel metal2 s 62458 0 62570 800 6 la2_data_out[13]
port 248 nsew signal bidirectional
rlabel metal3 s 0 22388 800 22628 6 la2_data_out[14]
port 249 nsew signal bidirectional
rlabel metal2 s 12226 0 12338 800 6 la2_data_out[15]
port 250 nsew signal bidirectional
rlabel metal3 s 73200 35988 74000 36228 6 la2_data_out[16]
port 251 nsew signal bidirectional
rlabel metal3 s 0 25788 800 26028 6 la2_data_out[17]
port 252 nsew signal bidirectional
rlabel metal3 s 73200 71348 74000 71588 6 la2_data_out[18]
port 253 nsew signal bidirectional
rlabel metal3 s 73200 61148 74000 61388 6 la2_data_out[19]
port 254 nsew signal bidirectional
rlabel metal3 s 73200 57748 74000 57988 6 la2_data_out[1]
port 255 nsew signal bidirectional
rlabel metal3 s 73200 57068 74000 57308 6 la2_data_out[20]
port 256 nsew signal bidirectional
rlabel metal2 s 36054 0 36166 800 6 la2_data_out[21]
port 257 nsew signal bidirectional
rlabel metal2 s 68254 73200 68366 74000 6 la2_data_out[22]
port 258 nsew signal bidirectional
rlabel metal2 s 1922 0 2034 800 6 la2_data_out[23]
port 259 nsew signal bidirectional
rlabel metal2 s 634 0 746 800 6 la2_data_out[24]
port 260 nsew signal bidirectional
rlabel metal2 s 4498 73200 4610 74000 6 la2_data_out[25]
port 261 nsew signal bidirectional
rlabel metal2 s 36698 0 36810 800 6 la2_data_out[26]
port 262 nsew signal bidirectional
rlabel metal2 s 73406 0 73518 800 6 la2_data_out[27]
port 263 nsew signal bidirectional
rlabel metal2 s 72762 73200 72874 74000 6 la2_data_out[28]
port 264 nsew signal bidirectional
rlabel metal3 s 73200 6068 74000 6308 6 la2_data_out[29]
port 265 nsew signal bidirectional
rlabel metal2 s 30902 73200 31014 74000 6 la2_data_out[2]
port 266 nsew signal bidirectional
rlabel metal3 s 0 49588 800 49828 6 la2_data_out[30]
port 267 nsew signal bidirectional
rlabel metal2 s 13514 0 13626 800 6 la2_data_out[31]
port 268 nsew signal bidirectional
rlabel metal2 s 30902 0 31014 800 6 la2_data_out[3]
port 269 nsew signal bidirectional
rlabel metal2 s 63746 73200 63858 74000 6 la2_data_out[4]
port 270 nsew signal bidirectional
rlabel metal3 s 0 19668 800 19908 6 la2_data_out[5]
port 271 nsew signal bidirectional
rlabel metal2 s 27038 0 27150 800 6 la2_data_out[6]
port 272 nsew signal bidirectional
rlabel metal3 s 0 57068 800 57308 6 la2_data_out[7]
port 273 nsew signal bidirectional
rlabel metal3 s 73200 33268 74000 33508 6 la2_data_out[8]
port 274 nsew signal bidirectional
rlabel metal3 s 73200 46868 74000 47108 6 la2_data_out[9]
port 275 nsew signal bidirectional
rlabel metal2 s 54730 0 54842 800 6 la2_oenb[0]
port 276 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la2_oenb[10]
port 277 nsew signal input
rlabel metal2 s 70186 0 70298 800 6 la2_oenb[11]
port 278 nsew signal input
rlabel metal3 s 73200 44148 74000 44388 6 la2_oenb[12]
port 279 nsew signal input
rlabel metal2 s 52154 73200 52266 74000 6 la2_oenb[13]
port 280 nsew signal input
rlabel metal3 s 0 628 800 868 6 la2_oenb[14]
port 281 nsew signal input
rlabel metal2 s 54086 0 54198 800 6 la2_oenb[15]
port 282 nsew signal input
rlabel metal2 s 67610 73200 67722 74000 6 la2_oenb[16]
port 283 nsew signal input
rlabel metal3 s 73200 4028 74000 4268 6 la2_oenb[17]
port 284 nsew signal input
rlabel metal2 s 46358 73200 46470 74000 6 la2_oenb[18]
port 285 nsew signal input
rlabel metal2 s 66322 0 66434 800 6 la2_oenb[19]
port 286 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 la2_oenb[1]
port 287 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la2_oenb[20]
port 288 nsew signal input
rlabel metal3 s 73200 34628 74000 34868 6 la2_oenb[21]
port 289 nsew signal input
rlabel metal2 s -10 73200 102 74000 6 la2_oenb[22]
port 290 nsew signal input
rlabel metal3 s 73200 45508 74000 45748 6 la2_oenb[23]
port 291 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la2_oenb[24]
port 292 nsew signal input
rlabel metal2 s 67610 0 67722 800 6 la2_oenb[25]
port 293 nsew signal input
rlabel metal2 s 24462 73200 24574 74000 6 la2_oenb[26]
port 294 nsew signal input
rlabel metal2 s 65034 73200 65146 74000 6 la2_oenb[27]
port 295 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la2_oenb[28]
port 296 nsew signal input
rlabel metal3 s 0 17628 800 17868 6 la2_oenb[29]
port 297 nsew signal input
rlabel metal2 s 28326 73200 28438 74000 6 la2_oenb[2]
port 298 nsew signal input
rlabel metal3 s 73200 10148 74000 10388 6 la2_oenb[30]
port 299 nsew signal input
rlabel metal2 s 17378 73200 17490 74000 6 la2_oenb[31]
port 300 nsew signal input
rlabel metal3 s 73200 23068 74000 23308 6 la2_oenb[3]
port 301 nsew signal input
rlabel metal2 s 50866 73200 50978 74000 6 la2_oenb[4]
port 302 nsew signal input
rlabel metal2 s 36054 73200 36166 74000 6 la2_oenb[5]
port 303 nsew signal input
rlabel metal2 s 7718 73200 7830 74000 6 la2_oenb[6]
port 304 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la2_oenb[7]
port 305 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la2_oenb[8]
port 306 nsew signal input
rlabel metal3 s 73200 52308 74000 52548 6 la2_oenb[9]
port 307 nsew signal input
rlabel metal3 s 73200 48228 74000 48468 6 la3_data_in[0]
port 308 nsew signal input
rlabel metal2 s 45070 0 45182 800 6 la3_data_in[10]
port 309 nsew signal input
rlabel metal3 s 0 43468 800 43708 6 la3_data_in[11]
port 310 nsew signal input
rlabel metal3 s 73200 21028 74000 21268 6 la3_data_in[12]
port 311 nsew signal input
rlabel metal2 s 68898 0 69010 800 6 la3_data_in[13]
port 312 nsew signal input
rlabel metal3 s 0 5388 800 5628 6 la3_data_in[14]
port 313 nsew signal input
rlabel metal3 s 0 42108 800 42348 6 la3_data_in[15]
port 314 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la3_data_in[16]
port 315 nsew signal input
rlabel metal2 s 57306 0 57418 800 6 la3_data_in[17]
port 316 nsew signal input
rlabel metal3 s 73200 14228 74000 14468 6 la3_data_in[18]
port 317 nsew signal input
rlabel metal2 s 11582 73200 11694 74000 6 la3_data_in[19]
port 318 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 la3_data_in[1]
port 319 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la3_data_in[20]
port 320 nsew signal input
rlabel metal2 s 27038 73200 27150 74000 6 la3_data_in[21]
port 321 nsew signal input
rlabel metal3 s 73200 41428 74000 41668 6 la3_data_in[22]
port 322 nsew signal input
rlabel metal3 s 73200 69988 74000 70228 6 la3_data_in[23]
port 323 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la3_data_in[24]
port 324 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la3_data_in[25]
port 325 nsew signal input
rlabel metal3 s 73200 29188 74000 29428 6 la3_data_in[26]
port 326 nsew signal input
rlabel metal2 s 55374 0 55486 800 6 la3_data_in[27]
port 327 nsew signal input
rlabel metal2 s 57950 73200 58062 74000 6 la3_data_in[28]
port 328 nsew signal input
rlabel metal2 s 53442 0 53554 800 6 la3_data_in[29]
port 329 nsew signal input
rlabel metal3 s 0 37348 800 37588 6 la3_data_in[2]
port 330 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la3_data_in[30]
port 331 nsew signal input
rlabel metal2 s 72118 0 72230 800 6 la3_data_in[31]
port 332 nsew signal input
rlabel metal3 s 73200 17628 74000 17868 6 la3_data_in[3]
port 333 nsew signal input
rlabel metal2 s 25106 73200 25218 74000 6 la3_data_in[4]
port 334 nsew signal input
rlabel metal3 s 73200 63188 74000 63428 6 la3_data_in[5]
port 335 nsew signal input
rlabel metal3 s 0 59788 800 60028 6 la3_data_in[6]
port 336 nsew signal input
rlabel metal3 s 0 65228 800 65468 6 la3_data_in[7]
port 337 nsew signal input
rlabel metal3 s 0 63188 800 63428 6 la3_data_in[8]
port 338 nsew signal input
rlabel metal2 s 2566 0 2678 800 6 la3_data_in[9]
port 339 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la3_data_out[0]
port 340 nsew signal bidirectional
rlabel metal3 s 73200 36668 74000 36908 6 la3_data_out[10]
port 341 nsew signal bidirectional
rlabel metal2 s 41206 0 41318 800 6 la3_data_out[11]
port 342 nsew signal bidirectional
rlabel metal3 s 0 12188 800 12428 6 la3_data_out[12]
port 343 nsew signal bidirectional
rlabel metal2 s 69542 73200 69654 74000 6 la3_data_out[13]
port 344 nsew signal bidirectional
rlabel metal2 s 6430 73200 6542 74000 6 la3_data_out[14]
port 345 nsew signal bidirectional
rlabel metal3 s 0 32588 800 32828 6 la3_data_out[15]
port 346 nsew signal bidirectional
rlabel metal3 s 73200 42788 74000 43028 6 la3_data_out[16]
port 347 nsew signal bidirectional
rlabel metal2 s 70830 73200 70942 74000 6 la3_data_out[17]
port 348 nsew signal bidirectional
rlabel metal3 s 0 45508 800 45748 6 la3_data_out[18]
port 349 nsew signal bidirectional
rlabel metal3 s 0 10148 800 10388 6 la3_data_out[19]
port 350 nsew signal bidirectional
rlabel metal3 s 73200 22388 74000 22628 6 la3_data_out[1]
port 351 nsew signal bidirectional
rlabel metal2 s 49578 0 49690 800 6 la3_data_out[20]
port 352 nsew signal bidirectional
rlabel metal2 s 62458 73200 62570 74000 6 la3_data_out[21]
port 353 nsew signal bidirectional
rlabel metal2 s 19954 73200 20066 74000 6 la3_data_out[22]
port 354 nsew signal bidirectional
rlabel metal2 s 22530 0 22642 800 6 la3_data_out[23]
port 355 nsew signal bidirectional
rlabel metal3 s 73200 43468 74000 43708 6 la3_data_out[24]
port 356 nsew signal bidirectional
rlabel metal2 s 59238 0 59350 800 6 la3_data_out[25]
port 357 nsew signal bidirectional
rlabel metal3 s 73200 20348 74000 20588 6 la3_data_out[26]
port 358 nsew signal bidirectional
rlabel metal3 s 0 40748 800 40988 6 la3_data_out[27]
port 359 nsew signal bidirectional
rlabel metal3 s 73200 628 74000 868 6 la3_data_out[28]
port 360 nsew signal bidirectional
rlabel metal2 s 10938 0 11050 800 6 la3_data_out[29]
port 361 nsew signal bidirectional
rlabel metal2 s 35410 0 35522 800 6 la3_data_out[2]
port 362 nsew signal bidirectional
rlabel metal3 s 73200 30548 74000 30788 6 la3_data_out[30]
port 363 nsew signal bidirectional
rlabel metal2 s 59238 73200 59350 74000 6 la3_data_out[31]
port 364 nsew signal bidirectional
rlabel metal3 s 73200 65228 74000 65468 6 la3_data_out[3]
port 365 nsew signal bidirectional
rlabel metal3 s 73200 1308 74000 1548 6 la3_data_out[4]
port 366 nsew signal bidirectional
rlabel metal2 s 5142 0 5254 800 6 la3_data_out[5]
port 367 nsew signal bidirectional
rlabel metal3 s 73200 40748 74000 40988 6 la3_data_out[6]
port 368 nsew signal bidirectional
rlabel metal2 s 1278 0 1390 800 6 la3_data_out[7]
port 369 nsew signal bidirectional
rlabel metal3 s 73200 67948 74000 68188 6 la3_data_out[8]
port 370 nsew signal bidirectional
rlabel metal2 s 56662 73200 56774 74000 6 la3_data_out[9]
port 371 nsew signal bidirectional
rlabel metal3 s 73200 6748 74000 6988 6 la3_oenb[0]
port 372 nsew signal input
rlabel metal2 s 53442 73200 53554 74000 6 la3_oenb[10]
port 373 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 la3_oenb[11]
port 374 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la3_oenb[12]
port 375 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la3_oenb[13]
port 376 nsew signal input
rlabel metal2 s -10 0 102 800 6 la3_oenb[14]
port 377 nsew signal input
rlabel metal2 s 56662 0 56774 800 6 la3_oenb[15]
port 378 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 la3_oenb[16]
port 379 nsew signal input
rlabel metal3 s 0 65908 800 66148 6 la3_oenb[17]
port 380 nsew signal input
rlabel metal2 s 21886 73200 21998 74000 6 la3_oenb[18]
port 381 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la3_oenb[19]
port 382 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 la3_oenb[1]
port 383 nsew signal input
rlabel metal2 s 4498 0 4610 800 6 la3_oenb[20]
port 384 nsew signal input
rlabel metal2 s 39274 73200 39386 74000 6 la3_oenb[21]
port 385 nsew signal input
rlabel metal2 s 23174 73200 23286 74000 6 la3_oenb[22]
port 386 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 la3_oenb[23]
port 387 nsew signal input
rlabel metal2 s 51510 73200 51622 74000 6 la3_oenb[24]
port 388 nsew signal input
rlabel metal3 s 73200 18988 74000 19228 6 la3_oenb[25]
port 389 nsew signal input
rlabel metal3 s 0 50268 800 50508 6 la3_oenb[26]
port 390 nsew signal input
rlabel metal3 s 73200 56388 74000 56628 6 la3_oenb[27]
port 391 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la3_oenb[28]
port 392 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la3_oenb[29]
port 393 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la3_oenb[2]
port 394 nsew signal input
rlabel metal3 s 73200 54348 74000 54588 6 la3_oenb[30]
port 395 nsew signal input
rlabel metal2 s 43138 0 43250 800 6 la3_oenb[31]
port 396 nsew signal input
rlabel metal2 s 49578 73200 49690 74000 6 la3_oenb[3]
port 397 nsew signal input
rlabel metal2 s 48290 73200 48402 74000 6 la3_oenb[4]
port 398 nsew signal input
rlabel metal3 s 0 69988 800 70228 6 la3_oenb[5]
port 399 nsew signal input
rlabel metal2 s 9650 73200 9762 74000 6 la3_oenb[6]
port 400 nsew signal input
rlabel metal2 s 51510 0 51622 800 6 la3_oenb[7]
port 401 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la3_oenb[8]
port 402 nsew signal input
rlabel metal3 s 0 62508 800 62748 6 la3_oenb[9]
port 403 nsew signal input
rlabel metal4 s 4208 2128 4528 71856 6 vccd1
port 404 nsew power input
rlabel metal4 s 34928 2128 35248 71856 6 vccd1
port 404 nsew power input
rlabel metal4 s 65648 2128 65968 71856 6 vccd1
port 404 nsew power input
rlabel metal4 s 19568 2128 19888 71856 6 vssd1
port 405 nsew ground input
rlabel metal4 s 50288 2128 50608 71856 6 vssd1
port 405 nsew ground input
rlabel metal3 s 73200 35308 74000 35548 6 wb_clk_i
port 406 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 74000 74000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6338560
string GDS_FILE /openlane/designs/wrapped_instrumented_adder_ripple/runs/RUN_2022.06.07_13.34.55/results/finishing/wrapped_instrumented_adder_ripple.magic.gds
string GDS_START 659876
<< end >>

